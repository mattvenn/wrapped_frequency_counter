magic
tech sky130A
magscale 1 2
timestamp 1671727933
<< viali >>
rect 23857 47141 23891 47175
rect 27353 47141 27387 47175
rect 10333 47073 10367 47107
rect 26157 47073 26191 47107
rect 2237 47005 2271 47039
rect 2881 47005 2915 47039
rect 5825 47005 5859 47039
rect 6561 47005 6595 47039
rect 7941 47005 7975 47039
rect 9321 47005 9355 47039
rect 13001 47005 13035 47039
rect 18337 47005 18371 47039
rect 22937 47005 22971 47039
rect 24041 47005 24075 47039
rect 26617 47005 26651 47039
rect 27445 47005 27479 47039
rect 27905 47005 27939 47039
rect 9505 46937 9539 46971
rect 26433 46937 26467 46971
rect 2789 46869 2823 46903
rect 6009 46869 6043 46903
rect 6745 46869 6779 46903
rect 26433 46665 26467 46699
rect 2513 46597 2547 46631
rect 2329 46529 2363 46563
rect 7021 46529 7055 46563
rect 12909 46529 12943 46563
rect 15853 46529 15887 46563
rect 18245 46529 18279 46563
rect 22845 46529 22879 46563
rect 26525 46529 26559 46563
rect 27813 46529 27847 46563
rect 2789 46461 2823 46495
rect 7205 46461 7239 46495
rect 8401 46461 8435 46495
rect 9321 46461 9355 46495
rect 9505 46461 9539 46495
rect 10977 46461 11011 46495
rect 13093 46461 13127 46495
rect 13553 46461 13587 46495
rect 16865 46461 16899 46495
rect 18429 46461 18463 46495
rect 18705 46461 18739 46495
rect 23029 46461 23063 46495
rect 23489 46461 23523 46495
rect 25881 46461 25915 46495
rect 1685 46325 1719 46359
rect 11713 46325 11747 46359
rect 15945 46325 15979 46359
rect 20545 46325 20579 46359
rect 27169 46325 27203 46359
rect 27905 46325 27939 46359
rect 7941 46121 7975 46155
rect 9505 46121 9539 46155
rect 10149 46121 10183 46155
rect 18429 46121 18463 46155
rect 23121 46121 23155 46155
rect 1593 45985 1627 46019
rect 4445 45985 4479 46019
rect 11345 45985 11379 46019
rect 11805 45985 11839 46019
rect 15945 45985 15979 46019
rect 16129 45985 16163 46019
rect 16773 45985 16807 46019
rect 20269 45985 20303 46019
rect 21281 45985 21315 46019
rect 26525 45985 26559 46019
rect 27721 45985 27755 46019
rect 3433 45917 3467 45951
rect 3985 45917 4019 45951
rect 8033 45917 8067 45951
rect 9413 45917 9447 45951
rect 10241 45917 10275 45951
rect 10701 45917 10735 45951
rect 14289 45917 14323 45951
rect 18337 45917 18371 45951
rect 23213 45917 23247 45951
rect 25237 45917 25271 45951
rect 25881 45917 25915 45951
rect 3249 45849 3283 45883
rect 4169 45849 4203 45883
rect 10793 45849 10827 45883
rect 11529 45849 11563 45883
rect 20453 45849 20487 45883
rect 25973 45849 26007 45883
rect 26709 45849 26743 45883
rect 13185 45577 13219 45611
rect 20453 45577 20487 45611
rect 4077 45509 4111 45543
rect 26433 45509 26467 45543
rect 1685 45441 1719 45475
rect 3985 45441 4019 45475
rect 9689 45441 9723 45475
rect 10425 45441 10459 45475
rect 13277 45441 13311 45475
rect 14197 45441 14231 45475
rect 20361 45441 20395 45475
rect 26617 45441 26651 45475
rect 1869 45373 1903 45407
rect 2145 45373 2179 45407
rect 14381 45373 14415 45407
rect 15209 45373 15243 45407
rect 26065 45373 26099 45407
rect 27905 45237 27939 45271
rect 2053 45033 2087 45067
rect 3341 45033 3375 45067
rect 27537 44897 27571 44931
rect 28365 44897 28399 44931
rect 2145 44829 2179 44863
rect 26065 44829 26099 44863
rect 28181 44761 28215 44795
rect 2145 44489 2179 44523
rect 14289 44489 14323 44523
rect 27905 44489 27939 44523
rect 24961 44421 24995 44455
rect 2237 44353 2271 44387
rect 14197 44353 14231 44387
rect 27169 44353 27203 44387
rect 27813 44353 27847 44387
rect 24777 44285 24811 44319
rect 26157 44285 26191 44319
rect 2973 44149 3007 44183
rect 27261 44149 27295 44183
rect 2513 43945 2547 43979
rect 21281 43809 21315 43843
rect 26249 43809 26283 43843
rect 26433 43809 26467 43843
rect 28089 43809 28123 43843
rect 1685 43741 1719 43775
rect 3341 43741 3375 43775
rect 19441 43741 19475 43775
rect 19625 43673 19659 43707
rect 3249 43605 3283 43639
rect 19533 43401 19567 43435
rect 3157 43333 3191 43367
rect 2237 43265 2271 43299
rect 2973 43265 3007 43299
rect 19441 43265 19475 43299
rect 26157 43265 26191 43299
rect 4169 43197 4203 43231
rect 2145 43061 2179 43095
rect 26249 43061 26283 43095
rect 27169 43061 27203 43095
rect 28089 43061 28123 43095
rect 1593 42721 1627 42755
rect 1777 42721 1811 42755
rect 2789 42721 2823 42755
rect 26525 42721 26559 42755
rect 28365 42721 28399 42755
rect 26709 42585 26743 42619
rect 2697 42177 2731 42211
rect 27721 42177 27755 42211
rect 1685 41973 1719 42007
rect 2605 41973 2639 42007
rect 3341 41973 3375 42007
rect 27813 41973 27847 42007
rect 3249 41633 3283 41667
rect 3433 41633 3467 41667
rect 27537 41633 27571 41667
rect 28181 41633 28215 41667
rect 28365 41633 28399 41667
rect 1593 41565 1627 41599
rect 1685 41089 1719 41123
rect 27445 41089 27479 41123
rect 1869 41021 1903 41055
rect 2789 41021 2823 41055
rect 27537 40885 27571 40919
rect 28273 40885 28307 40919
rect 27537 40545 27571 40579
rect 28181 40545 28215 40579
rect 28365 40545 28399 40579
rect 1961 40477 1995 40511
rect 2421 40477 2455 40511
rect 17785 40477 17819 40511
rect 18613 40477 18647 40511
rect 18797 40477 18831 40511
rect 1869 40341 1903 40375
rect 17693 40341 17727 40375
rect 18705 40341 18739 40375
rect 18321 40137 18355 40171
rect 1869 40069 1903 40103
rect 3525 40069 3559 40103
rect 18521 40069 18555 40103
rect 17233 40001 17267 40035
rect 17509 40001 17543 40035
rect 17693 40001 17727 40035
rect 19625 40001 19659 40035
rect 1685 39933 1719 39967
rect 17417 39933 17451 39967
rect 19809 39933 19843 39967
rect 17325 39865 17359 39899
rect 18153 39865 18187 39899
rect 17049 39797 17083 39831
rect 18337 39797 18371 39831
rect 19441 39797 19475 39831
rect 27353 39797 27387 39831
rect 27997 39797 28031 39831
rect 2329 39593 2363 39627
rect 17509 39593 17543 39627
rect 18521 39525 18555 39559
rect 19901 39457 19935 39491
rect 26525 39457 26559 39491
rect 28365 39457 28399 39491
rect 1593 39389 1627 39423
rect 2421 39389 2455 39423
rect 17693 39389 17727 39423
rect 17785 39389 17819 39423
rect 18429 39389 18463 39423
rect 18613 39389 18647 39423
rect 18705 39389 18739 39423
rect 18889 39389 18923 39423
rect 19717 39389 19751 39423
rect 19809 39389 19843 39423
rect 19993 39389 20027 39423
rect 20177 39389 20211 39423
rect 20821 39389 20855 39423
rect 17509 39321 17543 39355
rect 26709 39321 26743 39355
rect 1777 39253 1811 39287
rect 18245 39253 18279 39287
rect 19533 39253 19567 39287
rect 20729 39253 20763 39287
rect 19073 39049 19107 39083
rect 19993 39049 20027 39083
rect 18337 38981 18371 39015
rect 19241 38981 19275 39015
rect 19441 38981 19475 39015
rect 26433 38981 26467 39015
rect 27813 38981 27847 39015
rect 18245 38913 18279 38947
rect 19901 38913 19935 38947
rect 20085 38913 20119 38947
rect 26617 38913 26651 38947
rect 27721 38913 27755 38947
rect 22017 38845 22051 38879
rect 22201 38845 22235 38879
rect 23489 38845 23523 38879
rect 26157 38845 26191 38879
rect 2145 38777 2179 38811
rect 2789 38709 2823 38743
rect 19257 38709 19291 38743
rect 17693 38505 17727 38539
rect 21373 38505 21407 38539
rect 15485 38369 15519 38403
rect 28273 38369 28307 38403
rect 1685 38301 1719 38335
rect 2973 38301 3007 38335
rect 15112 38311 15146 38345
rect 15209 38301 15243 38335
rect 16129 38301 16163 38335
rect 16221 38301 16255 38335
rect 16313 38301 16347 38335
rect 16497 38301 16531 38335
rect 17417 38301 17451 38335
rect 17509 38301 17543 38335
rect 17785 38301 17819 38335
rect 18245 38301 18279 38335
rect 21281 38301 21315 38335
rect 26525 38301 26559 38335
rect 15301 38233 15335 38267
rect 15485 38233 15519 38267
rect 26709 38233 26743 38267
rect 2881 38165 2915 38199
rect 15945 38165 15979 38199
rect 17233 38165 17267 38199
rect 18337 38165 18371 38199
rect 27905 37961 27939 37995
rect 3801 37893 3835 37927
rect 4537 37893 4571 37927
rect 16313 37893 16347 37927
rect 17003 37893 17037 37927
rect 17141 37893 17175 37927
rect 17233 37893 17267 37927
rect 19809 37893 19843 37927
rect 3985 37825 4019 37859
rect 4629 37825 4663 37859
rect 16037 37825 16071 37859
rect 16865 37825 16899 37859
rect 17325 37825 17359 37859
rect 18245 37825 18279 37859
rect 18429 37825 18463 37859
rect 18613 37825 18647 37859
rect 18797 37825 18831 37859
rect 19533 37825 19567 37859
rect 27169 37825 27203 37859
rect 27813 37825 27847 37859
rect 2789 37757 2823 37791
rect 16313 37757 16347 37791
rect 18521 37757 18555 37791
rect 19809 37757 19843 37791
rect 16129 37689 16163 37723
rect 17509 37621 17543 37655
rect 18061 37621 18095 37655
rect 19625 37621 19659 37655
rect 17141 37417 17175 37451
rect 17325 37417 17359 37451
rect 19533 37417 19567 37451
rect 20085 37417 20119 37451
rect 24777 37349 24811 37383
rect 3249 37281 3283 37315
rect 15485 37281 15519 37315
rect 20545 37281 20579 37315
rect 21189 37281 21223 37315
rect 23489 37281 23523 37315
rect 26341 37281 26375 37315
rect 1593 37213 1627 37247
rect 3433 37213 3467 37247
rect 3985 37213 4019 37247
rect 18159 37213 18193 37247
rect 18331 37213 18365 37247
rect 19625 37213 19659 37247
rect 20269 37213 20303 37247
rect 20361 37213 20395 37247
rect 20637 37213 20671 37247
rect 21097 37213 21131 37247
rect 21281 37213 21315 37247
rect 23397 37213 23431 37247
rect 24593 37213 24627 37247
rect 25881 37213 25915 37247
rect 28365 37213 28399 37247
rect 4169 37145 4203 37179
rect 5825 37145 5859 37179
rect 15669 37145 15703 37179
rect 16957 37145 16991 37179
rect 17173 37145 17207 37179
rect 26065 37145 26099 37179
rect 15577 37077 15611 37111
rect 16037 37077 16071 37111
rect 18245 37077 18279 37111
rect 22937 37077 22971 37111
rect 23305 37077 23339 37111
rect 28181 37077 28215 37111
rect 5273 36873 5307 36907
rect 15945 36873 15979 36907
rect 20821 36873 20855 36907
rect 25973 36873 26007 36907
rect 27261 36873 27295 36907
rect 3249 36805 3283 36839
rect 3893 36805 3927 36839
rect 21373 36805 21407 36839
rect 22293 36805 22327 36839
rect 1869 36737 1903 36771
rect 4537 36737 4571 36771
rect 5365 36737 5399 36771
rect 19073 36737 19107 36771
rect 19257 36737 19291 36771
rect 20177 36737 20211 36771
rect 20637 36737 20671 36771
rect 21281 36737 21315 36771
rect 22661 36737 22695 36771
rect 25881 36737 25915 36771
rect 27169 36737 27203 36771
rect 2513 36669 2547 36703
rect 16037 36669 16071 36703
rect 16221 36669 16255 36703
rect 20343 36669 20377 36703
rect 20454 36669 20488 36703
rect 20545 36601 20579 36635
rect 1777 36533 1811 36567
rect 15577 36533 15611 36567
rect 19257 36533 19291 36567
rect 27905 36533 27939 36567
rect 19809 36329 19843 36363
rect 20821 36329 20855 36363
rect 1593 36193 1627 36227
rect 1777 36193 1811 36227
rect 2789 36193 2823 36227
rect 26525 36193 26559 36227
rect 4261 36125 4295 36159
rect 16957 36125 16991 36159
rect 17141 36125 17175 36159
rect 19993 36125 20027 36159
rect 20085 36125 20119 36159
rect 20361 36125 20395 36159
rect 20821 36125 20855 36159
rect 21005 36125 21039 36159
rect 22753 36125 22787 36159
rect 28365 36125 28399 36159
rect 4905 36057 4939 36091
rect 20177 36057 20211 36091
rect 22937 36057 22971 36091
rect 26709 36057 26743 36091
rect 17049 35989 17083 36023
rect 23121 35989 23155 36023
rect 27261 35785 27295 35819
rect 2329 35717 2363 35751
rect 12725 35717 12759 35751
rect 3157 35649 3191 35683
rect 3801 35649 3835 35683
rect 5181 35649 5215 35683
rect 11989 35649 12023 35683
rect 15761 35649 15795 35683
rect 15945 35649 15979 35683
rect 16865 35649 16899 35683
rect 18153 35649 18187 35683
rect 18409 35649 18443 35683
rect 23029 35649 23063 35683
rect 26433 35649 26467 35683
rect 27353 35649 27387 35683
rect 4445 35581 4479 35615
rect 5733 35581 5767 35615
rect 15577 35581 15611 35615
rect 25697 35581 25731 35615
rect 19533 35513 19567 35547
rect 17049 35445 17083 35479
rect 22845 35445 22879 35479
rect 25145 35445 25179 35479
rect 26249 35445 26283 35479
rect 27997 35445 28031 35479
rect 18245 35241 18279 35275
rect 20821 35241 20855 35275
rect 21281 35241 21315 35275
rect 2881 35105 2915 35139
rect 4353 35105 4387 35139
rect 1685 35037 1719 35071
rect 2605 35037 2639 35071
rect 4169 35037 4203 35071
rect 16865 35037 16899 35071
rect 17132 35037 17166 35071
rect 19441 35037 19475 35071
rect 19697 35037 19731 35071
rect 22394 35037 22428 35071
rect 22661 35037 22695 35071
rect 26433 35037 26467 35071
rect 28273 35037 28307 35071
rect 26188 34969 26222 35003
rect 28028 34969 28062 35003
rect 25053 34901 25087 34935
rect 26893 34901 26927 34935
rect 18429 34697 18463 34731
rect 20529 34697 20563 34731
rect 23949 34697 23983 34731
rect 25237 34697 25271 34731
rect 20729 34629 20763 34663
rect 22836 34629 22870 34663
rect 26372 34629 26406 34663
rect 27169 34629 27203 34663
rect 1685 34561 1719 34595
rect 4169 34561 4203 34595
rect 15577 34561 15611 34595
rect 15669 34561 15703 34595
rect 17049 34561 17083 34595
rect 17316 34561 17350 34595
rect 26617 34561 26651 34595
rect 27721 34561 27755 34595
rect 1869 34493 1903 34527
rect 2789 34493 2823 34527
rect 4813 34493 4847 34527
rect 22569 34493 22603 34527
rect 20361 34425 20395 34459
rect 15853 34357 15887 34391
rect 20545 34357 20579 34391
rect 2145 34153 2179 34187
rect 20545 34153 20579 34187
rect 24685 34017 24719 34051
rect 27537 34017 27571 34051
rect 28365 34017 28399 34051
rect 2237 33949 2271 33983
rect 4813 33949 4847 33983
rect 16037 33949 16071 33983
rect 20637 33949 20671 33983
rect 21281 33949 21315 33983
rect 23673 33949 23707 33983
rect 23765 33949 23799 33983
rect 23949 33949 23983 33983
rect 24041 33949 24075 33983
rect 24952 33949 24986 33983
rect 4169 33881 4203 33915
rect 21526 33881 21560 33915
rect 28181 33881 28215 33915
rect 16221 33813 16255 33847
rect 22661 33813 22695 33847
rect 23489 33813 23523 33847
rect 26065 33813 26099 33847
rect 16313 33609 16347 33643
rect 21281 33609 21315 33643
rect 26249 33609 26283 33643
rect 26617 33609 26651 33643
rect 27537 33609 27571 33643
rect 28089 33609 28123 33643
rect 18162 33541 18196 33575
rect 27169 33541 27203 33575
rect 15761 33473 15795 33507
rect 16037 33473 16071 33507
rect 16129 33473 16163 33507
rect 21189 33473 21223 33507
rect 21373 33473 21407 33507
rect 23837 33473 23871 33507
rect 27353 33473 27387 33507
rect 27997 33473 28031 33507
rect 18429 33405 18463 33439
rect 23581 33405 23615 33439
rect 26065 33405 26099 33439
rect 26157 33405 26191 33439
rect 17049 33337 17083 33371
rect 15853 33269 15887 33303
rect 24961 33269 24995 33303
rect 16313 33065 16347 33099
rect 23397 33065 23431 33099
rect 24869 33065 24903 33099
rect 17049 32997 17083 33031
rect 20269 32929 20303 32963
rect 27537 32929 27571 32963
rect 16037 32861 16071 32895
rect 17141 32861 17175 32895
rect 20085 32861 20119 32895
rect 20177 32861 20211 32895
rect 20361 32861 20395 32895
rect 20545 32861 20579 32895
rect 23581 32861 23615 32895
rect 23857 32861 23891 32895
rect 24041 32861 24075 32895
rect 25881 32861 25915 32895
rect 28365 32861 28399 32895
rect 25053 32793 25087 32827
rect 28181 32793 28215 32827
rect 16497 32725 16531 32759
rect 19901 32725 19935 32759
rect 24685 32725 24719 32759
rect 24853 32725 24887 32759
rect 25697 32725 25731 32759
rect 21281 32521 21315 32555
rect 18797 32453 18831 32487
rect 19594 32453 19628 32487
rect 18705 32385 18739 32419
rect 18889 32385 18923 32419
rect 21189 32385 21223 32419
rect 21373 32385 21407 32419
rect 23121 32385 23155 32419
rect 25881 32385 25915 32419
rect 27445 32385 27479 32419
rect 12725 32317 12759 32351
rect 12909 32317 12943 32351
rect 13829 32317 13863 32351
rect 19349 32317 19383 32351
rect 20729 32249 20763 32283
rect 23305 32181 23339 32215
rect 25973 32181 26007 32215
rect 27905 32181 27939 32215
rect 12909 31977 12943 32011
rect 19441 31977 19475 32011
rect 20729 31977 20763 32011
rect 22569 31977 22603 32011
rect 28181 31977 28215 32011
rect 16681 31909 16715 31943
rect 16497 31841 16531 31875
rect 16957 31841 16991 31875
rect 17509 31841 17543 31875
rect 23673 31841 23707 31875
rect 25789 31841 25823 31875
rect 25973 31841 26007 31875
rect 27537 31841 27571 31875
rect 12817 31773 12851 31807
rect 16313 31773 16347 31807
rect 16589 31773 16623 31807
rect 16773 31773 16807 31807
rect 17417 31773 17451 31807
rect 17601 31773 17635 31807
rect 19717 31773 19751 31807
rect 19809 31773 19843 31807
rect 19901 31773 19935 31807
rect 20085 31773 20119 31807
rect 20545 31773 20579 31807
rect 20729 31773 20763 31807
rect 21189 31773 21223 31807
rect 21456 31773 21490 31807
rect 23210 31773 23244 31807
rect 23581 31773 23615 31807
rect 28089 31773 28123 31807
rect 24777 31705 24811 31739
rect 24961 31705 24995 31739
rect 23029 31637 23063 31671
rect 23213 31637 23247 31671
rect 16113 31433 16147 31467
rect 16957 31433 16991 31467
rect 22109 31433 22143 31467
rect 23213 31433 23247 31467
rect 23857 31433 23891 31467
rect 16313 31365 16347 31399
rect 18622 31365 18656 31399
rect 22937 31365 22971 31399
rect 24225 31365 24259 31399
rect 16865 31297 16899 31331
rect 17049 31297 17083 31331
rect 20177 31297 20211 31331
rect 22017 31297 22051 31331
rect 22201 31297 22235 31331
rect 22661 31297 22695 31331
rect 22845 31297 22879 31331
rect 23029 31297 23063 31331
rect 24041 31297 24075 31331
rect 26617 31297 26651 31331
rect 27721 31297 27755 31331
rect 18889 31229 18923 31263
rect 26157 31229 26191 31263
rect 26433 31229 26467 31263
rect 27813 31229 27847 31263
rect 15945 31161 15979 31195
rect 17509 31161 17543 31195
rect 16129 31093 16163 31127
rect 20269 31093 20303 31127
rect 16037 30889 16071 30923
rect 22661 30889 22695 30923
rect 23121 30889 23155 30923
rect 25789 30889 25823 30923
rect 23305 30753 23339 30787
rect 28273 30753 28307 30787
rect 16129 30685 16163 30719
rect 16681 30685 16715 30719
rect 16773 30685 16807 30719
rect 18337 30685 18371 30719
rect 22477 30685 22511 30719
rect 22661 30685 22695 30719
rect 23397 30685 23431 30719
rect 24777 30685 24811 30719
rect 24869 30685 24903 30719
rect 26433 30685 26467 30719
rect 18705 30617 18739 30651
rect 23673 30617 23707 30651
rect 23765 30617 23799 30651
rect 25421 30617 25455 30651
rect 25605 30617 25639 30651
rect 26617 30617 26651 30651
rect 16957 30549 16991 30583
rect 24593 30549 24627 30583
rect 20177 30345 20211 30379
rect 27261 30345 27295 30379
rect 19165 30277 19199 30311
rect 22017 30277 22051 30311
rect 16129 30209 16163 30243
rect 16313 30209 16347 30243
rect 17049 30209 17083 30243
rect 17233 30209 17267 30243
rect 17509 30209 17543 30243
rect 19073 30209 19107 30243
rect 19349 30209 19383 30243
rect 19809 30209 19843 30243
rect 19993 30209 20027 30243
rect 20269 30209 20303 30243
rect 22201 30209 22235 30243
rect 22293 30209 22327 30243
rect 23489 30209 23523 30243
rect 23673 30209 23707 30243
rect 24501 30209 24535 30243
rect 26065 30209 26099 30243
rect 26157 30209 26191 30243
rect 26341 30209 26375 30243
rect 27353 30209 27387 30243
rect 28365 30209 28399 30243
rect 1593 30141 1627 30175
rect 1869 30141 1903 30175
rect 17325 30141 17359 30175
rect 25145 30141 25179 30175
rect 25237 30141 25271 30175
rect 25605 30141 25639 30175
rect 16313 30073 16347 30107
rect 17141 30073 17175 30107
rect 24317 30073 24351 30107
rect 28181 30073 28215 30107
rect 16865 30005 16899 30039
rect 19349 30005 19383 30039
rect 22017 30005 22051 30039
rect 23305 30005 23339 30039
rect 23581 30005 23615 30039
rect 24961 30005 24995 30039
rect 26525 30005 26559 30039
rect 17325 29801 17359 29835
rect 20821 29801 20855 29835
rect 24961 29801 24995 29835
rect 26065 29801 26099 29835
rect 25697 29733 25731 29767
rect 24869 29665 24903 29699
rect 27537 29665 27571 29699
rect 16681 29597 16715 29631
rect 16865 29597 16899 29631
rect 18705 29597 18739 29631
rect 19441 29597 19475 29631
rect 19697 29597 19731 29631
rect 22661 29597 22695 29631
rect 24593 29597 24627 29631
rect 25881 29597 25915 29631
rect 26065 29597 26099 29631
rect 26525 29597 26559 29631
rect 16773 29529 16807 29563
rect 18438 29529 18472 29563
rect 22394 29529 22428 29563
rect 26709 29529 26743 29563
rect 21281 29461 21315 29495
rect 25145 29461 25179 29495
rect 20637 29257 20671 29291
rect 22661 29257 22695 29291
rect 23213 29257 23247 29291
rect 23857 29257 23891 29291
rect 25973 29257 26007 29291
rect 27353 29257 27387 29291
rect 19993 29189 20027 29223
rect 20545 29121 20579 29155
rect 22385 29121 22419 29155
rect 23121 29121 23155 29155
rect 23305 29121 23339 29155
rect 23765 29121 23799 29155
rect 23949 29121 23983 29155
rect 25697 29121 25731 29155
rect 27445 29121 27479 29155
rect 22017 29053 22051 29087
rect 22477 29053 22511 29087
rect 25973 29053 26007 29087
rect 25789 28985 25823 29019
rect 27905 28985 27939 29019
rect 18705 28917 18739 28951
rect 16865 28713 16899 28747
rect 24685 28713 24719 28747
rect 22477 28577 22511 28611
rect 26525 28577 26559 28611
rect 27445 28577 27479 28611
rect 18245 28509 18279 28543
rect 20821 28509 20855 28543
rect 24593 28509 24627 28543
rect 24685 28509 24719 28543
rect 15669 28441 15703 28475
rect 15853 28441 15887 28475
rect 17978 28441 18012 28475
rect 23121 28441 23155 28475
rect 26709 28441 26743 28475
rect 16037 28373 16071 28407
rect 23213 28373 23247 28407
rect 24961 28373 24995 28407
rect 17049 28169 17083 28203
rect 22477 28169 22511 28203
rect 23397 28169 23431 28203
rect 27353 28169 27387 28203
rect 23565 28101 23599 28135
rect 23765 28101 23799 28135
rect 1593 28033 1627 28067
rect 16865 28033 16899 28067
rect 22201 28033 22235 28067
rect 22293 28033 22327 28067
rect 24317 28033 24351 28067
rect 24501 28033 24535 28067
rect 24593 28033 24627 28067
rect 25504 28033 25538 28067
rect 27445 28033 27479 28067
rect 14289 27965 14323 27999
rect 15945 27965 15979 27999
rect 16129 27965 16163 27999
rect 24409 27965 24443 27999
rect 25237 27965 25271 27999
rect 1777 27829 1811 27863
rect 23581 27829 23615 27863
rect 24777 27829 24811 27863
rect 26617 27829 26651 27863
rect 28089 27829 28123 27863
rect 15945 27625 15979 27659
rect 25789 27625 25823 27659
rect 14473 27557 14507 27591
rect 15393 27489 15427 27523
rect 23949 27489 23983 27523
rect 27537 27489 27571 27523
rect 28365 27489 28399 27523
rect 14381 27421 14415 27455
rect 15577 27421 15611 27455
rect 16497 27421 16531 27455
rect 19441 27421 19475 27455
rect 25145 27421 25179 27455
rect 25329 27421 25363 27455
rect 25421 27421 25455 27455
rect 25513 27421 25547 27455
rect 15485 27353 15519 27387
rect 19708 27353 19742 27387
rect 23682 27353 23716 27387
rect 28181 27353 28215 27387
rect 16681 27285 16715 27319
rect 20821 27285 20855 27319
rect 22569 27285 22603 27319
rect 16313 27081 16347 27115
rect 20269 27081 20303 27115
rect 23213 27081 23247 27115
rect 24501 27081 24535 27115
rect 27813 27081 27847 27115
rect 21189 27013 21223 27047
rect 21373 27013 21407 27047
rect 15945 26945 15979 26979
rect 16129 26945 16163 26979
rect 17305 26945 17339 26979
rect 18889 26945 18923 26979
rect 19145 26945 19179 26979
rect 21465 26945 21499 26979
rect 22661 26945 22695 26979
rect 23121 26945 23155 26979
rect 23305 26945 23339 26979
rect 24409 26945 24443 26979
rect 24685 26945 24719 26979
rect 27721 26945 27755 26979
rect 17049 26877 17083 26911
rect 22017 26877 22051 26911
rect 22385 26877 22419 26911
rect 22477 26877 22511 26911
rect 24685 26809 24719 26843
rect 18429 26741 18463 26775
rect 21189 26741 21223 26775
rect 16221 26537 16255 26571
rect 19809 26537 19843 26571
rect 22017 26537 22051 26571
rect 24041 26537 24075 26571
rect 24869 26469 24903 26503
rect 15577 26401 15611 26435
rect 20637 26401 20671 26435
rect 24593 26401 24627 26435
rect 2237 26333 2271 26367
rect 15853 26333 15887 26367
rect 19993 26333 20027 26367
rect 20904 26333 20938 26367
rect 23857 26333 23891 26367
rect 24041 26333 24075 26367
rect 27353 26333 27387 26367
rect 15761 26265 15795 26299
rect 27086 26265 27120 26299
rect 2145 26197 2179 26231
rect 25053 26197 25087 26231
rect 25973 26197 26007 26231
rect 16313 25993 16347 26027
rect 18245 25993 18279 26027
rect 19809 25993 19843 26027
rect 22937 25993 22971 26027
rect 25145 25993 25179 26027
rect 1869 25925 1903 25959
rect 17110 25925 17144 25959
rect 26617 25925 26651 25959
rect 16129 25857 16163 25891
rect 19993 25857 20027 25891
rect 20177 25857 20211 25891
rect 22845 25857 22879 25891
rect 23029 25857 23063 25891
rect 23489 25857 23523 25891
rect 23673 25857 23707 25891
rect 25329 25857 25363 25891
rect 25513 25857 25547 25891
rect 26433 25857 26467 25891
rect 27169 25857 27203 25891
rect 27353 25857 27387 25891
rect 1685 25789 1719 25823
rect 2789 25789 2823 25823
rect 16865 25789 16899 25823
rect 25605 25789 25639 25823
rect 26157 25789 26191 25823
rect 23581 25721 23615 25755
rect 27169 25721 27203 25755
rect 26249 25653 26283 25687
rect 1685 25449 1719 25483
rect 17049 25449 17083 25483
rect 18521 25449 18555 25483
rect 25789 25449 25823 25483
rect 21557 25381 21591 25415
rect 15577 25313 15611 25347
rect 25329 25313 25363 25347
rect 25421 25313 25455 25347
rect 26525 25313 26559 25347
rect 15853 25245 15887 25279
rect 18521 25245 18555 25279
rect 18705 25245 18739 25279
rect 21557 25245 21591 25279
rect 21741 25245 21775 25279
rect 21833 25245 21867 25279
rect 24041 25245 24075 25279
rect 25053 25245 25087 25279
rect 25237 25245 25271 25279
rect 25605 25245 25639 25279
rect 16681 25177 16715 25211
rect 16865 25177 16899 25211
rect 26709 25177 26743 25211
rect 28365 25177 28399 25211
rect 15761 25109 15795 25143
rect 16221 25109 16255 25143
rect 22569 25109 22603 25143
rect 20545 24905 20579 24939
rect 25421 24905 25455 24939
rect 27261 24905 27295 24939
rect 20913 24837 20947 24871
rect 1593 24769 1627 24803
rect 17417 24769 17451 24803
rect 17673 24769 17707 24803
rect 19901 24769 19935 24803
rect 21005 24769 21039 24803
rect 22201 24769 22235 24803
rect 22569 24769 22603 24803
rect 22845 24769 22879 24803
rect 23765 24769 23799 24803
rect 23857 24769 23891 24803
rect 24501 24769 24535 24803
rect 25605 24769 25639 24803
rect 25697 24769 25731 24803
rect 25881 24769 25915 24803
rect 27169 24769 27203 24803
rect 27813 24769 27847 24803
rect 20085 24701 20119 24735
rect 21189 24701 21223 24735
rect 22661 24701 22695 24735
rect 24593 24701 24627 24735
rect 24777 24701 24811 24735
rect 25789 24701 25823 24735
rect 18797 24633 18831 24667
rect 24041 24633 24075 24667
rect 1777 24565 1811 24599
rect 19717 24565 19751 24599
rect 24685 24565 24719 24599
rect 17325 24361 17359 24395
rect 21649 24361 21683 24395
rect 23673 24361 23707 24395
rect 24777 24361 24811 24395
rect 28365 24225 28399 24259
rect 17141 24157 17175 24191
rect 17325 24157 17359 24191
rect 19441 24157 19475 24191
rect 22762 24157 22796 24191
rect 23029 24157 23063 24191
rect 24685 24157 24719 24191
rect 24869 24157 24903 24191
rect 26525 24157 26559 24191
rect 19708 24089 19742 24123
rect 23489 24089 23523 24123
rect 23689 24089 23723 24123
rect 26709 24089 26743 24123
rect 20821 24021 20855 24055
rect 23857 24021 23891 24055
rect 19717 23817 19751 23851
rect 20453 23817 20487 23851
rect 20913 23817 20947 23851
rect 27353 23817 27387 23851
rect 17477 23749 17511 23783
rect 17693 23749 17727 23783
rect 20821 23749 20855 23783
rect 18337 23681 18371 23715
rect 18797 23681 18831 23715
rect 18981 23681 19015 23715
rect 19901 23681 19935 23715
rect 27445 23681 27479 23715
rect 27905 23681 27939 23715
rect 21097 23613 21131 23647
rect 17325 23545 17359 23579
rect 17509 23477 17543 23511
rect 18245 23477 18279 23511
rect 18981 23477 19015 23511
rect 26617 23477 26651 23511
rect 17233 23273 17267 23307
rect 17509 23205 17543 23239
rect 18337 23205 18371 23239
rect 23765 23205 23799 23239
rect 17693 23137 17727 23171
rect 19809 23137 19843 23171
rect 20545 23137 20579 23171
rect 25237 23137 25271 23171
rect 26525 23137 26559 23171
rect 28365 23137 28399 23171
rect 15669 23069 15703 23103
rect 15853 23069 15887 23103
rect 16405 23069 16439 23103
rect 16497 23069 16531 23103
rect 17417 23069 17451 23103
rect 17601 23069 17635 23103
rect 17877 23069 17911 23103
rect 18337 23069 18371 23103
rect 18521 23069 18555 23103
rect 19625 23069 19659 23103
rect 20729 23069 20763 23103
rect 23489 23069 23523 23103
rect 25145 23069 25179 23103
rect 16681 23001 16715 23035
rect 23765 23001 23799 23035
rect 26709 23001 26743 23035
rect 15761 22933 15795 22967
rect 19441 22933 19475 22967
rect 20913 22933 20947 22967
rect 23581 22933 23615 22967
rect 25513 22933 25547 22967
rect 18521 22729 18555 22763
rect 20729 22729 20763 22763
rect 21189 22729 21223 22763
rect 26525 22729 26559 22763
rect 27261 22729 27295 22763
rect 21097 22661 21131 22695
rect 17049 22593 17083 22627
rect 17141 22593 17175 22627
rect 17233 22593 17267 22627
rect 17509 22593 17543 22627
rect 18705 22593 18739 22627
rect 18889 22593 18923 22627
rect 18980 22593 19014 22627
rect 19165 22593 19199 22627
rect 19809 22593 19843 22627
rect 22753 22593 22787 22627
rect 22937 22593 22971 22627
rect 23857 22593 23891 22627
rect 24041 22593 24075 22627
rect 24317 22593 24351 22627
rect 25145 22593 25179 22627
rect 25401 22593 25435 22627
rect 27353 22593 27387 22627
rect 17325 22525 17359 22559
rect 21373 22525 21407 22559
rect 24133 22525 24167 22559
rect 18797 22457 18831 22491
rect 23949 22457 23983 22491
rect 16865 22389 16899 22423
rect 19717 22389 19751 22423
rect 22845 22389 22879 22423
rect 23673 22389 23707 22423
rect 28089 22389 28123 22423
rect 19625 22185 19659 22219
rect 25237 22185 25271 22219
rect 23949 22049 23983 22083
rect 27537 22049 27571 22083
rect 28365 22049 28399 22083
rect 16037 21981 16071 22015
rect 16221 21981 16255 22015
rect 20453 21981 20487 22015
rect 22293 21981 22327 22015
rect 22477 21981 22511 22015
rect 22569 21981 22603 22015
rect 23857 21981 23891 22015
rect 24041 21981 24075 22015
rect 24593 21981 24627 22015
rect 24777 21981 24811 22015
rect 24869 21981 24903 22015
rect 24961 21981 24995 22015
rect 19533 21913 19567 21947
rect 20720 21913 20754 21947
rect 28181 21913 28215 21947
rect 16129 21845 16163 21879
rect 21833 21845 21867 21879
rect 22391 21845 22425 21879
rect 18245 21641 18279 21675
rect 20729 21641 20763 21675
rect 22937 21641 22971 21675
rect 27905 21641 27939 21675
rect 17110 21573 17144 21607
rect 19533 21505 19567 21539
rect 20913 21505 20947 21539
rect 22661 21505 22695 21539
rect 23857 21505 23891 21539
rect 24961 21505 24995 21539
rect 25145 21505 25179 21539
rect 25237 21505 25271 21539
rect 25513 21505 25547 21539
rect 27353 21505 27387 21539
rect 27813 21505 27847 21539
rect 16865 21437 16899 21471
rect 22293 21437 22327 21471
rect 22753 21437 22787 21471
rect 23949 21437 23983 21471
rect 24225 21437 24259 21471
rect 25421 21437 25455 21471
rect 19809 21369 19843 21403
rect 24961 21301 24995 21335
rect 27261 21301 27295 21335
rect 20269 21029 20303 21063
rect 20913 20961 20947 20995
rect 23397 20961 23431 20995
rect 26525 20961 26559 20995
rect 28365 20961 28399 20995
rect 16037 20893 16071 20927
rect 18705 20893 18739 20927
rect 19441 20893 19475 20927
rect 19625 20893 19659 20927
rect 19809 20893 19843 20927
rect 23130 20893 23164 20927
rect 26709 20825 26743 20859
rect 16221 20757 16255 20791
rect 18889 20757 18923 20791
rect 20637 20757 20671 20791
rect 20729 20757 20763 20791
rect 22017 20757 22051 20791
rect 15853 20553 15887 20587
rect 27353 20553 27387 20587
rect 19524 20485 19558 20519
rect 25504 20485 25538 20519
rect 1961 20417 1995 20451
rect 15485 20417 15519 20451
rect 15669 20417 15703 20451
rect 16865 20417 16899 20451
rect 17121 20417 17155 20451
rect 19257 20417 19291 20451
rect 27169 20417 27203 20451
rect 25237 20349 25271 20383
rect 26617 20281 26651 20315
rect 1869 20213 1903 20247
rect 18245 20213 18279 20247
rect 20637 20213 20671 20247
rect 27905 20213 27939 20247
rect 15209 20009 15243 20043
rect 1777 19873 1811 19907
rect 2789 19873 2823 19907
rect 15761 19873 15795 19907
rect 26525 19873 26559 19907
rect 28365 19873 28399 19907
rect 1593 19805 1627 19839
rect 15577 19805 15611 19839
rect 21465 19805 21499 19839
rect 21649 19805 21683 19839
rect 21741 19805 21775 19839
rect 21833 19805 21867 19839
rect 24777 19805 24811 19839
rect 25053 19805 25087 19839
rect 25237 19805 25271 19839
rect 26709 19737 26743 19771
rect 15669 19669 15703 19703
rect 22109 19669 22143 19703
rect 24593 19669 24627 19703
rect 16957 19465 16991 19499
rect 18087 19465 18121 19499
rect 18705 19465 18739 19499
rect 22109 19465 22143 19499
rect 25605 19465 25639 19499
rect 27353 19465 27387 19499
rect 16221 19397 16255 19431
rect 17877 19397 17911 19431
rect 23222 19397 23256 19431
rect 1685 19329 1719 19363
rect 16129 19329 16163 19363
rect 16865 19329 16899 19363
rect 17141 19329 17175 19363
rect 18981 19329 19015 19363
rect 19073 19329 19107 19363
rect 19717 19329 19751 19363
rect 20637 19329 20671 19363
rect 20821 19329 20855 19363
rect 21281 19329 21315 19363
rect 21373 19329 21407 19363
rect 23489 19329 23523 19363
rect 24961 19329 24995 19363
rect 25145 19329 25179 19363
rect 25237 19329 25271 19363
rect 25329 19329 25363 19363
rect 27445 19329 27479 19363
rect 18890 19261 18924 19295
rect 19165 19261 19199 19295
rect 19993 19261 20027 19295
rect 20085 19261 20119 19295
rect 27905 19261 27939 19295
rect 17141 19193 17175 19227
rect 19901 19193 19935 19227
rect 20637 19193 20671 19227
rect 18061 19125 18095 19159
rect 18245 19125 18279 19159
rect 19809 19125 19843 19159
rect 19533 18921 19567 18955
rect 27721 18921 27755 18955
rect 17325 18853 17359 18887
rect 23397 18853 23431 18887
rect 22109 18785 22143 18819
rect 22293 18785 22327 18819
rect 23765 18785 23799 18819
rect 26341 18785 26375 18819
rect 1593 18717 1627 18751
rect 17049 18717 17083 18751
rect 17141 18717 17175 18751
rect 17417 18717 17451 18751
rect 18061 18717 18095 18751
rect 18521 18717 18555 18751
rect 18705 18717 18739 18751
rect 19441 18717 19475 18751
rect 19625 18717 19659 18751
rect 24777 18717 24811 18751
rect 28365 18717 28399 18751
rect 20453 18649 20487 18683
rect 24593 18649 24627 18683
rect 26608 18649 26642 18683
rect 1777 18581 1811 18615
rect 16865 18581 16899 18615
rect 17969 18581 18003 18615
rect 18521 18581 18555 18615
rect 23305 18581 23339 18615
rect 16865 18377 16899 18411
rect 17233 18377 17267 18411
rect 21189 18377 21223 18411
rect 24685 18377 24719 18411
rect 27997 18377 28031 18411
rect 19993 18309 20027 18343
rect 23397 18309 23431 18343
rect 15669 18241 15703 18275
rect 15853 18241 15887 18275
rect 17141 18241 17175 18275
rect 17325 18241 17359 18275
rect 17509 18241 17543 18275
rect 20821 18241 20855 18275
rect 21005 18241 21039 18275
rect 22753 18241 22787 18275
rect 22937 18241 22971 18275
rect 27353 18241 27387 18275
rect 27537 18241 27571 18275
rect 28181 18241 28215 18275
rect 17601 18173 17635 18207
rect 18245 18173 18279 18207
rect 27169 18173 27203 18207
rect 1685 18037 1719 18071
rect 16037 18037 16071 18071
rect 22937 18037 22971 18071
rect 15393 17833 15427 17867
rect 17233 17833 17267 17867
rect 17417 17833 17451 17867
rect 18429 17833 18463 17867
rect 19717 17833 19751 17867
rect 1593 17697 1627 17731
rect 2789 17697 2823 17731
rect 15853 17697 15887 17731
rect 15945 17697 15979 17731
rect 16865 17697 16899 17731
rect 24593 17697 24627 17731
rect 26525 17697 26559 17731
rect 28365 17697 28399 17731
rect 18797 17629 18831 17663
rect 19441 17629 19475 17663
rect 22661 17629 22695 17663
rect 23121 17629 23155 17663
rect 23305 17629 23339 17663
rect 23489 17629 23523 17663
rect 24860 17629 24894 17663
rect 1777 17561 1811 17595
rect 17233 17561 17267 17595
rect 19533 17561 19567 17595
rect 19717 17561 19751 17595
rect 28181 17561 28215 17595
rect 15761 17493 15795 17527
rect 18245 17493 18279 17527
rect 18429 17493 18463 17527
rect 22477 17493 22511 17527
rect 25973 17493 26007 17527
rect 1961 17289 1995 17323
rect 17969 17289 18003 17323
rect 19901 17289 19935 17323
rect 27169 17289 27203 17323
rect 27537 17289 27571 17323
rect 16037 17221 16071 17255
rect 25513 17221 25547 17255
rect 2053 17153 2087 17187
rect 15761 17153 15795 17187
rect 16865 17153 16899 17187
rect 17785 17153 17819 17187
rect 17969 17153 18003 17187
rect 18705 17153 18739 17187
rect 18981 17153 19015 17187
rect 19533 17153 19567 17187
rect 19717 17153 19751 17187
rect 22017 17153 22051 17187
rect 22201 17153 22235 17187
rect 22385 17153 22419 17187
rect 22845 17153 22879 17187
rect 23581 17153 23615 17187
rect 23837 17153 23871 17187
rect 25881 17153 25915 17187
rect 26433 17153 26467 17187
rect 18613 17085 18647 17119
rect 19073 17085 19107 17119
rect 27629 17085 27663 17119
rect 27721 17085 27755 17119
rect 18429 17017 18463 17051
rect 17049 16949 17083 16983
rect 23029 16949 23063 16983
rect 24961 16949 24995 16983
rect 26525 16949 26559 16983
rect 13277 16745 13311 16779
rect 18797 16745 18831 16779
rect 27169 16745 27203 16779
rect 27905 16745 27939 16779
rect 16865 16609 16899 16643
rect 21281 16609 21315 16643
rect 23305 16609 23339 16643
rect 25789 16609 25823 16643
rect 2145 16541 2179 16575
rect 13461 16541 13495 16575
rect 13737 16541 13771 16575
rect 17132 16541 17166 16575
rect 18889 16541 18923 16575
rect 19717 16541 19751 16575
rect 21373 16541 21407 16575
rect 23038 16541 23072 16575
rect 23765 16541 23799 16575
rect 23949 16541 23983 16575
rect 24869 16541 24903 16575
rect 25605 16541 25639 16575
rect 27353 16541 27387 16575
rect 27813 16541 27847 16575
rect 23857 16473 23891 16507
rect 2053 16405 2087 16439
rect 13645 16405 13679 16439
rect 18245 16405 18279 16439
rect 19533 16405 19567 16439
rect 20803 16405 20837 16439
rect 21281 16405 21315 16439
rect 21925 16405 21959 16439
rect 24685 16405 24719 16439
rect 25421 16405 25455 16439
rect 14105 16201 14139 16235
rect 20361 16201 20395 16235
rect 22017 16201 22051 16235
rect 22385 16201 22419 16235
rect 24777 16201 24811 16235
rect 1869 16133 1903 16167
rect 14381 16133 14415 16167
rect 16129 16133 16163 16167
rect 25482 16133 25516 16167
rect 14105 16065 14139 16099
rect 14197 16065 14231 16099
rect 15761 16065 15795 16099
rect 15945 16065 15979 16099
rect 20453 16065 20487 16099
rect 24593 16065 24627 16099
rect 27445 16065 27479 16099
rect 1685 15997 1719 16031
rect 2789 15997 2823 16031
rect 20637 15997 20671 16031
rect 22477 15997 22511 16031
rect 22569 15997 22603 16031
rect 25237 15997 25271 16031
rect 19993 15861 20027 15895
rect 26617 15861 26651 15895
rect 27537 15861 27571 15895
rect 28273 15861 28307 15895
rect 1685 15657 1719 15691
rect 13737 15657 13771 15691
rect 15761 15657 15795 15691
rect 25329 15657 25363 15691
rect 21373 15589 21407 15623
rect 20637 15521 20671 15555
rect 25881 15521 25915 15555
rect 27537 15521 27571 15555
rect 28181 15521 28215 15555
rect 28365 15521 28399 15555
rect 13553 15453 13587 15487
rect 13737 15453 13771 15487
rect 14473 15453 14507 15487
rect 14657 15453 14691 15487
rect 16037 15453 16071 15487
rect 20729 15453 20763 15487
rect 21649 15453 21683 15487
rect 25697 15453 25731 15487
rect 14565 15385 14599 15419
rect 21925 15385 21959 15419
rect 15577 15317 15611 15351
rect 20159 15317 20193 15351
rect 20637 15317 20671 15351
rect 21833 15317 21867 15351
rect 25789 15317 25823 15351
rect 13645 15113 13679 15147
rect 14381 15113 14415 15147
rect 15025 15113 15059 15147
rect 15669 15113 15703 15147
rect 16313 15113 16347 15147
rect 2053 14977 2087 15011
rect 13461 14977 13495 15011
rect 14197 14977 14231 15011
rect 14473 14977 14507 15011
rect 14933 14977 14967 15011
rect 15209 14977 15243 15011
rect 17049 14977 17083 15011
rect 19340 14977 19374 15011
rect 23590 14977 23624 15011
rect 23857 14977 23891 15011
rect 27445 14977 27479 15011
rect 13277 14909 13311 14943
rect 15853 14909 15887 14943
rect 15945 14909 15979 14943
rect 19073 14909 19107 14943
rect 15209 14841 15243 14875
rect 1961 14773 1995 14807
rect 14197 14773 14231 14807
rect 16957 14773 16991 14807
rect 20453 14773 20487 14807
rect 22477 14773 22511 14807
rect 27353 14773 27387 14807
rect 27905 14773 27939 14807
rect 14289 14569 14323 14603
rect 15945 14569 15979 14603
rect 20821 14569 20855 14603
rect 12449 14501 12483 14535
rect 18245 14501 18279 14535
rect 1777 14433 1811 14467
rect 2789 14433 2823 14467
rect 9689 14433 9723 14467
rect 11437 14433 11471 14467
rect 12909 14433 12943 14467
rect 24593 14433 24627 14467
rect 26525 14433 26559 14467
rect 26709 14433 26743 14467
rect 1593 14365 1627 14399
rect 8401 14365 8435 14399
rect 12265 14365 12299 14399
rect 12449 14365 12483 14399
rect 13185 14365 13219 14399
rect 13369 14365 13403 14399
rect 14427 14365 14461 14399
rect 14565 14365 14599 14399
rect 14840 14365 14874 14399
rect 14933 14365 14967 14399
rect 15485 14365 15519 14399
rect 15577 14365 15611 14399
rect 15761 14365 15795 14399
rect 16865 14365 16899 14399
rect 18889 14365 18923 14399
rect 19441 14365 19475 14399
rect 21281 14365 21315 14399
rect 28365 14365 28399 14399
rect 11253 14297 11287 14331
rect 14657 14297 14691 14331
rect 17110 14297 17144 14331
rect 19708 14297 19742 14331
rect 21548 14297 21582 14331
rect 24838 14297 24872 14331
rect 8493 14229 8527 14263
rect 13093 14229 13127 14263
rect 18705 14229 18739 14263
rect 22661 14229 22695 14263
rect 25973 14229 26007 14263
rect 15301 14025 15335 14059
rect 16313 14025 16347 14059
rect 17233 14025 17267 14059
rect 19625 14025 19659 14059
rect 28181 14025 28215 14059
rect 9965 13957 9999 13991
rect 11069 13957 11103 13991
rect 13369 13957 13403 13991
rect 15485 13957 15519 13991
rect 15669 13957 15703 13991
rect 22262 13957 22296 13991
rect 1685 13889 1719 13923
rect 10149 13889 10183 13923
rect 10977 13889 11011 13923
rect 14749 13889 14783 13923
rect 16129 13889 16163 13923
rect 17325 13889 17359 13923
rect 18245 13889 18279 13923
rect 18512 13889 18546 13923
rect 22017 13889 22051 13923
rect 24225 13889 24259 13923
rect 24492 13889 24526 13923
rect 27353 13889 27387 13923
rect 28365 13889 28399 13923
rect 2513 13821 2547 13855
rect 8309 13821 8343 13855
rect 11713 13821 11747 13855
rect 13553 13821 13587 13855
rect 14289 13821 14323 13855
rect 14473 13821 14507 13855
rect 14565 13821 14599 13855
rect 14657 13821 14691 13855
rect 17417 13821 17451 13855
rect 16865 13685 16899 13719
rect 23397 13685 23431 13719
rect 25605 13685 25639 13719
rect 27261 13685 27295 13719
rect 9781 13481 9815 13515
rect 14381 13481 14415 13515
rect 16589 13481 16623 13515
rect 1593 13345 1627 13379
rect 3433 13345 3467 13379
rect 16957 13345 16991 13379
rect 26709 13345 26743 13379
rect 28089 13345 28123 13379
rect 9689 13277 9723 13311
rect 14289 13277 14323 13311
rect 14473 13277 14507 13311
rect 14933 13277 14967 13311
rect 15117 13277 15151 13311
rect 16773 13277 16807 13311
rect 26525 13277 26559 13311
rect 3249 13209 3283 13243
rect 15025 13209 15059 13243
rect 2053 12937 2087 12971
rect 19441 12937 19475 12971
rect 24777 12937 24811 12971
rect 2145 12801 2179 12835
rect 19625 12801 19659 12835
rect 22569 12801 22603 12835
rect 22753 12801 22787 12835
rect 24133 12801 24167 12835
rect 24317 12801 24351 12835
rect 24409 12801 24443 12835
rect 24501 12801 24535 12835
rect 27445 12801 27479 12835
rect 27905 12665 27939 12699
rect 22753 12597 22787 12631
rect 27353 12597 27387 12631
rect 19625 12393 19659 12427
rect 21557 12393 21591 12427
rect 24593 12393 24627 12427
rect 25697 12393 25731 12427
rect 21005 12257 21039 12291
rect 23489 12257 23523 12291
rect 23581 12257 23615 12291
rect 26525 12257 26559 12291
rect 26709 12257 26743 12291
rect 28365 12257 28399 12291
rect 19441 12189 19475 12223
rect 20729 12189 20763 12223
rect 21741 12189 21775 12223
rect 22385 12189 22419 12223
rect 22477 12189 22511 12223
rect 22845 12189 22879 12223
rect 23673 12189 23707 12223
rect 23765 12189 23799 12223
rect 24869 12189 24903 12223
rect 24961 12189 24995 12223
rect 25053 12189 25087 12223
rect 25237 12189 25271 12223
rect 25973 12189 26007 12223
rect 25697 12121 25731 12155
rect 25881 12121 25915 12155
rect 20361 12053 20395 12087
rect 20821 12053 20855 12087
rect 22201 12053 22235 12087
rect 22569 12053 22603 12087
rect 22753 12053 22787 12087
rect 23305 12053 23339 12087
rect 19441 11849 19475 11883
rect 20821 11849 20855 11883
rect 22017 11849 22051 11883
rect 23121 11849 23155 11883
rect 24225 11849 24259 11883
rect 25329 11849 25363 11883
rect 19625 11713 19659 11747
rect 22293 11713 22327 11747
rect 22385 11713 22419 11747
rect 22477 11713 22511 11747
rect 22661 11713 22695 11747
rect 23397 11713 23431 11747
rect 23489 11713 23523 11747
rect 23581 11713 23615 11747
rect 23765 11713 23799 11747
rect 24501 11713 24535 11747
rect 24593 11713 24627 11747
rect 25421 11713 25455 11747
rect 1685 11645 1719 11679
rect 1869 11645 1903 11679
rect 2789 11645 2823 11679
rect 19809 11645 19843 11679
rect 20913 11645 20947 11679
rect 21005 11645 21039 11679
rect 24409 11645 24443 11679
rect 24685 11645 24719 11679
rect 20453 11509 20487 11543
rect 1685 11305 1719 11339
rect 2421 11305 2455 11339
rect 19533 11305 19567 11339
rect 22385 11305 22419 11339
rect 23581 11305 23615 11339
rect 25145 11305 25179 11339
rect 21649 11169 21683 11203
rect 23305 11169 23339 11203
rect 23397 11169 23431 11203
rect 24685 11169 24719 11203
rect 24777 11169 24811 11203
rect 27537 11169 27571 11203
rect 2513 11101 2547 11135
rect 19717 11101 19751 11135
rect 19901 11101 19935 11135
rect 21557 11101 21591 11135
rect 22293 11101 22327 11135
rect 22937 11101 22971 11135
rect 24869 11101 24903 11135
rect 24961 11101 24995 11135
rect 28365 11101 28399 11135
rect 21465 11033 21499 11067
rect 23029 11033 23063 11067
rect 28181 11033 28215 11067
rect 21097 10965 21131 10999
rect 23213 10965 23247 10999
rect 21097 10761 21131 10795
rect 22753 10761 22787 10795
rect 22385 10693 22419 10727
rect 22601 10693 22635 10727
rect 20729 10625 20763 10659
rect 20913 10625 20947 10659
rect 26433 10625 26467 10659
rect 28089 10625 28123 10659
rect 22569 10421 22603 10455
rect 26525 10421 26559 10455
rect 27169 10421 27203 10455
rect 26525 10081 26559 10115
rect 26709 10081 26743 10115
rect 28365 10081 28399 10115
rect 1777 10013 1811 10047
rect 3065 10013 3099 10047
rect 27721 9605 27755 9639
rect 2513 9537 2547 9571
rect 3065 9537 3099 9571
rect 25973 9537 26007 9571
rect 27629 9537 27663 9571
rect 3249 9469 3283 9503
rect 4169 9469 4203 9503
rect 1685 9333 1719 9367
rect 2421 9333 2455 9367
rect 25881 9333 25915 9367
rect 4077 9129 4111 9163
rect 1593 8993 1627 9027
rect 1777 8993 1811 9027
rect 2789 8993 2823 9027
rect 25605 8993 25639 9027
rect 25789 8993 25823 9027
rect 4169 8925 4203 8959
rect 28089 8925 28123 8959
rect 27445 8857 27479 8891
rect 1685 8449 1719 8483
rect 4813 8449 4847 8483
rect 9321 8449 9355 8483
rect 27721 8449 27755 8483
rect 1869 8381 1903 8415
rect 2789 8381 2823 8415
rect 9413 8313 9447 8347
rect 3985 8245 4019 8279
rect 4721 8245 4755 8279
rect 26617 8245 26651 8279
rect 27813 8245 27847 8279
rect 2145 8041 2179 8075
rect 3985 7905 4019 7939
rect 4169 7905 4203 7939
rect 5549 7905 5583 7939
rect 27537 7905 27571 7939
rect 28181 7905 28215 7939
rect 28365 7905 28399 7939
rect 2237 7837 2271 7871
rect 2237 7361 2271 7395
rect 26617 7361 26651 7395
rect 27629 7361 27663 7395
rect 26157 7293 26191 7327
rect 26433 7293 26467 7327
rect 27721 7293 27755 7327
rect 2145 7157 2179 7191
rect 3065 7157 3099 7191
rect 1777 6817 1811 6851
rect 2789 6817 2823 6851
rect 24593 6817 24627 6851
rect 25145 6817 25179 6851
rect 1593 6749 1627 6783
rect 23857 6749 23891 6783
rect 27629 6749 27663 6783
rect 23949 6681 23983 6715
rect 24777 6681 24811 6715
rect 26433 6341 26467 6375
rect 27537 6341 27571 6375
rect 1685 6273 1719 6307
rect 2329 6273 2363 6307
rect 2973 6273 3007 6307
rect 26617 6273 26651 6307
rect 27445 6273 27479 6307
rect 2421 6205 2455 6239
rect 3157 6205 3191 6239
rect 4169 6205 4203 6239
rect 26157 6205 26191 6239
rect 3065 5729 3099 5763
rect 25881 5729 25915 5763
rect 1593 5661 1627 5695
rect 4721 5661 4755 5695
rect 25329 5661 25363 5695
rect 26433 5661 26467 5695
rect 1777 5593 1811 5627
rect 26617 5593 26651 5627
rect 28273 5593 28307 5627
rect 2421 5321 2455 5355
rect 26433 5321 26467 5355
rect 1685 5185 1719 5219
rect 2513 5185 2547 5219
rect 5365 5185 5399 5219
rect 26341 5185 26375 5219
rect 27169 5185 27203 5219
rect 2973 5117 3007 5151
rect 3157 5117 3191 5151
rect 4813 5117 4847 5151
rect 5457 4981 5491 5015
rect 27905 4981 27939 5015
rect 2973 4777 3007 4811
rect 5457 4641 5491 4675
rect 5825 4641 5859 4675
rect 23949 4641 23983 4675
rect 27445 4641 27479 4675
rect 1593 4573 1627 4607
rect 2421 4573 2455 4607
rect 3985 4573 4019 4607
rect 4813 4573 4847 4607
rect 5273 4573 5307 4607
rect 28365 4573 28399 4607
rect 22109 4505 22143 4539
rect 23765 4505 23799 4539
rect 28181 4505 28215 4539
rect 2329 4437 2363 4471
rect 27813 4233 27847 4267
rect 1961 4097 1995 4131
rect 2421 4097 2455 4131
rect 2513 4097 2547 4131
rect 3249 4097 3283 4131
rect 3709 4097 3743 4131
rect 6745 4097 6779 4131
rect 10517 4097 10551 4131
rect 18705 4097 18739 4131
rect 21281 4097 21315 4131
rect 22201 4097 22235 4131
rect 22293 4097 22327 4131
rect 27721 4097 27755 4131
rect 3893 4029 3927 4063
rect 4353 4029 4387 4063
rect 12817 4029 12851 4063
rect 13001 4029 13035 4063
rect 13645 4029 13679 4063
rect 1869 3893 1903 3927
rect 3157 3893 3191 3927
rect 6653 3893 6687 3927
rect 7757 3893 7791 3927
rect 10609 3893 10643 3927
rect 18797 3893 18831 3927
rect 20453 3893 20487 3927
rect 21189 3893 21223 3927
rect 4261 3689 4295 3723
rect 12909 3689 12943 3723
rect 1593 3553 1627 3587
rect 1777 3553 1811 3587
rect 2053 3553 2087 3587
rect 5917 3553 5951 3587
rect 6469 3553 6503 3587
rect 10609 3553 10643 3587
rect 10977 3553 11011 3587
rect 20361 3553 20395 3587
rect 20545 3553 20579 3587
rect 21281 3553 21315 3587
rect 27537 3553 27571 3587
rect 4353 3485 4387 3519
rect 5273 3485 5307 3519
rect 5733 3485 5767 3519
rect 8217 3485 8251 3519
rect 9321 3485 9355 3519
rect 9965 3485 9999 3519
rect 10425 3485 10459 3519
rect 13553 3485 13587 3519
rect 14289 3485 14323 3519
rect 16221 3485 16255 3519
rect 16681 3485 16715 3519
rect 17693 3485 17727 3519
rect 18153 3485 18187 3519
rect 19441 3485 19475 3519
rect 26065 3485 26099 3519
rect 26525 3485 26559 3519
rect 26709 3417 26743 3451
rect 8125 3349 8159 3383
rect 13645 3349 13679 3383
rect 16773 3349 16807 3383
rect 18245 3349 18279 3383
rect 12909 3145 12943 3179
rect 27261 3145 27295 3179
rect 1961 3077 1995 3111
rect 4353 3077 4387 3111
rect 7113 3077 7147 3111
rect 9413 3077 9447 3111
rect 14197 3077 14231 3111
rect 17049 3077 17083 3111
rect 19349 3077 19383 3111
rect 26433 3077 26467 3111
rect 4169 3009 4203 3043
rect 9229 3009 9263 3043
rect 12817 3009 12851 3043
rect 14013 3009 14047 3043
rect 16865 3009 16899 3043
rect 19165 3009 19199 3043
rect 26617 3009 26651 3043
rect 27353 3009 27387 3043
rect 28089 3009 28123 3043
rect 1777 2941 1811 2975
rect 2789 2941 2823 2975
rect 4813 2941 4847 2975
rect 6929 2941 6963 2975
rect 8401 2941 8435 2975
rect 9689 2941 9723 2975
rect 14749 2941 14783 2975
rect 17325 2941 17359 2975
rect 19625 2941 19659 2975
rect 26157 2941 26191 2975
rect 1869 2601 1903 2635
rect 17601 2601 17635 2635
rect 26433 2601 26467 2635
rect 27813 2601 27847 2635
rect 16865 2533 16899 2567
rect 4445 2465 4479 2499
rect 9413 2465 9447 2499
rect 19441 2465 19475 2499
rect 19625 2465 19659 2499
rect 19993 2465 20027 2499
rect 2605 2397 2639 2431
rect 3433 2397 3467 2431
rect 3985 2397 4019 2431
rect 9137 2397 9171 2431
rect 17785 2397 17819 2431
rect 26617 2397 26651 2431
rect 27721 2397 27755 2431
rect 2697 2329 2731 2363
rect 4169 2329 4203 2363
rect 17049 2329 17083 2363
<< metal1 >>
rect 1104 47354 28888 47376
rect 1104 47302 4423 47354
rect 4475 47302 4487 47354
rect 4539 47302 4551 47354
rect 4603 47302 4615 47354
rect 4667 47302 4679 47354
rect 4731 47302 11369 47354
rect 11421 47302 11433 47354
rect 11485 47302 11497 47354
rect 11549 47302 11561 47354
rect 11613 47302 11625 47354
rect 11677 47302 18315 47354
rect 18367 47302 18379 47354
rect 18431 47302 18443 47354
rect 18495 47302 18507 47354
rect 18559 47302 18571 47354
rect 18623 47302 25261 47354
rect 25313 47302 25325 47354
rect 25377 47302 25389 47354
rect 25441 47302 25453 47354
rect 25505 47302 25517 47354
rect 25569 47302 28888 47354
rect 1104 47280 28888 47302
rect 23750 47132 23756 47184
rect 23808 47172 23814 47184
rect 23845 47175 23903 47181
rect 23845 47172 23857 47175
rect 23808 47144 23857 47172
rect 23808 47132 23814 47144
rect 23845 47141 23857 47144
rect 23891 47141 23903 47175
rect 23845 47135 23903 47141
rect 25038 47132 25044 47184
rect 25096 47172 25102 47184
rect 27341 47175 27399 47181
rect 27341 47172 27353 47175
rect 25096 47144 27353 47172
rect 25096 47132 25102 47144
rect 27341 47141 27353 47144
rect 27387 47141 27399 47175
rect 27341 47135 27399 47141
rect 10318 47104 10324 47116
rect 10279 47076 10324 47104
rect 10318 47064 10324 47076
rect 10376 47064 10382 47116
rect 26145 47107 26203 47113
rect 26145 47073 26157 47107
rect 26191 47104 26203 47107
rect 28350 47104 28356 47116
rect 26191 47076 28356 47104
rect 26191 47073 26203 47076
rect 26145 47067 26203 47073
rect 28350 47064 28356 47076
rect 28408 47064 28414 47116
rect 2222 47036 2228 47048
rect 2183 47008 2228 47036
rect 2222 46996 2228 47008
rect 2280 46996 2286 47048
rect 2866 47036 2872 47048
rect 2779 47008 2872 47036
rect 2866 46996 2872 47008
rect 2924 47036 2930 47048
rect 5810 47036 5816 47048
rect 2924 47008 4200 47036
rect 5771 47008 5816 47036
rect 2924 46996 2930 47008
rect 4172 46968 4200 47008
rect 5810 46996 5816 47008
rect 5868 46996 5874 47048
rect 6454 46996 6460 47048
rect 6512 47036 6518 47048
rect 6549 47039 6607 47045
rect 6549 47036 6561 47039
rect 6512 47008 6561 47036
rect 6512 46996 6518 47008
rect 6549 47005 6561 47008
rect 6595 47005 6607 47039
rect 6549 46999 6607 47005
rect 7006 46996 7012 47048
rect 7064 47036 7070 47048
rect 7929 47039 7987 47045
rect 7929 47036 7941 47039
rect 7064 47008 7941 47036
rect 7064 46996 7070 47008
rect 7929 47005 7941 47008
rect 7975 47005 7987 47039
rect 9306 47036 9312 47048
rect 9267 47008 9312 47036
rect 7929 46999 7987 47005
rect 9306 46996 9312 47008
rect 9364 46996 9370 47048
rect 12894 46996 12900 47048
rect 12952 47036 12958 47048
rect 12989 47039 13047 47045
rect 12989 47036 13001 47039
rect 12952 47008 13001 47036
rect 12952 46996 12958 47008
rect 12989 47005 13001 47008
rect 13035 47005 13047 47039
rect 12989 46999 13047 47005
rect 18230 46996 18236 47048
rect 18288 47036 18294 47048
rect 18325 47039 18383 47045
rect 18325 47036 18337 47039
rect 18288 47008 18337 47036
rect 18288 46996 18294 47008
rect 18325 47005 18337 47008
rect 18371 47005 18383 47039
rect 18325 46999 18383 47005
rect 22830 46996 22836 47048
rect 22888 47036 22894 47048
rect 22925 47039 22983 47045
rect 22925 47036 22937 47039
rect 22888 47008 22937 47036
rect 22888 46996 22894 47008
rect 22925 47005 22937 47008
rect 22971 47005 22983 47039
rect 24026 47036 24032 47048
rect 23987 47008 24032 47036
rect 22925 46999 22983 47005
rect 24026 46996 24032 47008
rect 24084 46996 24090 47048
rect 26602 46996 26608 47048
rect 26660 47036 26666 47048
rect 26660 47008 26705 47036
rect 26660 46996 26666 47008
rect 27338 46996 27344 47048
rect 27396 47036 27402 47048
rect 27433 47039 27491 47045
rect 27433 47036 27445 47039
rect 27396 47008 27445 47036
rect 27396 46996 27402 47008
rect 27433 47005 27445 47008
rect 27479 47005 27491 47039
rect 27890 47036 27896 47048
rect 27851 47008 27896 47036
rect 27433 46999 27491 47005
rect 27890 46996 27896 47008
rect 27948 46996 27954 47048
rect 9214 46968 9220 46980
rect 4172 46940 9220 46968
rect 9214 46928 9220 46940
rect 9272 46928 9278 46980
rect 9490 46968 9496 46980
rect 9451 46940 9496 46968
rect 9490 46928 9496 46940
rect 9548 46928 9554 46980
rect 26418 46968 26424 46980
rect 26379 46940 26424 46968
rect 26418 46928 26424 46940
rect 26476 46928 26482 46980
rect 2774 46900 2780 46912
rect 2735 46872 2780 46900
rect 2774 46860 2780 46872
rect 2832 46860 2838 46912
rect 5994 46900 6000 46912
rect 5955 46872 6000 46900
rect 5994 46860 6000 46872
rect 6052 46860 6058 46912
rect 6730 46900 6736 46912
rect 6691 46872 6736 46900
rect 6730 46860 6736 46872
rect 6788 46860 6794 46912
rect 19978 46860 19984 46912
rect 20036 46900 20042 46912
rect 23474 46900 23480 46912
rect 20036 46872 23480 46900
rect 20036 46860 20042 46872
rect 23474 46860 23480 46872
rect 23532 46860 23538 46912
rect 1104 46810 29048 46832
rect 1104 46758 7896 46810
rect 7948 46758 7960 46810
rect 8012 46758 8024 46810
rect 8076 46758 8088 46810
rect 8140 46758 8152 46810
rect 8204 46758 14842 46810
rect 14894 46758 14906 46810
rect 14958 46758 14970 46810
rect 15022 46758 15034 46810
rect 15086 46758 15098 46810
rect 15150 46758 21788 46810
rect 21840 46758 21852 46810
rect 21904 46758 21916 46810
rect 21968 46758 21980 46810
rect 22032 46758 22044 46810
rect 22096 46758 28734 46810
rect 28786 46758 28798 46810
rect 28850 46758 28862 46810
rect 28914 46758 28926 46810
rect 28978 46758 28990 46810
rect 29042 46758 29048 46810
rect 1104 46736 29048 46758
rect 26418 46696 26424 46708
rect 26379 46668 26424 46696
rect 26418 46656 26424 46668
rect 26476 46656 26482 46708
rect 2501 46631 2559 46637
rect 2501 46597 2513 46631
rect 2547 46628 2559 46631
rect 2774 46628 2780 46640
rect 2547 46600 2780 46628
rect 2547 46597 2559 46600
rect 2501 46591 2559 46597
rect 2774 46588 2780 46600
rect 2832 46588 2838 46640
rect 2222 46520 2228 46572
rect 2280 46560 2286 46572
rect 2317 46563 2375 46569
rect 2317 46560 2329 46563
rect 2280 46532 2329 46560
rect 2280 46520 2286 46532
rect 2317 46529 2329 46532
rect 2363 46529 2375 46563
rect 7006 46560 7012 46572
rect 6967 46532 7012 46560
rect 2317 46523 2375 46529
rect 7006 46520 7012 46532
rect 7064 46520 7070 46572
rect 12894 46560 12900 46572
rect 12855 46532 12900 46560
rect 12894 46520 12900 46532
rect 12952 46520 12958 46572
rect 15838 46560 15844 46572
rect 15799 46532 15844 46560
rect 15838 46520 15844 46532
rect 15896 46520 15902 46572
rect 18230 46560 18236 46572
rect 18191 46532 18236 46560
rect 18230 46520 18236 46532
rect 18288 46520 18294 46572
rect 22830 46560 22836 46572
rect 22791 46532 22836 46560
rect 22830 46520 22836 46532
rect 22888 46520 22894 46572
rect 26513 46563 26571 46569
rect 26513 46529 26525 46563
rect 26559 46560 26571 46563
rect 26559 46532 26740 46560
rect 26559 46529 26571 46532
rect 26513 46523 26571 46529
rect 1946 46452 1952 46504
rect 2004 46492 2010 46504
rect 2777 46495 2835 46501
rect 2777 46492 2789 46495
rect 2004 46464 2789 46492
rect 2004 46452 2010 46464
rect 2777 46461 2789 46464
rect 2823 46461 2835 46495
rect 2777 46455 2835 46461
rect 7193 46495 7251 46501
rect 7193 46461 7205 46495
rect 7239 46492 7251 46495
rect 7926 46492 7932 46504
rect 7239 46464 7932 46492
rect 7239 46461 7251 46464
rect 7193 46455 7251 46461
rect 7926 46452 7932 46464
rect 7984 46452 7990 46504
rect 8386 46492 8392 46504
rect 8347 46464 8392 46492
rect 8386 46452 8392 46464
rect 8444 46452 8450 46504
rect 9309 46495 9367 46501
rect 9309 46461 9321 46495
rect 9355 46461 9367 46495
rect 9309 46455 9367 46461
rect 9493 46495 9551 46501
rect 9493 46461 9505 46495
rect 9539 46492 9551 46495
rect 10134 46492 10140 46504
rect 9539 46464 10140 46492
rect 9539 46461 9551 46464
rect 9493 46455 9551 46461
rect 9324 46424 9352 46455
rect 10134 46452 10140 46464
rect 10192 46452 10198 46504
rect 10962 46492 10968 46504
rect 10923 46464 10968 46492
rect 10962 46452 10968 46464
rect 11020 46452 11026 46504
rect 13078 46492 13084 46504
rect 13039 46464 13084 46492
rect 13078 46452 13084 46464
rect 13136 46452 13142 46504
rect 13538 46492 13544 46504
rect 13499 46464 13544 46492
rect 13538 46452 13544 46464
rect 13596 46452 13602 46504
rect 15930 46452 15936 46504
rect 15988 46492 15994 46504
rect 16853 46495 16911 46501
rect 16853 46492 16865 46495
rect 15988 46464 16865 46492
rect 15988 46452 15994 46464
rect 16853 46461 16865 46464
rect 16899 46461 16911 46495
rect 16853 46455 16911 46461
rect 18138 46452 18144 46504
rect 18196 46492 18202 46504
rect 18417 46495 18475 46501
rect 18417 46492 18429 46495
rect 18196 46464 18429 46492
rect 18196 46452 18202 46464
rect 18417 46461 18429 46464
rect 18463 46461 18475 46495
rect 18690 46492 18696 46504
rect 18651 46464 18696 46492
rect 18417 46455 18475 46461
rect 18690 46452 18696 46464
rect 18748 46452 18754 46504
rect 23017 46495 23075 46501
rect 23017 46461 23029 46495
rect 23063 46492 23075 46495
rect 23106 46492 23112 46504
rect 23063 46464 23112 46492
rect 23063 46461 23075 46464
rect 23017 46455 23075 46461
rect 23106 46452 23112 46464
rect 23164 46452 23170 46504
rect 23198 46452 23204 46504
rect 23256 46492 23262 46504
rect 23477 46495 23535 46501
rect 23477 46492 23489 46495
rect 23256 46464 23489 46492
rect 23256 46452 23262 46464
rect 23477 46461 23489 46464
rect 23523 46461 23535 46495
rect 23477 46455 23535 46461
rect 25869 46495 25927 46501
rect 25869 46461 25881 46495
rect 25915 46492 25927 46495
rect 26602 46492 26608 46504
rect 25915 46464 26608 46492
rect 25915 46461 25927 46464
rect 25869 46455 25927 46461
rect 26602 46452 26608 46464
rect 26660 46452 26666 46504
rect 10410 46424 10416 46436
rect 9324 46396 10416 46424
rect 10410 46384 10416 46396
rect 10468 46384 10474 46436
rect 17218 46384 17224 46436
rect 17276 46424 17282 46436
rect 26712 46424 26740 46532
rect 27430 46520 27436 46572
rect 27488 46560 27494 46572
rect 27801 46563 27859 46569
rect 27801 46560 27813 46563
rect 27488 46532 27813 46560
rect 27488 46520 27494 46532
rect 27801 46529 27813 46532
rect 27847 46529 27859 46563
rect 27801 46523 27859 46529
rect 28534 46424 28540 46436
rect 17276 46396 28540 46424
rect 17276 46384 17282 46396
rect 28534 46384 28540 46396
rect 28592 46384 28598 46436
rect 1670 46356 1676 46368
rect 1631 46328 1676 46356
rect 1670 46316 1676 46328
rect 1728 46316 1734 46368
rect 11698 46356 11704 46368
rect 11659 46328 11704 46356
rect 11698 46316 11704 46328
rect 11756 46316 11762 46368
rect 15933 46359 15991 46365
rect 15933 46325 15945 46359
rect 15979 46356 15991 46359
rect 16114 46356 16120 46368
rect 15979 46328 16120 46356
rect 15979 46325 15991 46328
rect 15933 46319 15991 46325
rect 16114 46316 16120 46328
rect 16172 46316 16178 46368
rect 20254 46316 20260 46368
rect 20312 46356 20318 46368
rect 20533 46359 20591 46365
rect 20533 46356 20545 46359
rect 20312 46328 20545 46356
rect 20312 46316 20318 46328
rect 20533 46325 20545 46328
rect 20579 46325 20591 46359
rect 20533 46319 20591 46325
rect 26510 46316 26516 46368
rect 26568 46356 26574 46368
rect 27157 46359 27215 46365
rect 27157 46356 27169 46359
rect 26568 46328 27169 46356
rect 26568 46316 26574 46328
rect 27157 46325 27169 46328
rect 27203 46325 27215 46359
rect 27157 46319 27215 46325
rect 27246 46316 27252 46368
rect 27304 46356 27310 46368
rect 27893 46359 27951 46365
rect 27893 46356 27905 46359
rect 27304 46328 27905 46356
rect 27304 46316 27310 46328
rect 27893 46325 27905 46328
rect 27939 46325 27951 46359
rect 27893 46319 27951 46325
rect 1104 46266 28888 46288
rect 1104 46214 4423 46266
rect 4475 46214 4487 46266
rect 4539 46214 4551 46266
rect 4603 46214 4615 46266
rect 4667 46214 4679 46266
rect 4731 46214 11369 46266
rect 11421 46214 11433 46266
rect 11485 46214 11497 46266
rect 11549 46214 11561 46266
rect 11613 46214 11625 46266
rect 11677 46214 18315 46266
rect 18367 46214 18379 46266
rect 18431 46214 18443 46266
rect 18495 46214 18507 46266
rect 18559 46214 18571 46266
rect 18623 46214 25261 46266
rect 25313 46214 25325 46266
rect 25377 46214 25389 46266
rect 25441 46214 25453 46266
rect 25505 46214 25517 46266
rect 25569 46214 28888 46266
rect 1104 46192 28888 46214
rect 7926 46152 7932 46164
rect 7887 46124 7932 46152
rect 7926 46112 7932 46124
rect 7984 46112 7990 46164
rect 9490 46152 9496 46164
rect 9451 46124 9496 46152
rect 9490 46112 9496 46124
rect 9548 46112 9554 46164
rect 10134 46152 10140 46164
rect 10095 46124 10140 46152
rect 10134 46112 10140 46124
rect 10192 46112 10198 46164
rect 17218 46152 17224 46164
rect 10244 46124 17224 46152
rect 1026 45976 1032 46028
rect 1084 46016 1090 46028
rect 1581 46019 1639 46025
rect 1581 46016 1593 46019
rect 1084 45988 1593 46016
rect 1084 45976 1090 45988
rect 1581 45985 1593 45988
rect 1627 45985 1639 46019
rect 1581 45979 1639 45985
rect 2590 45976 2596 46028
rect 2648 46016 2654 46028
rect 4433 46019 4491 46025
rect 4433 46016 4445 46019
rect 2648 45988 4445 46016
rect 2648 45976 2654 45988
rect 4433 45985 4445 45988
rect 4479 45985 4491 46019
rect 10244 46016 10272 46124
rect 17218 46112 17224 46124
rect 17276 46112 17282 46164
rect 18138 46112 18144 46164
rect 18196 46152 18202 46164
rect 18417 46155 18475 46161
rect 18417 46152 18429 46155
rect 18196 46124 18429 46152
rect 18196 46112 18202 46124
rect 18417 46121 18429 46124
rect 18463 46121 18475 46155
rect 23106 46152 23112 46164
rect 23067 46124 23112 46152
rect 18417 46115 18475 46121
rect 23106 46112 23112 46124
rect 23164 46112 23170 46164
rect 27430 46084 27436 46096
rect 4433 45979 4491 45985
rect 8036 45988 10272 46016
rect 10704 46056 27436 46084
rect 3418 45908 3424 45960
rect 3476 45948 3482 45960
rect 3970 45948 3976 45960
rect 3476 45920 3521 45948
rect 3931 45920 3976 45948
rect 3476 45908 3482 45920
rect 3970 45908 3976 45920
rect 4028 45908 4034 45960
rect 7742 45908 7748 45960
rect 7800 45948 7806 45960
rect 8036 45957 8064 45988
rect 10704 45960 10732 46056
rect 11333 46019 11391 46025
rect 11333 45985 11345 46019
rect 11379 46016 11391 46019
rect 11698 46016 11704 46028
rect 11379 45988 11704 46016
rect 11379 45985 11391 45988
rect 11333 45979 11391 45985
rect 11698 45976 11704 45988
rect 11756 45976 11762 46028
rect 11790 45976 11796 46028
rect 11848 46016 11854 46028
rect 15930 46016 15936 46028
rect 11848 45988 11893 46016
rect 15891 45988 15936 46016
rect 11848 45976 11854 45988
rect 15930 45976 15936 45988
rect 15988 45976 15994 46028
rect 16114 46016 16120 46028
rect 16075 45988 16120 46016
rect 16114 45976 16120 45988
rect 16172 45976 16178 46028
rect 16758 46016 16764 46028
rect 16719 45988 16764 46016
rect 16758 45976 16764 45988
rect 16816 45976 16822 46028
rect 20254 46016 20260 46028
rect 20215 45988 20260 46016
rect 20254 45976 20260 45988
rect 20312 45976 20318 46028
rect 21266 46016 21272 46028
rect 21227 45988 21272 46016
rect 21266 45976 21272 45988
rect 21324 45976 21330 46028
rect 8021 45951 8079 45957
rect 8021 45948 8033 45951
rect 7800 45920 8033 45948
rect 7800 45908 7806 45920
rect 8021 45917 8033 45920
rect 8067 45917 8079 45951
rect 8021 45911 8079 45917
rect 9214 45908 9220 45960
rect 9272 45948 9278 45960
rect 9401 45951 9459 45957
rect 9401 45948 9413 45951
rect 9272 45920 9413 45948
rect 9272 45908 9278 45920
rect 9401 45917 9413 45920
rect 9447 45948 9459 45951
rect 10229 45951 10287 45957
rect 10229 45948 10241 45951
rect 9447 45920 10241 45948
rect 9447 45917 9459 45920
rect 9401 45911 9459 45917
rect 10229 45917 10241 45920
rect 10275 45917 10287 45951
rect 10686 45948 10692 45960
rect 10599 45920 10692 45948
rect 10229 45911 10287 45917
rect 3234 45880 3240 45892
rect 3195 45852 3240 45880
rect 3234 45840 3240 45852
rect 3292 45840 3298 45892
rect 4154 45880 4160 45892
rect 4115 45852 4160 45880
rect 4154 45840 4160 45852
rect 4212 45840 4218 45892
rect 10244 45812 10272 45911
rect 10686 45908 10692 45920
rect 10744 45908 10750 45960
rect 14182 45908 14188 45960
rect 14240 45948 14246 45960
rect 14277 45951 14335 45957
rect 14277 45948 14289 45951
rect 14240 45920 14289 45948
rect 14240 45908 14246 45920
rect 14277 45917 14289 45920
rect 14323 45917 14335 45951
rect 18322 45948 18328 45960
rect 18283 45920 18328 45948
rect 14277 45911 14335 45917
rect 18322 45908 18328 45920
rect 18380 45908 18386 45960
rect 23198 45948 23204 45960
rect 23159 45920 23204 45948
rect 23198 45908 23204 45920
rect 23256 45908 23262 45960
rect 24946 45908 24952 45960
rect 25004 45948 25010 45960
rect 25884 45957 25912 46056
rect 27430 46044 27436 46056
rect 27488 46044 27494 46096
rect 26510 46016 26516 46028
rect 26471 45988 26516 46016
rect 26510 45976 26516 45988
rect 26568 45976 26574 46028
rect 27706 46016 27712 46028
rect 27667 45988 27712 46016
rect 27706 45976 27712 45988
rect 27764 45976 27770 46028
rect 25225 45951 25283 45957
rect 25225 45948 25237 45951
rect 25004 45920 25237 45948
rect 25004 45908 25010 45920
rect 25225 45917 25237 45920
rect 25271 45917 25283 45951
rect 25225 45911 25283 45917
rect 25869 45951 25927 45957
rect 25869 45917 25881 45951
rect 25915 45917 25927 45951
rect 25869 45911 25927 45917
rect 10781 45883 10839 45889
rect 10781 45849 10793 45883
rect 10827 45880 10839 45883
rect 11517 45883 11575 45889
rect 11517 45880 11529 45883
rect 10827 45852 11529 45880
rect 10827 45849 10839 45852
rect 10781 45843 10839 45849
rect 11517 45849 11529 45852
rect 11563 45849 11575 45883
rect 20438 45880 20444 45892
rect 20399 45852 20444 45880
rect 11517 45843 11575 45849
rect 20438 45840 20444 45852
rect 20496 45840 20502 45892
rect 21266 45840 21272 45892
rect 21324 45880 21330 45892
rect 22554 45880 22560 45892
rect 21324 45852 22560 45880
rect 21324 45840 21330 45852
rect 22554 45840 22560 45852
rect 22612 45840 22618 45892
rect 25961 45883 26019 45889
rect 25961 45849 25973 45883
rect 26007 45880 26019 45883
rect 26697 45883 26755 45889
rect 26697 45880 26709 45883
rect 26007 45852 26709 45880
rect 26007 45849 26019 45852
rect 25961 45843 26019 45849
rect 26697 45849 26709 45852
rect 26743 45849 26755 45883
rect 26697 45843 26755 45849
rect 12710 45812 12716 45824
rect 10244 45784 12716 45812
rect 12710 45772 12716 45784
rect 12768 45812 12774 45824
rect 13262 45812 13268 45824
rect 12768 45784 13268 45812
rect 12768 45772 12774 45784
rect 13262 45772 13268 45784
rect 13320 45772 13326 45824
rect 15838 45772 15844 45824
rect 15896 45812 15902 45824
rect 20346 45812 20352 45824
rect 15896 45784 20352 45812
rect 15896 45772 15902 45784
rect 20346 45772 20352 45784
rect 20404 45772 20410 45824
rect 1104 45722 29048 45744
rect 1104 45670 7896 45722
rect 7948 45670 7960 45722
rect 8012 45670 8024 45722
rect 8076 45670 8088 45722
rect 8140 45670 8152 45722
rect 8204 45670 14842 45722
rect 14894 45670 14906 45722
rect 14958 45670 14970 45722
rect 15022 45670 15034 45722
rect 15086 45670 15098 45722
rect 15150 45670 21788 45722
rect 21840 45670 21852 45722
rect 21904 45670 21916 45722
rect 21968 45670 21980 45722
rect 22032 45670 22044 45722
rect 22096 45670 28734 45722
rect 28786 45670 28798 45722
rect 28850 45670 28862 45722
rect 28914 45670 28926 45722
rect 28978 45670 28990 45722
rect 29042 45670 29048 45722
rect 1104 45648 29048 45670
rect 13078 45568 13084 45620
rect 13136 45608 13142 45620
rect 13173 45611 13231 45617
rect 13173 45608 13185 45611
rect 13136 45580 13185 45608
rect 13136 45568 13142 45580
rect 13173 45577 13185 45580
rect 13219 45577 13231 45611
rect 13173 45571 13231 45577
rect 18322 45568 18328 45620
rect 18380 45608 18386 45620
rect 20438 45608 20444 45620
rect 18380 45580 20300 45608
rect 20399 45580 20444 45608
rect 18380 45568 18386 45580
rect 4065 45543 4123 45549
rect 4065 45509 4077 45543
rect 4111 45540 4123 45543
rect 4154 45540 4160 45552
rect 4111 45512 4160 45540
rect 4111 45509 4123 45512
rect 4065 45503 4123 45509
rect 4154 45500 4160 45512
rect 4212 45500 4218 45552
rect 18340 45540 18368 45568
rect 14016 45512 18368 45540
rect 20272 45540 20300 45580
rect 20438 45568 20444 45580
rect 20496 45568 20502 45620
rect 27706 45608 27712 45620
rect 20548 45580 27712 45608
rect 20548 45540 20576 45580
rect 27706 45568 27712 45580
rect 27764 45568 27770 45620
rect 20272 45512 20576 45540
rect 26421 45543 26479 45549
rect 1670 45472 1676 45484
rect 1631 45444 1676 45472
rect 1670 45432 1676 45444
rect 1728 45432 1734 45484
rect 3973 45475 4031 45481
rect 3973 45441 3985 45475
rect 4019 45441 4031 45475
rect 3973 45435 4031 45441
rect 1857 45407 1915 45413
rect 1857 45373 1869 45407
rect 1903 45404 1915 45407
rect 2038 45404 2044 45416
rect 1903 45376 2044 45404
rect 1903 45373 1915 45376
rect 1857 45367 1915 45373
rect 2038 45364 2044 45376
rect 2096 45364 2102 45416
rect 2133 45407 2191 45413
rect 2133 45373 2145 45407
rect 2179 45373 2191 45407
rect 2133 45367 2191 45373
rect 14 45296 20 45348
rect 72 45336 78 45348
rect 2148 45336 2176 45367
rect 2498 45364 2504 45416
rect 2556 45404 2562 45416
rect 3988 45404 4016 45435
rect 9306 45432 9312 45484
rect 9364 45472 9370 45484
rect 9677 45475 9735 45481
rect 9677 45472 9689 45475
rect 9364 45444 9689 45472
rect 9364 45432 9370 45444
rect 9677 45441 9689 45444
rect 9723 45441 9735 45475
rect 10410 45472 10416 45484
rect 10371 45444 10416 45472
rect 9677 45435 9735 45441
rect 10410 45432 10416 45444
rect 10468 45432 10474 45484
rect 13262 45472 13268 45484
rect 13175 45444 13268 45472
rect 13262 45432 13268 45444
rect 13320 45472 13326 45484
rect 14016 45472 14044 45512
rect 26421 45509 26433 45543
rect 26467 45540 26479 45543
rect 27246 45540 27252 45552
rect 26467 45512 27252 45540
rect 26467 45509 26479 45512
rect 26421 45503 26479 45509
rect 27246 45500 27252 45512
rect 27304 45500 27310 45552
rect 14182 45472 14188 45484
rect 13320 45444 14044 45472
rect 14143 45444 14188 45472
rect 13320 45432 13326 45444
rect 14182 45432 14188 45444
rect 14240 45432 14246 45484
rect 20346 45472 20352 45484
rect 20307 45444 20352 45472
rect 20346 45432 20352 45444
rect 20404 45432 20410 45484
rect 26605 45475 26663 45481
rect 26605 45441 26617 45475
rect 26651 45472 26663 45475
rect 27890 45472 27896 45484
rect 26651 45444 27896 45472
rect 26651 45441 26663 45444
rect 26605 45435 26663 45441
rect 27890 45432 27896 45444
rect 27948 45432 27954 45484
rect 14366 45404 14372 45416
rect 2556 45376 6914 45404
rect 14327 45376 14372 45404
rect 2556 45364 2562 45376
rect 72 45308 2176 45336
rect 6886 45336 6914 45376
rect 14366 45364 14372 45376
rect 14424 45364 14430 45416
rect 15194 45404 15200 45416
rect 15155 45376 15200 45404
rect 15194 45364 15200 45376
rect 15252 45364 15258 45416
rect 26050 45404 26056 45416
rect 26011 45376 26056 45404
rect 26050 45364 26056 45376
rect 26108 45364 26114 45416
rect 27982 45336 27988 45348
rect 6886 45308 27988 45336
rect 72 45296 78 45308
rect 27982 45296 27988 45308
rect 28040 45296 28046 45348
rect 20346 45228 20352 45280
rect 20404 45268 20410 45280
rect 21634 45268 21640 45280
rect 20404 45240 21640 45268
rect 20404 45228 20410 45240
rect 21634 45228 21640 45240
rect 21692 45268 21698 45280
rect 27338 45268 27344 45280
rect 21692 45240 27344 45268
rect 21692 45228 21698 45240
rect 27338 45228 27344 45240
rect 27396 45228 27402 45280
rect 27893 45271 27951 45277
rect 27893 45237 27905 45271
rect 27939 45268 27951 45271
rect 28350 45268 28356 45280
rect 27939 45240 28356 45268
rect 27939 45237 27951 45240
rect 27893 45231 27951 45237
rect 28350 45228 28356 45240
rect 28408 45228 28414 45280
rect 1104 45178 28888 45200
rect 1104 45126 4423 45178
rect 4475 45126 4487 45178
rect 4539 45126 4551 45178
rect 4603 45126 4615 45178
rect 4667 45126 4679 45178
rect 4731 45126 11369 45178
rect 11421 45126 11433 45178
rect 11485 45126 11497 45178
rect 11549 45126 11561 45178
rect 11613 45126 11625 45178
rect 11677 45126 18315 45178
rect 18367 45126 18379 45178
rect 18431 45126 18443 45178
rect 18495 45126 18507 45178
rect 18559 45126 18571 45178
rect 18623 45126 25261 45178
rect 25313 45126 25325 45178
rect 25377 45126 25389 45178
rect 25441 45126 25453 45178
rect 25505 45126 25517 45178
rect 25569 45126 28888 45178
rect 1104 45104 28888 45126
rect 2038 45064 2044 45076
rect 1999 45036 2044 45064
rect 2038 45024 2044 45036
rect 2096 45024 2102 45076
rect 3329 45067 3387 45073
rect 3329 45033 3341 45067
rect 3375 45064 3387 45067
rect 3970 45064 3976 45076
rect 3375 45036 3976 45064
rect 3375 45033 3387 45036
rect 3329 45027 3387 45033
rect 3970 45024 3976 45036
rect 4028 45024 4034 45076
rect 27522 44928 27528 44940
rect 27483 44900 27528 44928
rect 27522 44888 27528 44900
rect 27580 44888 27586 44940
rect 28350 44928 28356 44940
rect 28311 44900 28356 44928
rect 28350 44888 28356 44900
rect 28408 44888 28414 44940
rect 2133 44863 2191 44869
rect 2133 44829 2145 44863
rect 2179 44860 2191 44863
rect 2498 44860 2504 44872
rect 2179 44832 2504 44860
rect 2179 44829 2191 44832
rect 2133 44823 2191 44829
rect 2498 44820 2504 44832
rect 2556 44820 2562 44872
rect 5166 44820 5172 44872
rect 5224 44860 5230 44872
rect 23198 44860 23204 44872
rect 5224 44832 23204 44860
rect 5224 44820 5230 44832
rect 23198 44820 23204 44832
rect 23256 44820 23262 44872
rect 26053 44863 26111 44869
rect 26053 44829 26065 44863
rect 26099 44860 26111 44863
rect 26234 44860 26240 44872
rect 26099 44832 26240 44860
rect 26099 44829 26111 44832
rect 26053 44823 26111 44829
rect 26234 44820 26240 44832
rect 26292 44820 26298 44872
rect 27890 44752 27896 44804
rect 27948 44792 27954 44804
rect 28169 44795 28227 44801
rect 28169 44792 28181 44795
rect 27948 44764 28181 44792
rect 27948 44752 27954 44764
rect 28169 44761 28181 44764
rect 28215 44761 28227 44795
rect 28169 44755 28227 44761
rect 1104 44634 29048 44656
rect 1104 44582 7896 44634
rect 7948 44582 7960 44634
rect 8012 44582 8024 44634
rect 8076 44582 8088 44634
rect 8140 44582 8152 44634
rect 8204 44582 14842 44634
rect 14894 44582 14906 44634
rect 14958 44582 14970 44634
rect 15022 44582 15034 44634
rect 15086 44582 15098 44634
rect 15150 44582 21788 44634
rect 21840 44582 21852 44634
rect 21904 44582 21916 44634
rect 21968 44582 21980 44634
rect 22032 44582 22044 44634
rect 22096 44582 28734 44634
rect 28786 44582 28798 44634
rect 28850 44582 28862 44634
rect 28914 44582 28926 44634
rect 28978 44582 28990 44634
rect 29042 44582 29048 44634
rect 1104 44560 29048 44582
rect 2133 44523 2191 44529
rect 2133 44489 2145 44523
rect 2179 44520 2191 44523
rect 3234 44520 3240 44532
rect 2179 44492 3240 44520
rect 2179 44489 2191 44492
rect 2133 44483 2191 44489
rect 3234 44480 3240 44492
rect 3292 44480 3298 44532
rect 14277 44523 14335 44529
rect 14277 44489 14289 44523
rect 14323 44520 14335 44523
rect 14366 44520 14372 44532
rect 14323 44492 14372 44520
rect 14323 44489 14335 44492
rect 14277 44483 14335 44489
rect 14366 44480 14372 44492
rect 14424 44480 14430 44532
rect 27890 44520 27896 44532
rect 27851 44492 27896 44520
rect 27890 44480 27896 44492
rect 27948 44480 27954 44532
rect 24949 44455 25007 44461
rect 24949 44421 24961 44455
rect 24995 44452 25007 44455
rect 25038 44452 25044 44464
rect 24995 44424 25044 44452
rect 24995 44421 25007 44424
rect 24949 44415 25007 44421
rect 25038 44412 25044 44424
rect 25096 44412 25102 44464
rect 2225 44387 2283 44393
rect 2225 44353 2237 44387
rect 2271 44384 2283 44387
rect 4338 44384 4344 44396
rect 2271 44356 4344 44384
rect 2271 44353 2283 44356
rect 2225 44347 2283 44353
rect 4338 44344 4344 44356
rect 4396 44384 4402 44396
rect 5166 44384 5172 44396
rect 4396 44356 5172 44384
rect 4396 44344 4402 44356
rect 5166 44344 5172 44356
rect 5224 44344 5230 44396
rect 14185 44387 14243 44393
rect 14185 44353 14197 44387
rect 14231 44384 14243 44387
rect 14366 44384 14372 44396
rect 14231 44356 14372 44384
rect 14231 44353 14243 44356
rect 14185 44347 14243 44353
rect 14366 44344 14372 44356
rect 14424 44384 14430 44396
rect 19334 44384 19340 44396
rect 14424 44356 19340 44384
rect 14424 44344 14430 44356
rect 19334 44344 19340 44356
rect 19392 44344 19398 44396
rect 27154 44384 27160 44396
rect 27115 44356 27160 44384
rect 27154 44344 27160 44356
rect 27212 44344 27218 44396
rect 27801 44387 27859 44393
rect 27801 44353 27813 44387
rect 27847 44384 27859 44387
rect 27982 44384 27988 44396
rect 27847 44356 27988 44384
rect 27847 44353 27859 44356
rect 27801 44347 27859 44353
rect 27982 44344 27988 44356
rect 28040 44344 28046 44396
rect 24765 44319 24823 44325
rect 24765 44285 24777 44319
rect 24811 44316 24823 44319
rect 24946 44316 24952 44328
rect 24811 44288 24952 44316
rect 24811 44285 24823 44288
rect 24765 44279 24823 44285
rect 24946 44276 24952 44288
rect 25004 44276 25010 44328
rect 26142 44316 26148 44328
rect 26103 44288 26148 44316
rect 26142 44276 26148 44288
rect 26200 44276 26206 44328
rect 2958 44180 2964 44192
rect 2919 44152 2964 44180
rect 2958 44140 2964 44152
rect 3016 44140 3022 44192
rect 26418 44140 26424 44192
rect 26476 44180 26482 44192
rect 27249 44183 27307 44189
rect 27249 44180 27261 44183
rect 26476 44152 27261 44180
rect 26476 44140 26482 44152
rect 27249 44149 27261 44152
rect 27295 44149 27307 44183
rect 27249 44143 27307 44149
rect 1104 44090 28888 44112
rect 1104 44038 4423 44090
rect 4475 44038 4487 44090
rect 4539 44038 4551 44090
rect 4603 44038 4615 44090
rect 4667 44038 4679 44090
rect 4731 44038 11369 44090
rect 11421 44038 11433 44090
rect 11485 44038 11497 44090
rect 11549 44038 11561 44090
rect 11613 44038 11625 44090
rect 11677 44038 18315 44090
rect 18367 44038 18379 44090
rect 18431 44038 18443 44090
rect 18495 44038 18507 44090
rect 18559 44038 18571 44090
rect 18623 44038 25261 44090
rect 25313 44038 25325 44090
rect 25377 44038 25389 44090
rect 25441 44038 25453 44090
rect 25505 44038 25517 44090
rect 25569 44038 28888 44090
rect 1104 44016 28888 44038
rect 2501 43979 2559 43985
rect 2501 43945 2513 43979
rect 2547 43976 2559 43979
rect 3418 43976 3424 43988
rect 2547 43948 3424 43976
rect 2547 43945 2559 43948
rect 2501 43939 2559 43945
rect 3418 43936 3424 43948
rect 3476 43936 3482 43988
rect 21266 43840 21272 43852
rect 21227 43812 21272 43840
rect 21266 43800 21272 43812
rect 21324 43800 21330 43852
rect 26234 43800 26240 43852
rect 26292 43840 26298 43852
rect 26292 43812 26337 43840
rect 26292 43800 26298 43812
rect 26418 43800 26424 43852
rect 26476 43840 26482 43852
rect 28074 43840 28080 43852
rect 26476 43812 26521 43840
rect 28035 43812 28080 43840
rect 26476 43800 26482 43812
rect 28074 43800 28080 43812
rect 28132 43800 28138 43852
rect 1578 43732 1584 43784
rect 1636 43772 1642 43784
rect 1673 43775 1731 43781
rect 1673 43772 1685 43775
rect 1636 43744 1685 43772
rect 1636 43732 1642 43744
rect 1673 43741 1685 43744
rect 1719 43741 1731 43775
rect 1673 43735 1731 43741
rect 3329 43775 3387 43781
rect 3329 43741 3341 43775
rect 3375 43772 3387 43775
rect 5074 43772 5080 43784
rect 3375 43744 5080 43772
rect 3375 43741 3387 43744
rect 3329 43735 3387 43741
rect 5074 43732 5080 43744
rect 5132 43772 5138 43784
rect 10686 43772 10692 43784
rect 5132 43744 10692 43772
rect 5132 43732 5138 43744
rect 10686 43732 10692 43744
rect 10744 43732 10750 43784
rect 19426 43772 19432 43784
rect 19387 43744 19432 43772
rect 19426 43732 19432 43744
rect 19484 43732 19490 43784
rect 19610 43704 19616 43716
rect 19571 43676 19616 43704
rect 19610 43664 19616 43676
rect 19668 43664 19674 43716
rect 3142 43596 3148 43648
rect 3200 43636 3206 43648
rect 3237 43639 3295 43645
rect 3237 43636 3249 43639
rect 3200 43608 3249 43636
rect 3200 43596 3206 43608
rect 3237 43605 3249 43608
rect 3283 43605 3295 43639
rect 3237 43599 3295 43605
rect 1104 43546 29048 43568
rect 1104 43494 7896 43546
rect 7948 43494 7960 43546
rect 8012 43494 8024 43546
rect 8076 43494 8088 43546
rect 8140 43494 8152 43546
rect 8204 43494 14842 43546
rect 14894 43494 14906 43546
rect 14958 43494 14970 43546
rect 15022 43494 15034 43546
rect 15086 43494 15098 43546
rect 15150 43494 21788 43546
rect 21840 43494 21852 43546
rect 21904 43494 21916 43546
rect 21968 43494 21980 43546
rect 22032 43494 22044 43546
rect 22096 43494 28734 43546
rect 28786 43494 28798 43546
rect 28850 43494 28862 43546
rect 28914 43494 28926 43546
rect 28978 43494 28990 43546
rect 29042 43494 29048 43546
rect 1104 43472 29048 43494
rect 3050 43392 3056 43444
rect 3108 43432 3114 43444
rect 15838 43432 15844 43444
rect 3108 43404 15844 43432
rect 3108 43392 3114 43404
rect 15838 43392 15844 43404
rect 15896 43392 15902 43444
rect 19521 43435 19579 43441
rect 19521 43401 19533 43435
rect 19567 43432 19579 43435
rect 19610 43432 19616 43444
rect 19567 43404 19616 43432
rect 19567 43401 19579 43404
rect 19521 43395 19579 43401
rect 19610 43392 19616 43404
rect 19668 43392 19674 43444
rect 3142 43364 3148 43376
rect 3103 43336 3148 43364
rect 3142 43324 3148 43336
rect 3200 43324 3206 43376
rect 2225 43299 2283 43305
rect 2225 43265 2237 43299
rect 2271 43265 2283 43299
rect 2958 43296 2964 43308
rect 2919 43268 2964 43296
rect 2225 43259 2283 43265
rect 2240 43228 2268 43259
rect 2958 43256 2964 43268
rect 3016 43256 3022 43308
rect 19334 43256 19340 43308
rect 19392 43296 19398 43308
rect 19429 43299 19487 43305
rect 19429 43296 19441 43299
rect 19392 43268 19441 43296
rect 19392 43256 19398 43268
rect 19429 43265 19441 43268
rect 19475 43296 19487 43299
rect 26145 43299 26203 43305
rect 26145 43296 26157 43299
rect 19475 43268 26157 43296
rect 19475 43265 19487 43268
rect 19429 43259 19487 43265
rect 26145 43265 26157 43268
rect 26191 43296 26203 43299
rect 27154 43296 27160 43308
rect 26191 43268 27160 43296
rect 26191 43265 26203 43268
rect 26145 43259 26203 43265
rect 27154 43256 27160 43268
rect 27212 43256 27218 43308
rect 4154 43228 4160 43240
rect 2240 43200 3096 43228
rect 4115 43200 4160 43228
rect 3068 43172 3096 43200
rect 4154 43188 4160 43200
rect 4212 43188 4218 43240
rect 3050 43120 3056 43172
rect 3108 43120 3114 43172
rect 1762 43052 1768 43104
rect 1820 43092 1826 43104
rect 2133 43095 2191 43101
rect 2133 43092 2145 43095
rect 1820 43064 2145 43092
rect 1820 43052 1826 43064
rect 2133 43061 2145 43064
rect 2179 43061 2191 43095
rect 2133 43055 2191 43061
rect 26237 43095 26295 43101
rect 26237 43061 26249 43095
rect 26283 43092 26295 43095
rect 26694 43092 26700 43104
rect 26283 43064 26700 43092
rect 26283 43061 26295 43064
rect 26237 43055 26295 43061
rect 26694 43052 26700 43064
rect 26752 43052 26758 43104
rect 27154 43092 27160 43104
rect 27115 43064 27160 43092
rect 27154 43052 27160 43064
rect 27212 43052 27218 43104
rect 28074 43092 28080 43104
rect 28035 43064 28080 43092
rect 28074 43052 28080 43064
rect 28132 43052 28138 43104
rect 1104 43002 28888 43024
rect 1104 42950 4423 43002
rect 4475 42950 4487 43002
rect 4539 42950 4551 43002
rect 4603 42950 4615 43002
rect 4667 42950 4679 43002
rect 4731 42950 11369 43002
rect 11421 42950 11433 43002
rect 11485 42950 11497 43002
rect 11549 42950 11561 43002
rect 11613 42950 11625 43002
rect 11677 42950 18315 43002
rect 18367 42950 18379 43002
rect 18431 42950 18443 43002
rect 18495 42950 18507 43002
rect 18559 42950 18571 43002
rect 18623 42950 25261 43002
rect 25313 42950 25325 43002
rect 25377 42950 25389 43002
rect 25441 42950 25453 43002
rect 25505 42950 25517 43002
rect 25569 42950 28888 43002
rect 1104 42928 28888 42950
rect 1578 42752 1584 42764
rect 1539 42724 1584 42752
rect 1578 42712 1584 42724
rect 1636 42712 1642 42764
rect 1762 42752 1768 42764
rect 1723 42724 1768 42752
rect 1762 42712 1768 42724
rect 1820 42712 1826 42764
rect 2774 42752 2780 42764
rect 2735 42724 2780 42752
rect 2774 42712 2780 42724
rect 2832 42712 2838 42764
rect 26513 42755 26571 42761
rect 26513 42721 26525 42755
rect 26559 42752 26571 42755
rect 27154 42752 27160 42764
rect 26559 42724 27160 42752
rect 26559 42721 26571 42724
rect 26513 42715 26571 42721
rect 27154 42712 27160 42724
rect 27212 42712 27218 42764
rect 28350 42752 28356 42764
rect 28311 42724 28356 42752
rect 28350 42712 28356 42724
rect 28408 42712 28414 42764
rect 26694 42616 26700 42628
rect 26655 42588 26700 42616
rect 26694 42576 26700 42588
rect 26752 42576 26758 42628
rect 1104 42458 29048 42480
rect 1104 42406 7896 42458
rect 7948 42406 7960 42458
rect 8012 42406 8024 42458
rect 8076 42406 8088 42458
rect 8140 42406 8152 42458
rect 8204 42406 14842 42458
rect 14894 42406 14906 42458
rect 14958 42406 14970 42458
rect 15022 42406 15034 42458
rect 15086 42406 15098 42458
rect 15150 42406 21788 42458
rect 21840 42406 21852 42458
rect 21904 42406 21916 42458
rect 21968 42406 21980 42458
rect 22032 42406 22044 42458
rect 22096 42406 28734 42458
rect 28786 42406 28798 42458
rect 28850 42406 28862 42458
rect 28914 42406 28926 42458
rect 28978 42406 28990 42458
rect 29042 42406 29048 42458
rect 1104 42384 29048 42406
rect 2685 42211 2743 42217
rect 2685 42177 2697 42211
rect 2731 42208 2743 42211
rect 2866 42208 2872 42220
rect 2731 42180 2872 42208
rect 2731 42177 2743 42180
rect 2685 42171 2743 42177
rect 2866 42168 2872 42180
rect 2924 42168 2930 42220
rect 27706 42208 27712 42220
rect 27667 42180 27712 42208
rect 27706 42168 27712 42180
rect 27764 42168 27770 42220
rect 1670 42004 1676 42016
rect 1631 41976 1676 42004
rect 1670 41964 1676 41976
rect 1728 41964 1734 42016
rect 2593 42007 2651 42013
rect 2593 41973 2605 42007
rect 2639 42004 2651 42007
rect 3234 42004 3240 42016
rect 2639 41976 3240 42004
rect 2639 41973 2651 41976
rect 2593 41967 2651 41973
rect 3234 41964 3240 41976
rect 3292 41964 3298 42016
rect 3329 42007 3387 42013
rect 3329 41973 3341 42007
rect 3375 42004 3387 42007
rect 3418 42004 3424 42016
rect 3375 41976 3424 42004
rect 3375 41973 3387 41976
rect 3329 41967 3387 41973
rect 3418 41964 3424 41976
rect 3476 41964 3482 42016
rect 27801 42007 27859 42013
rect 27801 41973 27813 42007
rect 27847 42004 27859 42007
rect 28166 42004 28172 42016
rect 27847 41976 28172 42004
rect 27847 41973 27859 41976
rect 27801 41967 27859 41973
rect 28166 41964 28172 41976
rect 28224 41964 28230 42016
rect 1104 41914 28888 41936
rect 1104 41862 4423 41914
rect 4475 41862 4487 41914
rect 4539 41862 4551 41914
rect 4603 41862 4615 41914
rect 4667 41862 4679 41914
rect 4731 41862 11369 41914
rect 11421 41862 11433 41914
rect 11485 41862 11497 41914
rect 11549 41862 11561 41914
rect 11613 41862 11625 41914
rect 11677 41862 18315 41914
rect 18367 41862 18379 41914
rect 18431 41862 18443 41914
rect 18495 41862 18507 41914
rect 18559 41862 18571 41914
rect 18623 41862 25261 41914
rect 25313 41862 25325 41914
rect 25377 41862 25389 41914
rect 25441 41862 25453 41914
rect 25505 41862 25517 41914
rect 25569 41862 28888 41914
rect 1104 41840 28888 41862
rect 28074 41692 28080 41744
rect 28132 41732 28138 41744
rect 28132 41704 28396 41732
rect 28132 41692 28138 41704
rect 3234 41664 3240 41676
rect 3195 41636 3240 41664
rect 3234 41624 3240 41636
rect 3292 41624 3298 41676
rect 3418 41664 3424 41676
rect 3379 41636 3424 41664
rect 3418 41624 3424 41636
rect 3476 41624 3482 41676
rect 27522 41664 27528 41676
rect 27483 41636 27528 41664
rect 27522 41624 27528 41636
rect 27580 41624 27586 41676
rect 28166 41664 28172 41676
rect 28127 41636 28172 41664
rect 28166 41624 28172 41636
rect 28224 41624 28230 41676
rect 28368 41673 28396 41704
rect 28353 41667 28411 41673
rect 28353 41633 28365 41667
rect 28399 41633 28411 41667
rect 28353 41627 28411 41633
rect 1578 41596 1584 41608
rect 1539 41568 1584 41596
rect 1578 41556 1584 41568
rect 1636 41556 1642 41608
rect 1104 41370 29048 41392
rect 1104 41318 7896 41370
rect 7948 41318 7960 41370
rect 8012 41318 8024 41370
rect 8076 41318 8088 41370
rect 8140 41318 8152 41370
rect 8204 41318 14842 41370
rect 14894 41318 14906 41370
rect 14958 41318 14970 41370
rect 15022 41318 15034 41370
rect 15086 41318 15098 41370
rect 15150 41318 21788 41370
rect 21840 41318 21852 41370
rect 21904 41318 21916 41370
rect 21968 41318 21980 41370
rect 22032 41318 22044 41370
rect 22096 41318 28734 41370
rect 28786 41318 28798 41370
rect 28850 41318 28862 41370
rect 28914 41318 28926 41370
rect 28978 41318 28990 41370
rect 29042 41318 29048 41370
rect 1104 41296 29048 41318
rect 1670 41120 1676 41132
rect 1631 41092 1676 41120
rect 1670 41080 1676 41092
rect 1728 41080 1734 41132
rect 27430 41120 27436 41132
rect 27391 41092 27436 41120
rect 27430 41080 27436 41092
rect 27488 41080 27494 41132
rect 1857 41055 1915 41061
rect 1857 41021 1869 41055
rect 1903 41052 1915 41055
rect 2314 41052 2320 41064
rect 1903 41024 2320 41052
rect 1903 41021 1915 41024
rect 1857 41015 1915 41021
rect 2314 41012 2320 41024
rect 2372 41012 2378 41064
rect 2774 41052 2780 41064
rect 2735 41024 2780 41052
rect 2774 41012 2780 41024
rect 2832 41012 2838 41064
rect 27525 40919 27583 40925
rect 27525 40885 27537 40919
rect 27571 40916 27583 40919
rect 28166 40916 28172 40928
rect 27571 40888 28172 40916
rect 27571 40885 27583 40888
rect 27525 40879 27583 40885
rect 28166 40876 28172 40888
rect 28224 40876 28230 40928
rect 28261 40919 28319 40925
rect 28261 40885 28273 40919
rect 28307 40916 28319 40919
rect 28350 40916 28356 40928
rect 28307 40888 28356 40916
rect 28307 40885 28319 40888
rect 28261 40879 28319 40885
rect 28350 40876 28356 40888
rect 28408 40876 28414 40928
rect 1104 40826 28888 40848
rect 1104 40774 4423 40826
rect 4475 40774 4487 40826
rect 4539 40774 4551 40826
rect 4603 40774 4615 40826
rect 4667 40774 4679 40826
rect 4731 40774 11369 40826
rect 11421 40774 11433 40826
rect 11485 40774 11497 40826
rect 11549 40774 11561 40826
rect 11613 40774 11625 40826
rect 11677 40774 18315 40826
rect 18367 40774 18379 40826
rect 18431 40774 18443 40826
rect 18495 40774 18507 40826
rect 18559 40774 18571 40826
rect 18623 40774 25261 40826
rect 25313 40774 25325 40826
rect 25377 40774 25389 40826
rect 25441 40774 25453 40826
rect 25505 40774 25517 40826
rect 25569 40774 28888 40826
rect 1104 40752 28888 40774
rect 27522 40576 27528 40588
rect 27483 40548 27528 40576
rect 27522 40536 27528 40548
rect 27580 40536 27586 40588
rect 28166 40576 28172 40588
rect 28127 40548 28172 40576
rect 28166 40536 28172 40548
rect 28224 40536 28230 40588
rect 28350 40576 28356 40588
rect 28311 40548 28356 40576
rect 28350 40536 28356 40548
rect 28408 40536 28414 40588
rect 1946 40508 1952 40520
rect 1907 40480 1952 40508
rect 1946 40468 1952 40480
rect 2004 40468 2010 40520
rect 2406 40508 2412 40520
rect 2367 40480 2412 40508
rect 2406 40468 2412 40480
rect 2464 40468 2470 40520
rect 17773 40511 17831 40517
rect 17773 40477 17785 40511
rect 17819 40508 17831 40511
rect 17862 40508 17868 40520
rect 17819 40480 17868 40508
rect 17819 40477 17831 40480
rect 17773 40471 17831 40477
rect 17862 40468 17868 40480
rect 17920 40468 17926 40520
rect 18598 40508 18604 40520
rect 18559 40480 18604 40508
rect 18598 40468 18604 40480
rect 18656 40468 18662 40520
rect 18785 40511 18843 40517
rect 18785 40477 18797 40511
rect 18831 40477 18843 40511
rect 18785 40471 18843 40477
rect 18230 40400 18236 40452
rect 18288 40440 18294 40452
rect 18800 40440 18828 40471
rect 18288 40412 18828 40440
rect 18288 40400 18294 40412
rect 1854 40372 1860 40384
rect 1815 40344 1860 40372
rect 1854 40332 1860 40344
rect 1912 40332 1918 40384
rect 17494 40332 17500 40384
rect 17552 40372 17558 40384
rect 17681 40375 17739 40381
rect 17681 40372 17693 40375
rect 17552 40344 17693 40372
rect 17552 40332 17558 40344
rect 17681 40341 17693 40344
rect 17727 40341 17739 40375
rect 18690 40372 18696 40384
rect 18651 40344 18696 40372
rect 17681 40335 17739 40341
rect 18690 40332 18696 40344
rect 18748 40332 18754 40384
rect 1104 40282 29048 40304
rect 1104 40230 7896 40282
rect 7948 40230 7960 40282
rect 8012 40230 8024 40282
rect 8076 40230 8088 40282
rect 8140 40230 8152 40282
rect 8204 40230 14842 40282
rect 14894 40230 14906 40282
rect 14958 40230 14970 40282
rect 15022 40230 15034 40282
rect 15086 40230 15098 40282
rect 15150 40230 21788 40282
rect 21840 40230 21852 40282
rect 21904 40230 21916 40282
rect 21968 40230 21980 40282
rect 22032 40230 22044 40282
rect 22096 40230 28734 40282
rect 28786 40230 28798 40282
rect 28850 40230 28862 40282
rect 28914 40230 28926 40282
rect 28978 40230 28990 40282
rect 29042 40230 29048 40282
rect 1104 40208 29048 40230
rect 18309 40171 18367 40177
rect 18309 40137 18321 40171
rect 18355 40168 18367 40171
rect 18598 40168 18604 40180
rect 18355 40140 18604 40168
rect 18355 40137 18367 40140
rect 18309 40131 18367 40137
rect 18598 40128 18604 40140
rect 18656 40168 18662 40180
rect 19242 40168 19248 40180
rect 18656 40140 19248 40168
rect 18656 40128 18662 40140
rect 19242 40128 19248 40140
rect 19300 40128 19306 40180
rect 1854 40100 1860 40112
rect 1815 40072 1860 40100
rect 1854 40060 1860 40072
rect 1912 40060 1918 40112
rect 3510 40100 3516 40112
rect 3471 40072 3516 40100
rect 3510 40060 3516 40072
rect 3568 40060 3574 40112
rect 17862 40060 17868 40112
rect 17920 40100 17926 40112
rect 18509 40103 18567 40109
rect 18509 40100 18521 40103
rect 17920 40072 18521 40100
rect 17920 40060 17926 40072
rect 18509 40069 18521 40072
rect 18555 40069 18567 40103
rect 18509 40063 18567 40069
rect 17218 40032 17224 40044
rect 17179 40004 17224 40032
rect 17218 39992 17224 40004
rect 17276 39992 17282 40044
rect 17494 40032 17500 40044
rect 17455 40004 17500 40032
rect 17494 39992 17500 40004
rect 17552 39992 17558 40044
rect 17681 40035 17739 40041
rect 17681 40001 17693 40035
rect 17727 40032 17739 40035
rect 18874 40032 18880 40044
rect 17727 40004 18880 40032
rect 17727 40001 17739 40004
rect 17681 39995 17739 40001
rect 18874 39992 18880 40004
rect 18932 39992 18938 40044
rect 19610 40032 19616 40044
rect 19571 40004 19616 40032
rect 19610 39992 19616 40004
rect 19668 39992 19674 40044
rect 1673 39967 1731 39973
rect 1673 39933 1685 39967
rect 1719 39964 1731 39967
rect 2406 39964 2412 39976
rect 1719 39936 2412 39964
rect 1719 39933 1731 39936
rect 1673 39927 1731 39933
rect 2406 39924 2412 39936
rect 2464 39924 2470 39976
rect 16298 39924 16304 39976
rect 16356 39964 16362 39976
rect 17405 39967 17463 39973
rect 17405 39964 17417 39967
rect 16356 39936 17417 39964
rect 16356 39924 16362 39936
rect 17405 39933 17417 39936
rect 17451 39964 17463 39967
rect 19797 39967 19855 39973
rect 17451 39936 18184 39964
rect 17451 39933 17463 39936
rect 17405 39927 17463 39933
rect 17310 39896 17316 39908
rect 17271 39868 17316 39896
rect 17310 39856 17316 39868
rect 17368 39856 17374 39908
rect 18156 39905 18184 39936
rect 19797 39933 19809 39967
rect 19843 39964 19855 39967
rect 20898 39964 20904 39976
rect 19843 39936 20904 39964
rect 19843 39933 19855 39936
rect 19797 39927 19855 39933
rect 20898 39924 20904 39936
rect 20956 39924 20962 39976
rect 18141 39899 18199 39905
rect 18141 39865 18153 39899
rect 18187 39865 18199 39899
rect 18141 39859 18199 39865
rect 17034 39828 17040 39840
rect 16995 39800 17040 39828
rect 17034 39788 17040 39800
rect 17092 39788 17098 39840
rect 18230 39788 18236 39840
rect 18288 39828 18294 39840
rect 18325 39831 18383 39837
rect 18325 39828 18337 39831
rect 18288 39800 18337 39828
rect 18288 39788 18294 39800
rect 18325 39797 18337 39800
rect 18371 39797 18383 39831
rect 18325 39791 18383 39797
rect 19242 39788 19248 39840
rect 19300 39828 19306 39840
rect 19429 39831 19487 39837
rect 19429 39828 19441 39831
rect 19300 39800 19441 39828
rect 19300 39788 19306 39800
rect 19429 39797 19441 39800
rect 19475 39797 19487 39831
rect 19429 39791 19487 39797
rect 26510 39788 26516 39840
rect 26568 39828 26574 39840
rect 27341 39831 27399 39837
rect 27341 39828 27353 39831
rect 26568 39800 27353 39828
rect 26568 39788 26574 39800
rect 27341 39797 27353 39800
rect 27387 39797 27399 39831
rect 27341 39791 27399 39797
rect 27522 39788 27528 39840
rect 27580 39828 27586 39840
rect 27985 39831 28043 39837
rect 27985 39828 27997 39831
rect 27580 39800 27997 39828
rect 27580 39788 27586 39800
rect 27985 39797 27997 39800
rect 28031 39797 28043 39831
rect 27985 39791 28043 39797
rect 1104 39738 28888 39760
rect 1104 39686 4423 39738
rect 4475 39686 4487 39738
rect 4539 39686 4551 39738
rect 4603 39686 4615 39738
rect 4667 39686 4679 39738
rect 4731 39686 11369 39738
rect 11421 39686 11433 39738
rect 11485 39686 11497 39738
rect 11549 39686 11561 39738
rect 11613 39686 11625 39738
rect 11677 39686 18315 39738
rect 18367 39686 18379 39738
rect 18431 39686 18443 39738
rect 18495 39686 18507 39738
rect 18559 39686 18571 39738
rect 18623 39686 25261 39738
rect 25313 39686 25325 39738
rect 25377 39686 25389 39738
rect 25441 39686 25453 39738
rect 25505 39686 25517 39738
rect 25569 39686 28888 39738
rect 1104 39664 28888 39686
rect 2314 39624 2320 39636
rect 2275 39596 2320 39624
rect 2314 39584 2320 39596
rect 2372 39584 2378 39636
rect 17310 39584 17316 39636
rect 17368 39624 17374 39636
rect 17497 39627 17555 39633
rect 17497 39624 17509 39627
rect 17368 39596 17509 39624
rect 17368 39584 17374 39596
rect 17497 39593 17509 39596
rect 17543 39593 17555 39627
rect 17497 39587 17555 39593
rect 18230 39556 18236 39568
rect 17696 39528 18236 39556
rect 1946 39448 1952 39500
rect 2004 39488 2010 39500
rect 2004 39460 2452 39488
rect 2004 39448 2010 39460
rect 2424 39429 2452 39460
rect 17696 39429 17724 39528
rect 18230 39516 18236 39528
rect 18288 39516 18294 39568
rect 18509 39559 18567 39565
rect 18509 39525 18521 39559
rect 18555 39556 18567 39559
rect 18690 39556 18696 39568
rect 18555 39528 18696 39556
rect 18555 39525 18567 39528
rect 18509 39519 18567 39525
rect 18690 39516 18696 39528
rect 18748 39516 18754 39568
rect 18874 39516 18880 39568
rect 18932 39556 18938 39568
rect 18932 39528 20208 39556
rect 18932 39516 18938 39528
rect 19242 39488 19248 39500
rect 17788 39460 19248 39488
rect 17788 39429 17816 39460
rect 19242 39448 19248 39460
rect 19300 39488 19306 39500
rect 19889 39491 19947 39497
rect 19889 39488 19901 39491
rect 19300 39460 19901 39488
rect 19300 39448 19306 39460
rect 19889 39457 19901 39460
rect 19935 39457 19947 39491
rect 19889 39451 19947 39457
rect 1581 39423 1639 39429
rect 1581 39389 1593 39423
rect 1627 39420 1639 39423
rect 2409 39423 2467 39429
rect 1627 39392 2360 39420
rect 1627 39389 1639 39392
rect 1581 39383 1639 39389
rect 2332 39352 2360 39392
rect 2409 39389 2421 39423
rect 2455 39389 2467 39423
rect 2409 39383 2467 39389
rect 17681 39423 17739 39429
rect 17681 39389 17693 39423
rect 17727 39389 17739 39423
rect 17681 39383 17739 39389
rect 17773 39423 17831 39429
rect 17773 39389 17785 39423
rect 17819 39389 17831 39423
rect 17773 39383 17831 39389
rect 18417 39423 18475 39429
rect 18417 39389 18429 39423
rect 18463 39389 18475 39423
rect 18598 39420 18604 39432
rect 18559 39392 18604 39420
rect 18417 39383 18475 39389
rect 2866 39352 2872 39364
rect 2332 39324 2872 39352
rect 2866 39312 2872 39324
rect 2924 39312 2930 39364
rect 17497 39355 17555 39361
rect 17497 39321 17509 39355
rect 17543 39352 17555 39355
rect 17862 39352 17868 39364
rect 17543 39324 17868 39352
rect 17543 39321 17555 39324
rect 17497 39315 17555 39321
rect 17862 39312 17868 39324
rect 17920 39312 17926 39364
rect 18432 39352 18460 39383
rect 18598 39380 18604 39392
rect 18656 39380 18662 39432
rect 18690 39380 18696 39432
rect 18748 39420 18754 39432
rect 18748 39392 18793 39420
rect 18748 39380 18754 39392
rect 18874 39380 18880 39432
rect 18932 39420 18938 39432
rect 19705 39423 19763 39429
rect 18932 39392 18977 39420
rect 18932 39380 18938 39392
rect 19705 39389 19717 39423
rect 19751 39389 19763 39423
rect 19705 39383 19763 39389
rect 19720 39352 19748 39383
rect 19794 39380 19800 39432
rect 19852 39420 19858 39432
rect 20180 39429 20208 39528
rect 26510 39488 26516 39500
rect 26471 39460 26516 39488
rect 26510 39448 26516 39460
rect 26568 39448 26574 39500
rect 28353 39491 28411 39497
rect 28353 39457 28365 39491
rect 28399 39488 28411 39491
rect 28626 39488 28632 39500
rect 28399 39460 28632 39488
rect 28399 39457 28411 39460
rect 28353 39451 28411 39457
rect 28626 39448 28632 39460
rect 28684 39448 28690 39500
rect 19981 39423 20039 39429
rect 19852 39392 19897 39420
rect 19852 39380 19858 39392
rect 19981 39389 19993 39423
rect 20027 39389 20039 39423
rect 19981 39383 20039 39389
rect 20165 39423 20223 39429
rect 20165 39389 20177 39423
rect 20211 39420 20223 39423
rect 20254 39420 20260 39432
rect 20211 39392 20260 39420
rect 20211 39389 20223 39392
rect 20165 39383 20223 39389
rect 17972 39324 19748 39352
rect 19996 39352 20024 39383
rect 20254 39380 20260 39392
rect 20312 39380 20318 39432
rect 20809 39423 20867 39429
rect 20809 39389 20821 39423
rect 20855 39420 20867 39423
rect 20898 39420 20904 39432
rect 20855 39392 20904 39420
rect 20855 39389 20867 39392
rect 20809 39383 20867 39389
rect 20898 39380 20904 39392
rect 20956 39380 20962 39432
rect 26697 39355 26755 39361
rect 19996 39324 20668 39352
rect 1765 39287 1823 39293
rect 1765 39253 1777 39287
rect 1811 39284 1823 39287
rect 3142 39284 3148 39296
rect 1811 39256 3148 39284
rect 1811 39253 1823 39256
rect 1765 39247 1823 39253
rect 3142 39244 3148 39256
rect 3200 39244 3206 39296
rect 17218 39244 17224 39296
rect 17276 39284 17282 39296
rect 17972 39284 18000 39324
rect 17276 39256 18000 39284
rect 17276 39244 17282 39256
rect 18138 39244 18144 39296
rect 18196 39284 18202 39296
rect 18233 39287 18291 39293
rect 18233 39284 18245 39287
rect 18196 39256 18245 39284
rect 18196 39244 18202 39256
rect 18233 39253 18245 39256
rect 18279 39253 18291 39287
rect 18233 39247 18291 39253
rect 19242 39244 19248 39296
rect 19300 39284 19306 39296
rect 19521 39287 19579 39293
rect 19521 39284 19533 39287
rect 19300 39256 19533 39284
rect 19300 39244 19306 39256
rect 19521 39253 19533 39256
rect 19567 39253 19579 39287
rect 19720 39284 19748 39324
rect 20640 39296 20668 39324
rect 26697 39321 26709 39355
rect 26743 39352 26755 39355
rect 27890 39352 27896 39364
rect 26743 39324 27896 39352
rect 26743 39321 26755 39324
rect 26697 39315 26755 39321
rect 27890 39312 27896 39324
rect 27948 39312 27954 39364
rect 19978 39284 19984 39296
rect 19720 39256 19984 39284
rect 19521 39247 19579 39253
rect 19978 39244 19984 39256
rect 20036 39244 20042 39296
rect 20622 39244 20628 39296
rect 20680 39284 20686 39296
rect 20717 39287 20775 39293
rect 20717 39284 20729 39287
rect 20680 39256 20729 39284
rect 20680 39244 20686 39256
rect 20717 39253 20729 39256
rect 20763 39253 20775 39287
rect 20717 39247 20775 39253
rect 1104 39194 29048 39216
rect 1104 39142 7896 39194
rect 7948 39142 7960 39194
rect 8012 39142 8024 39194
rect 8076 39142 8088 39194
rect 8140 39142 8152 39194
rect 8204 39142 14842 39194
rect 14894 39142 14906 39194
rect 14958 39142 14970 39194
rect 15022 39142 15034 39194
rect 15086 39142 15098 39194
rect 15150 39142 21788 39194
rect 21840 39142 21852 39194
rect 21904 39142 21916 39194
rect 21968 39142 21980 39194
rect 22032 39142 22044 39194
rect 22096 39142 28734 39194
rect 28786 39142 28798 39194
rect 28850 39142 28862 39194
rect 28914 39142 28926 39194
rect 28978 39142 28990 39194
rect 29042 39142 29048 39194
rect 1104 39120 29048 39142
rect 18598 39040 18604 39092
rect 18656 39080 18662 39092
rect 19061 39083 19119 39089
rect 19061 39080 19073 39083
rect 18656 39052 19073 39080
rect 18656 39040 18662 39052
rect 19061 39049 19073 39052
rect 19107 39049 19119 39083
rect 19061 39043 19119 39049
rect 19168 39052 19472 39080
rect 18046 38972 18052 39024
rect 18104 39012 18110 39024
rect 18325 39015 18383 39021
rect 18325 39012 18337 39015
rect 18104 38984 18337 39012
rect 18104 38972 18110 38984
rect 18325 38981 18337 38984
rect 18371 39012 18383 39015
rect 18690 39012 18696 39024
rect 18371 38984 18696 39012
rect 18371 38981 18383 38984
rect 18325 38975 18383 38981
rect 18690 38972 18696 38984
rect 18748 38972 18754 39024
rect 18230 38944 18236 38956
rect 18191 38916 18236 38944
rect 18230 38904 18236 38916
rect 18288 38944 18294 38956
rect 19168 38944 19196 39052
rect 19444 39021 19472 39052
rect 19794 39040 19800 39092
rect 19852 39080 19858 39092
rect 19981 39083 20039 39089
rect 19981 39080 19993 39083
rect 19852 39052 19993 39080
rect 19852 39040 19858 39052
rect 19981 39049 19993 39052
rect 20027 39049 20039 39083
rect 19981 39043 20039 39049
rect 19229 39015 19287 39021
rect 19229 38981 19241 39015
rect 19275 39012 19287 39015
rect 19429 39015 19487 39021
rect 19275 38984 19380 39012
rect 19275 38981 19287 38984
rect 19229 38975 19287 38981
rect 18288 38916 19196 38944
rect 19352 38944 19380 38984
rect 19429 38981 19441 39015
rect 19475 38981 19487 39015
rect 19429 38975 19487 38981
rect 26421 39015 26479 39021
rect 26421 38981 26433 39015
rect 26467 39012 26479 39015
rect 27801 39015 27859 39021
rect 27801 39012 27813 39015
rect 26467 38984 27813 39012
rect 26467 38981 26479 38984
rect 26421 38975 26479 38981
rect 27801 38981 27813 38984
rect 27847 38981 27859 39015
rect 27801 38975 27859 38981
rect 19610 38944 19616 38956
rect 19352 38916 19616 38944
rect 18288 38904 18294 38916
rect 19610 38904 19616 38916
rect 19668 38944 19674 38956
rect 19889 38947 19947 38953
rect 19889 38944 19901 38947
rect 19668 38916 19901 38944
rect 19668 38904 19674 38916
rect 19889 38913 19901 38916
rect 19935 38913 19947 38947
rect 19889 38907 19947 38913
rect 20073 38947 20131 38953
rect 20073 38913 20085 38947
rect 20119 38944 20131 38947
rect 20898 38944 20904 38956
rect 20119 38916 20904 38944
rect 20119 38913 20131 38916
rect 20073 38907 20131 38913
rect 19904 38876 19932 38907
rect 20438 38876 20444 38888
rect 19904 38848 20444 38876
rect 20438 38836 20444 38848
rect 20496 38836 20502 38888
rect 2133 38811 2191 38817
rect 2133 38777 2145 38811
rect 2179 38808 2191 38811
rect 3418 38808 3424 38820
rect 2179 38780 3424 38808
rect 2179 38777 2191 38780
rect 2133 38771 2191 38777
rect 3418 38768 3424 38780
rect 3476 38768 3482 38820
rect 2777 38743 2835 38749
rect 2777 38709 2789 38743
rect 2823 38740 2835 38743
rect 3970 38740 3976 38752
rect 2823 38712 3976 38740
rect 2823 38709 2835 38712
rect 2777 38703 2835 38709
rect 3970 38700 3976 38712
rect 4028 38700 4034 38752
rect 18782 38700 18788 38752
rect 18840 38740 18846 38752
rect 19245 38743 19303 38749
rect 19245 38740 19257 38743
rect 18840 38712 19257 38740
rect 18840 38700 18846 38712
rect 19245 38709 19257 38712
rect 19291 38740 19303 38743
rect 20548 38740 20576 38916
rect 20898 38904 20904 38916
rect 20956 38904 20962 38956
rect 26605 38947 26663 38953
rect 26605 38913 26617 38947
rect 26651 38944 26663 38947
rect 27522 38944 27528 38956
rect 26651 38916 27528 38944
rect 26651 38913 26663 38916
rect 26605 38907 26663 38913
rect 27522 38904 27528 38916
rect 27580 38904 27586 38956
rect 27706 38904 27712 38956
rect 27764 38944 27770 38956
rect 28626 38944 28632 38956
rect 27764 38916 28632 38944
rect 27764 38904 27770 38916
rect 28626 38904 28632 38916
rect 28684 38904 28690 38956
rect 22005 38879 22063 38885
rect 22005 38845 22017 38879
rect 22051 38845 22063 38879
rect 22186 38876 22192 38888
rect 22147 38848 22192 38876
rect 22005 38839 22063 38845
rect 22020 38808 22048 38839
rect 22186 38836 22192 38848
rect 22244 38836 22250 38888
rect 23474 38876 23480 38888
rect 23435 38848 23480 38876
rect 23474 38836 23480 38848
rect 23532 38836 23538 38888
rect 26142 38876 26148 38888
rect 26103 38848 26148 38876
rect 26142 38836 26148 38848
rect 26200 38836 26206 38888
rect 23106 38808 23112 38820
rect 22020 38780 23112 38808
rect 23106 38768 23112 38780
rect 23164 38768 23170 38820
rect 19291 38712 20576 38740
rect 19291 38709 19303 38712
rect 19245 38703 19303 38709
rect 1104 38650 28888 38672
rect 1104 38598 4423 38650
rect 4475 38598 4487 38650
rect 4539 38598 4551 38650
rect 4603 38598 4615 38650
rect 4667 38598 4679 38650
rect 4731 38598 11369 38650
rect 11421 38598 11433 38650
rect 11485 38598 11497 38650
rect 11549 38598 11561 38650
rect 11613 38598 11625 38650
rect 11677 38598 18315 38650
rect 18367 38598 18379 38650
rect 18431 38598 18443 38650
rect 18495 38598 18507 38650
rect 18559 38598 18571 38650
rect 18623 38598 25261 38650
rect 25313 38598 25325 38650
rect 25377 38598 25389 38650
rect 25441 38598 25453 38650
rect 25505 38598 25517 38650
rect 25569 38598 28888 38650
rect 1104 38576 28888 38598
rect 15286 38496 15292 38548
rect 15344 38536 15350 38548
rect 17681 38539 17739 38545
rect 17681 38536 17693 38539
rect 15344 38508 17693 38536
rect 15344 38496 15350 38508
rect 16114 38468 16120 38480
rect 15120 38440 16120 38468
rect 15120 38351 15148 38440
rect 16114 38428 16120 38440
rect 16172 38428 16178 38480
rect 15470 38400 15476 38412
rect 15431 38372 15476 38400
rect 15470 38360 15476 38372
rect 15528 38360 15534 38412
rect 15838 38360 15844 38412
rect 15896 38400 15902 38412
rect 15896 38372 16252 38400
rect 15896 38360 15902 38372
rect 15100 38345 15158 38351
rect 1670 38332 1676 38344
rect 1631 38304 1676 38332
rect 1670 38292 1676 38304
rect 1728 38292 1734 38344
rect 2961 38335 3019 38341
rect 2961 38301 2973 38335
rect 3007 38332 3019 38335
rect 5534 38332 5540 38344
rect 3007 38304 5540 38332
rect 3007 38301 3019 38304
rect 2961 38295 3019 38301
rect 5534 38292 5540 38304
rect 5592 38292 5598 38344
rect 15100 38311 15112 38345
rect 15146 38311 15158 38345
rect 15100 38305 15158 38311
rect 15197 38335 15255 38341
rect 15197 38301 15209 38335
rect 15243 38332 15255 38335
rect 15856 38332 15884 38360
rect 16114 38332 16120 38344
rect 15243 38304 15884 38332
rect 16075 38304 16120 38332
rect 15243 38301 15255 38304
rect 15197 38295 15255 38301
rect 16114 38292 16120 38304
rect 16172 38292 16178 38344
rect 16224 38341 16252 38372
rect 16316 38341 16344 38508
rect 17681 38505 17693 38508
rect 17727 38505 17739 38539
rect 17681 38499 17739 38505
rect 21361 38539 21419 38545
rect 21361 38505 21373 38539
rect 21407 38536 21419 38539
rect 22186 38536 22192 38548
rect 21407 38508 22192 38536
rect 21407 38505 21419 38508
rect 21361 38499 21419 38505
rect 22186 38496 22192 38508
rect 22244 38496 22250 38548
rect 27706 38400 27712 38412
rect 26206 38372 27712 38400
rect 16209 38335 16267 38341
rect 16209 38301 16221 38335
rect 16255 38301 16267 38335
rect 16209 38295 16267 38301
rect 16301 38335 16359 38341
rect 16301 38301 16313 38335
rect 16347 38301 16359 38335
rect 16301 38295 16359 38301
rect 16485 38335 16543 38341
rect 16485 38301 16497 38335
rect 16531 38332 16543 38335
rect 17310 38332 17316 38344
rect 16531 38304 17316 38332
rect 16531 38301 16543 38304
rect 16485 38295 16543 38301
rect 15286 38264 15292 38276
rect 15247 38236 15292 38264
rect 15286 38224 15292 38236
rect 15344 38224 15350 38276
rect 15473 38267 15531 38273
rect 15473 38233 15485 38267
rect 15519 38264 15531 38267
rect 16500 38264 16528 38295
rect 17310 38292 17316 38304
rect 17368 38292 17374 38344
rect 17405 38335 17463 38341
rect 17405 38301 17417 38335
rect 17451 38301 17463 38335
rect 17405 38295 17463 38301
rect 17497 38335 17555 38341
rect 17497 38301 17509 38335
rect 17543 38301 17555 38335
rect 17497 38295 17555 38301
rect 15519 38236 16528 38264
rect 15519 38233 15531 38236
rect 15473 38227 15531 38233
rect 2869 38199 2927 38205
rect 2869 38165 2881 38199
rect 2915 38196 2927 38199
rect 3234 38196 3240 38208
rect 2915 38168 3240 38196
rect 2915 38165 2927 38168
rect 2869 38159 2927 38165
rect 3234 38156 3240 38168
rect 3292 38156 3298 38208
rect 15933 38199 15991 38205
rect 15933 38165 15945 38199
rect 15979 38196 15991 38199
rect 16022 38196 16028 38208
rect 15979 38168 16028 38196
rect 15979 38165 15991 38168
rect 15933 38159 15991 38165
rect 16022 38156 16028 38168
rect 16080 38156 16086 38208
rect 17126 38156 17132 38208
rect 17184 38196 17190 38208
rect 17221 38199 17279 38205
rect 17221 38196 17233 38199
rect 17184 38168 17233 38196
rect 17184 38156 17190 38168
rect 17221 38165 17233 38168
rect 17267 38165 17279 38199
rect 17420 38196 17448 38295
rect 17512 38264 17540 38295
rect 17586 38292 17592 38344
rect 17644 38332 17650 38344
rect 17773 38335 17831 38341
rect 17773 38332 17785 38335
rect 17644 38304 17785 38332
rect 17644 38292 17650 38304
rect 17773 38301 17785 38304
rect 17819 38301 17831 38335
rect 17773 38295 17831 38301
rect 17954 38292 17960 38344
rect 18012 38332 18018 38344
rect 18233 38335 18291 38341
rect 18233 38332 18245 38335
rect 18012 38304 18245 38332
rect 18012 38292 18018 38304
rect 18233 38301 18245 38304
rect 18279 38301 18291 38335
rect 18233 38295 18291 38301
rect 21269 38335 21327 38341
rect 21269 38301 21281 38335
rect 21315 38332 21327 38335
rect 21634 38332 21640 38344
rect 21315 38304 21640 38332
rect 21315 38301 21327 38304
rect 21269 38295 21327 38301
rect 21634 38292 21640 38304
rect 21692 38332 21698 38344
rect 26206 38332 26234 38372
rect 27706 38360 27712 38372
rect 27764 38360 27770 38412
rect 28258 38400 28264 38412
rect 28219 38372 28264 38400
rect 28258 38360 28264 38372
rect 28316 38360 28322 38412
rect 26510 38332 26516 38344
rect 21692 38304 26234 38332
rect 26471 38304 26516 38332
rect 21692 38292 21698 38304
rect 26510 38292 26516 38304
rect 26568 38292 26574 38344
rect 18046 38264 18052 38276
rect 17512 38236 18052 38264
rect 18046 38224 18052 38236
rect 18104 38224 18110 38276
rect 26694 38264 26700 38276
rect 26655 38236 26700 38264
rect 26694 38224 26700 38236
rect 26752 38224 26758 38276
rect 17954 38196 17960 38208
rect 17420 38168 17960 38196
rect 17221 38159 17279 38165
rect 17954 38156 17960 38168
rect 18012 38156 18018 38208
rect 18325 38199 18383 38205
rect 18325 38165 18337 38199
rect 18371 38196 18383 38199
rect 18414 38196 18420 38208
rect 18371 38168 18420 38196
rect 18371 38165 18383 38168
rect 18325 38159 18383 38165
rect 18414 38156 18420 38168
rect 18472 38156 18478 38208
rect 1104 38106 29048 38128
rect 1104 38054 7896 38106
rect 7948 38054 7960 38106
rect 8012 38054 8024 38106
rect 8076 38054 8088 38106
rect 8140 38054 8152 38106
rect 8204 38054 14842 38106
rect 14894 38054 14906 38106
rect 14958 38054 14970 38106
rect 15022 38054 15034 38106
rect 15086 38054 15098 38106
rect 15150 38054 21788 38106
rect 21840 38054 21852 38106
rect 21904 38054 21916 38106
rect 21968 38054 21980 38106
rect 22032 38054 22044 38106
rect 22096 38054 28734 38106
rect 28786 38054 28798 38106
rect 28850 38054 28862 38106
rect 28914 38054 28926 38106
rect 28978 38054 28990 38106
rect 29042 38054 29048 38106
rect 1104 38032 29048 38054
rect 15470 37952 15476 38004
rect 15528 37992 15534 38004
rect 27890 37992 27896 38004
rect 15528 37964 17172 37992
rect 27851 37964 27896 37992
rect 15528 37952 15534 37964
rect 17144 37933 17172 37964
rect 27890 37952 27896 37964
rect 27948 37952 27954 38004
rect 3789 37927 3847 37933
rect 3789 37893 3801 37927
rect 3835 37924 3847 37927
rect 4525 37927 4583 37933
rect 4525 37924 4537 37927
rect 3835 37896 4537 37924
rect 3835 37893 3847 37896
rect 3789 37887 3847 37893
rect 4525 37893 4537 37896
rect 4571 37893 4583 37927
rect 4525 37887 4583 37893
rect 16301 37927 16359 37933
rect 16301 37893 16313 37927
rect 16347 37924 16359 37927
rect 16991 37927 17049 37933
rect 16991 37924 17003 37927
rect 16347 37896 17003 37924
rect 16347 37893 16359 37896
rect 16301 37887 16359 37893
rect 16991 37893 17003 37896
rect 17037 37893 17049 37927
rect 16991 37887 17049 37893
rect 17129 37927 17187 37933
rect 17129 37893 17141 37927
rect 17175 37893 17187 37927
rect 17129 37887 17187 37893
rect 17221 37927 17279 37933
rect 17221 37893 17233 37927
rect 17267 37924 17279 37927
rect 19797 37927 19855 37933
rect 19797 37924 19809 37927
rect 17267 37896 19809 37924
rect 17267 37893 17279 37896
rect 17221 37887 17279 37893
rect 19797 37893 19809 37896
rect 19843 37893 19855 37927
rect 19797 37887 19855 37893
rect 3970 37816 3976 37868
rect 4028 37856 4034 37868
rect 4617 37859 4675 37865
rect 4028 37828 4073 37856
rect 4028 37816 4034 37828
rect 4617 37825 4629 37859
rect 4663 37856 4675 37859
rect 4890 37856 4896 37868
rect 4663 37828 4896 37856
rect 4663 37825 4675 37828
rect 4617 37819 4675 37825
rect 4890 37816 4896 37828
rect 4948 37816 4954 37868
rect 16022 37856 16028 37868
rect 15983 37828 16028 37856
rect 16022 37816 16028 37828
rect 16080 37816 16086 37868
rect 16390 37816 16396 37868
rect 16448 37856 16454 37868
rect 16853 37859 16911 37865
rect 16853 37856 16865 37859
rect 16448 37828 16865 37856
rect 16448 37816 16454 37828
rect 16853 37825 16865 37828
rect 16899 37825 16911 37859
rect 16853 37819 16911 37825
rect 2774 37788 2780 37800
rect 2735 37760 2780 37788
rect 2774 37748 2780 37760
rect 2832 37748 2838 37800
rect 16301 37791 16359 37797
rect 16301 37757 16313 37791
rect 16347 37788 16359 37791
rect 16574 37788 16580 37800
rect 16347 37760 16580 37788
rect 16347 37757 16359 37760
rect 16301 37751 16359 37757
rect 16574 37748 16580 37760
rect 16632 37748 16638 37800
rect 16868 37788 16896 37819
rect 17310 37816 17316 37868
rect 17368 37856 17374 37868
rect 18230 37856 18236 37868
rect 17368 37828 17413 37856
rect 18191 37828 18236 37856
rect 17368 37816 17374 37828
rect 18230 37816 18236 37828
rect 18288 37816 18294 37868
rect 18414 37856 18420 37868
rect 18375 37828 18420 37856
rect 18414 37816 18420 37828
rect 18472 37816 18478 37868
rect 18601 37859 18659 37865
rect 18601 37825 18613 37859
rect 18647 37856 18659 37859
rect 18690 37856 18696 37868
rect 18647 37828 18696 37856
rect 18647 37825 18659 37828
rect 18601 37819 18659 37825
rect 18690 37816 18696 37828
rect 18748 37816 18754 37868
rect 18785 37859 18843 37865
rect 18785 37825 18797 37859
rect 18831 37825 18843 37859
rect 19518 37856 19524 37868
rect 19479 37828 19524 37856
rect 18785 37819 18843 37825
rect 16868 37760 18460 37788
rect 16117 37723 16175 37729
rect 16117 37689 16129 37723
rect 16163 37720 16175 37723
rect 17126 37720 17132 37732
rect 16163 37692 17132 37720
rect 16163 37689 16175 37692
rect 16117 37683 16175 37689
rect 17126 37680 17132 37692
rect 17184 37680 17190 37732
rect 18432 37720 18460 37760
rect 18506 37748 18512 37800
rect 18564 37788 18570 37800
rect 18564 37760 18609 37788
rect 18564 37748 18570 37760
rect 18800 37720 18828 37819
rect 19518 37816 19524 37828
rect 19576 37816 19582 37868
rect 26510 37816 26516 37868
rect 26568 37856 26574 37868
rect 27157 37859 27215 37865
rect 27157 37856 27169 37859
rect 26568 37828 27169 37856
rect 26568 37816 26574 37828
rect 27157 37825 27169 37828
rect 27203 37825 27215 37859
rect 27798 37856 27804 37868
rect 27759 37828 27804 37856
rect 27157 37819 27215 37825
rect 27798 37816 27804 37828
rect 27856 37816 27862 37868
rect 19797 37791 19855 37797
rect 19797 37757 19809 37791
rect 19843 37788 19855 37791
rect 20070 37788 20076 37800
rect 19843 37760 20076 37788
rect 19843 37757 19855 37760
rect 19797 37751 19855 37757
rect 20070 37748 20076 37760
rect 20128 37748 20134 37800
rect 18432 37692 18828 37720
rect 16942 37612 16948 37664
rect 17000 37652 17006 37664
rect 17497 37655 17555 37661
rect 17497 37652 17509 37655
rect 17000 37624 17509 37652
rect 17000 37612 17006 37624
rect 17497 37621 17509 37624
rect 17543 37621 17555 37655
rect 17497 37615 17555 37621
rect 17586 37612 17592 37664
rect 17644 37652 17650 37664
rect 18049 37655 18107 37661
rect 18049 37652 18061 37655
rect 17644 37624 18061 37652
rect 17644 37612 17650 37624
rect 18049 37621 18061 37624
rect 18095 37621 18107 37655
rect 18049 37615 18107 37621
rect 18230 37612 18236 37664
rect 18288 37652 18294 37664
rect 19150 37652 19156 37664
rect 18288 37624 19156 37652
rect 18288 37612 18294 37624
rect 19150 37612 19156 37624
rect 19208 37612 19214 37664
rect 19610 37652 19616 37664
rect 19571 37624 19616 37652
rect 19610 37612 19616 37624
rect 19668 37612 19674 37664
rect 1104 37562 28888 37584
rect 1104 37510 4423 37562
rect 4475 37510 4487 37562
rect 4539 37510 4551 37562
rect 4603 37510 4615 37562
rect 4667 37510 4679 37562
rect 4731 37510 11369 37562
rect 11421 37510 11433 37562
rect 11485 37510 11497 37562
rect 11549 37510 11561 37562
rect 11613 37510 11625 37562
rect 11677 37510 18315 37562
rect 18367 37510 18379 37562
rect 18431 37510 18443 37562
rect 18495 37510 18507 37562
rect 18559 37510 18571 37562
rect 18623 37510 25261 37562
rect 25313 37510 25325 37562
rect 25377 37510 25389 37562
rect 25441 37510 25453 37562
rect 25505 37510 25517 37562
rect 25569 37510 28888 37562
rect 1104 37488 28888 37510
rect 17126 37448 17132 37460
rect 17087 37420 17132 37448
rect 17126 37408 17132 37420
rect 17184 37408 17190 37460
rect 17310 37448 17316 37460
rect 17271 37420 17316 37448
rect 17310 37408 17316 37420
rect 17368 37408 17374 37460
rect 17420 37420 18552 37448
rect 16206 37380 16212 37392
rect 15488 37352 16212 37380
rect 15488 37324 15516 37352
rect 16206 37340 16212 37352
rect 16264 37380 16270 37392
rect 17420 37380 17448 37420
rect 18524 37380 18552 37420
rect 18690 37408 18696 37460
rect 18748 37448 18754 37460
rect 19521 37451 19579 37457
rect 19521 37448 19533 37451
rect 18748 37420 19533 37448
rect 18748 37408 18754 37420
rect 19521 37417 19533 37420
rect 19567 37417 19579 37451
rect 20070 37448 20076 37460
rect 20031 37420 20076 37448
rect 19521 37411 19579 37417
rect 20070 37408 20076 37420
rect 20128 37408 20134 37460
rect 20438 37408 20444 37460
rect 20496 37448 20502 37460
rect 20714 37448 20720 37460
rect 20496 37420 20720 37448
rect 20496 37408 20502 37420
rect 20714 37408 20720 37420
rect 20772 37408 20778 37460
rect 24762 37380 24768 37392
rect 16264 37352 17448 37380
rect 17512 37352 18184 37380
rect 18524 37352 23520 37380
rect 24723 37352 24768 37380
rect 16264 37340 16270 37352
rect 3234 37312 3240 37324
rect 3195 37284 3240 37312
rect 3234 37272 3240 37284
rect 3292 37272 3298 37324
rect 15470 37312 15476 37324
rect 15383 37284 15476 37312
rect 15470 37272 15476 37284
rect 15528 37272 15534 37324
rect 1578 37244 1584 37256
rect 1539 37216 1584 37244
rect 1578 37204 1584 37216
rect 1636 37204 1642 37256
rect 3418 37204 3424 37256
rect 3476 37244 3482 37256
rect 3973 37247 4031 37253
rect 3476 37216 3521 37244
rect 3476 37204 3482 37216
rect 3973 37213 3985 37247
rect 4019 37213 4031 37247
rect 17512 37244 17540 37352
rect 18156 37312 18184 37352
rect 20530 37312 20536 37324
rect 18156 37284 19334 37312
rect 3973 37207 4031 37213
rect 6886 37216 17540 37244
rect 3142 37136 3148 37188
rect 3200 37176 3206 37188
rect 3988 37176 4016 37207
rect 4154 37176 4160 37188
rect 3200 37148 4016 37176
rect 4115 37148 4160 37176
rect 3200 37136 3206 37148
rect 4154 37136 4160 37148
rect 4212 37136 4218 37188
rect 5813 37179 5871 37185
rect 5813 37145 5825 37179
rect 5859 37176 5871 37179
rect 6886 37176 6914 37216
rect 18138 37204 18144 37256
rect 18196 37253 18202 37256
rect 18322 37253 18328 37256
rect 18196 37244 18205 37253
rect 18319 37244 18328 37253
rect 18196 37216 18241 37244
rect 18283 37216 18328 37244
rect 18196 37207 18205 37216
rect 18319 37207 18328 37216
rect 18196 37204 18202 37207
rect 18322 37204 18328 37207
rect 18380 37204 18386 37256
rect 5859 37148 6914 37176
rect 15657 37179 15715 37185
rect 5859 37145 5871 37148
rect 5813 37139 5871 37145
rect 15657 37145 15669 37179
rect 15703 37176 15715 37179
rect 16114 37176 16120 37188
rect 15703 37148 16120 37176
rect 15703 37145 15715 37148
rect 15657 37139 15715 37145
rect 16114 37136 16120 37148
rect 16172 37136 16178 37188
rect 16574 37136 16580 37188
rect 16632 37176 16638 37188
rect 16945 37179 17003 37185
rect 16945 37176 16957 37179
rect 16632 37148 16957 37176
rect 16632 37136 16638 37148
rect 16945 37145 16957 37148
rect 16991 37145 17003 37179
rect 16945 37139 17003 37145
rect 17161 37179 17219 37185
rect 17161 37145 17173 37179
rect 17207 37176 17219 37179
rect 17586 37176 17592 37188
rect 17207 37148 17592 37176
rect 17207 37145 17219 37148
rect 17161 37139 17219 37145
rect 17586 37136 17592 37148
rect 17644 37136 17650 37188
rect 19306 37176 19334 37284
rect 19628 37284 20536 37312
rect 19628 37253 19656 37284
rect 20530 37272 20536 37284
rect 20588 37272 20594 37324
rect 21177 37315 21235 37321
rect 21177 37281 21189 37315
rect 21223 37312 21235 37315
rect 22370 37312 22376 37324
rect 21223 37284 22376 37312
rect 21223 37281 21235 37284
rect 21177 37275 21235 37281
rect 22370 37272 22376 37284
rect 22428 37272 22434 37324
rect 23492 37321 23520 37352
rect 24762 37340 24768 37352
rect 24820 37340 24826 37392
rect 26050 37340 26056 37392
rect 26108 37380 26114 37392
rect 26108 37352 26372 37380
rect 26108 37340 26114 37352
rect 23477 37315 23535 37321
rect 23477 37281 23489 37315
rect 23523 37312 23535 37315
rect 26234 37312 26240 37324
rect 23523 37284 26240 37312
rect 23523 37281 23535 37284
rect 23477 37275 23535 37281
rect 26234 37272 26240 37284
rect 26292 37272 26298 37324
rect 26344 37321 26372 37352
rect 26329 37315 26387 37321
rect 26329 37281 26341 37315
rect 26375 37281 26387 37315
rect 26329 37275 26387 37281
rect 19613 37247 19671 37253
rect 19613 37213 19625 37247
rect 19659 37213 19671 37247
rect 19613 37207 19671 37213
rect 20162 37204 20168 37256
rect 20220 37244 20226 37256
rect 20257 37247 20315 37253
rect 20257 37244 20269 37247
rect 20220 37216 20269 37244
rect 20220 37204 20226 37216
rect 20257 37213 20269 37216
rect 20303 37213 20315 37247
rect 20257 37207 20315 37213
rect 20349 37247 20407 37253
rect 20349 37213 20361 37247
rect 20395 37244 20407 37247
rect 20438 37244 20444 37256
rect 20395 37216 20444 37244
rect 20395 37213 20407 37216
rect 20349 37207 20407 37213
rect 20438 37204 20444 37216
rect 20496 37204 20502 37256
rect 20622 37244 20628 37256
rect 20583 37216 20628 37244
rect 20622 37204 20628 37216
rect 20680 37204 20686 37256
rect 20806 37204 20812 37256
rect 20864 37244 20870 37256
rect 21085 37247 21143 37253
rect 21085 37244 21097 37247
rect 20864 37216 21097 37244
rect 20864 37204 20870 37216
rect 21085 37213 21097 37216
rect 21131 37213 21143 37247
rect 21085 37207 21143 37213
rect 21269 37247 21327 37253
rect 21269 37213 21281 37247
rect 21315 37244 21327 37247
rect 21450 37244 21456 37256
rect 21315 37216 21456 37244
rect 21315 37213 21327 37216
rect 21269 37207 21327 37213
rect 21450 37204 21456 37216
rect 21508 37204 21514 37256
rect 23385 37247 23443 37253
rect 23385 37213 23397 37247
rect 23431 37244 23443 37247
rect 23750 37244 23756 37256
rect 23431 37216 23756 37244
rect 23431 37213 23443 37216
rect 23385 37207 23443 37213
rect 23750 37204 23756 37216
rect 23808 37204 23814 37256
rect 24486 37204 24492 37256
rect 24544 37244 24550 37256
rect 24581 37247 24639 37253
rect 24581 37244 24593 37247
rect 24544 37216 24593 37244
rect 24544 37204 24550 37216
rect 24581 37213 24593 37216
rect 24627 37213 24639 37247
rect 24581 37207 24639 37213
rect 24762 37204 24768 37256
rect 24820 37244 24826 37256
rect 25869 37247 25927 37253
rect 25869 37244 25881 37247
rect 24820 37216 25881 37244
rect 24820 37204 24826 37216
rect 25869 37213 25881 37216
rect 25915 37213 25927 37247
rect 28350 37244 28356 37256
rect 28311 37216 28356 37244
rect 25869 37207 25927 37213
rect 28350 37204 28356 37216
rect 28408 37204 28414 37256
rect 26050 37176 26056 37188
rect 19306 37148 23428 37176
rect 26011 37148 26056 37176
rect 6730 37068 6736 37120
rect 6788 37108 6794 37120
rect 15565 37111 15623 37117
rect 15565 37108 15577 37111
rect 6788 37080 15577 37108
rect 6788 37068 6794 37080
rect 15565 37077 15577 37080
rect 15611 37077 15623 37111
rect 16022 37108 16028 37120
rect 15983 37080 16028 37108
rect 15565 37071 15623 37077
rect 16022 37068 16028 37080
rect 16080 37068 16086 37120
rect 18230 37068 18236 37120
rect 18288 37108 18294 37120
rect 18288 37080 18333 37108
rect 18288 37068 18294 37080
rect 19058 37068 19064 37120
rect 19116 37108 19122 37120
rect 21450 37108 21456 37120
rect 19116 37080 21456 37108
rect 19116 37068 19122 37080
rect 21450 37068 21456 37080
rect 21508 37068 21514 37120
rect 22738 37068 22744 37120
rect 22796 37108 22802 37120
rect 22925 37111 22983 37117
rect 22925 37108 22937 37111
rect 22796 37080 22937 37108
rect 22796 37068 22802 37080
rect 22925 37077 22937 37080
rect 22971 37077 22983 37111
rect 23290 37108 23296 37120
rect 23251 37080 23296 37108
rect 22925 37071 22983 37077
rect 23290 37068 23296 37080
rect 23348 37068 23354 37120
rect 23400 37108 23428 37148
rect 26050 37136 26056 37148
rect 26108 37136 26114 37188
rect 26326 37108 26332 37120
rect 23400 37080 26332 37108
rect 26326 37068 26332 37080
rect 26384 37068 26390 37120
rect 28166 37108 28172 37120
rect 28127 37080 28172 37108
rect 28166 37068 28172 37080
rect 28224 37068 28230 37120
rect 1104 37018 29048 37040
rect 1104 36966 7896 37018
rect 7948 36966 7960 37018
rect 8012 36966 8024 37018
rect 8076 36966 8088 37018
rect 8140 36966 8152 37018
rect 8204 36966 14842 37018
rect 14894 36966 14906 37018
rect 14958 36966 14970 37018
rect 15022 36966 15034 37018
rect 15086 36966 15098 37018
rect 15150 36966 21788 37018
rect 21840 36966 21852 37018
rect 21904 36966 21916 37018
rect 21968 36966 21980 37018
rect 22032 36966 22044 37018
rect 22096 36966 28734 37018
rect 28786 36966 28798 37018
rect 28850 36966 28862 37018
rect 28914 36966 28926 37018
rect 28978 36966 28990 37018
rect 29042 36966 29048 37018
rect 1104 36944 29048 36966
rect 4154 36864 4160 36916
rect 4212 36904 4218 36916
rect 5261 36907 5319 36913
rect 5261 36904 5273 36907
rect 4212 36876 5273 36904
rect 4212 36864 4218 36876
rect 5261 36873 5273 36876
rect 5307 36873 5319 36907
rect 5261 36867 5319 36873
rect 15933 36907 15991 36913
rect 15933 36873 15945 36907
rect 15979 36904 15991 36907
rect 17954 36904 17960 36916
rect 15979 36876 17960 36904
rect 15979 36873 15991 36876
rect 15933 36867 15991 36873
rect 17954 36864 17960 36876
rect 18012 36864 18018 36916
rect 19978 36864 19984 36916
rect 20036 36904 20042 36916
rect 20622 36904 20628 36916
rect 20036 36876 20628 36904
rect 20036 36864 20042 36876
rect 20622 36864 20628 36876
rect 20680 36864 20686 36916
rect 20806 36904 20812 36916
rect 20767 36876 20812 36904
rect 20806 36864 20812 36876
rect 20864 36864 20870 36916
rect 23474 36864 23480 36916
rect 23532 36904 23538 36916
rect 23934 36904 23940 36916
rect 23532 36876 23940 36904
rect 23532 36864 23538 36876
rect 23934 36864 23940 36876
rect 23992 36864 23998 36916
rect 25961 36907 26019 36913
rect 25961 36873 25973 36907
rect 26007 36904 26019 36907
rect 26050 36904 26056 36916
rect 26007 36876 26056 36904
rect 26007 36873 26019 36876
rect 25961 36867 26019 36873
rect 26050 36864 26056 36876
rect 26108 36864 26114 36916
rect 26694 36864 26700 36916
rect 26752 36904 26758 36916
rect 27249 36907 27307 36913
rect 27249 36904 27261 36907
rect 26752 36876 27261 36904
rect 26752 36864 26758 36876
rect 27249 36873 27261 36876
rect 27295 36873 27307 36907
rect 27249 36867 27307 36873
rect 3142 36796 3148 36848
rect 3200 36836 3206 36848
rect 3237 36839 3295 36845
rect 3237 36836 3249 36839
rect 3200 36808 3249 36836
rect 3200 36796 3206 36808
rect 3237 36805 3249 36808
rect 3283 36805 3295 36839
rect 3237 36799 3295 36805
rect 3881 36839 3939 36845
rect 3881 36805 3893 36839
rect 3927 36836 3939 36839
rect 4338 36836 4344 36848
rect 3927 36808 4344 36836
rect 3927 36805 3939 36808
rect 3881 36799 3939 36805
rect 4338 36796 4344 36808
rect 4396 36836 4402 36848
rect 4982 36836 4988 36848
rect 4396 36808 4988 36836
rect 4396 36796 4402 36808
rect 4982 36796 4988 36808
rect 5040 36796 5046 36848
rect 20254 36796 20260 36848
rect 20312 36796 20318 36848
rect 20438 36796 20444 36848
rect 20496 36836 20502 36848
rect 21361 36839 21419 36845
rect 21361 36836 21373 36839
rect 20496 36808 21373 36836
rect 20496 36796 20502 36808
rect 21361 36805 21373 36808
rect 21407 36805 21419 36839
rect 21361 36799 21419 36805
rect 21450 36796 21456 36848
rect 21508 36836 21514 36848
rect 22281 36839 22339 36845
rect 22281 36836 22293 36839
rect 21508 36808 22293 36836
rect 21508 36796 21514 36808
rect 22281 36805 22293 36808
rect 22327 36805 22339 36839
rect 27798 36836 27804 36848
rect 22281 36799 22339 36805
rect 26206 36808 27804 36836
rect 1857 36771 1915 36777
rect 1857 36737 1869 36771
rect 1903 36737 1915 36771
rect 1857 36731 1915 36737
rect 1872 36632 1900 36731
rect 4246 36728 4252 36780
rect 4304 36768 4310 36780
rect 4525 36771 4583 36777
rect 4525 36768 4537 36771
rect 4304 36740 4537 36768
rect 4304 36728 4310 36740
rect 4525 36737 4537 36740
rect 4571 36737 4583 36771
rect 4525 36731 4583 36737
rect 5353 36771 5411 36777
rect 5353 36737 5365 36771
rect 5399 36737 5411 36771
rect 5353 36731 5411 36737
rect 2501 36703 2559 36709
rect 2501 36669 2513 36703
rect 2547 36700 2559 36703
rect 2590 36700 2596 36712
rect 2547 36672 2596 36700
rect 2547 36669 2559 36672
rect 2501 36663 2559 36669
rect 2590 36660 2596 36672
rect 2648 36660 2654 36712
rect 4338 36660 4344 36712
rect 4396 36700 4402 36712
rect 5368 36700 5396 36731
rect 5994 36728 6000 36780
rect 6052 36768 6058 36780
rect 19058 36768 19064 36780
rect 6052 36740 12434 36768
rect 19019 36740 19064 36768
rect 6052 36728 6058 36740
rect 4396 36672 5396 36700
rect 12406 36700 12434 36740
rect 19058 36728 19064 36740
rect 19116 36728 19122 36780
rect 19242 36768 19248 36780
rect 19203 36740 19248 36768
rect 19242 36728 19248 36740
rect 19300 36728 19306 36780
rect 20165 36771 20223 36777
rect 20165 36737 20177 36771
rect 20211 36768 20223 36771
rect 20272 36768 20300 36796
rect 20622 36768 20628 36780
rect 20211 36740 20300 36768
rect 20583 36740 20628 36768
rect 20211 36737 20223 36740
rect 20165 36731 20223 36737
rect 20622 36728 20628 36740
rect 20680 36728 20686 36780
rect 21266 36768 21272 36780
rect 21227 36740 21272 36768
rect 21266 36728 21272 36740
rect 21324 36728 21330 36780
rect 22649 36771 22707 36777
rect 22649 36737 22661 36771
rect 22695 36768 22707 36771
rect 23474 36768 23480 36780
rect 22695 36740 23480 36768
rect 22695 36737 22707 36740
rect 22649 36731 22707 36737
rect 23474 36728 23480 36740
rect 23532 36728 23538 36780
rect 25869 36771 25927 36777
rect 25869 36737 25881 36771
rect 25915 36768 25927 36771
rect 25958 36768 25964 36780
rect 25915 36740 25964 36768
rect 25915 36737 25927 36740
rect 25869 36731 25927 36737
rect 25958 36728 25964 36740
rect 26016 36768 26022 36780
rect 26206 36768 26234 36808
rect 27798 36796 27804 36808
rect 27856 36796 27862 36848
rect 26016 36740 26234 36768
rect 26016 36728 26022 36740
rect 26970 36728 26976 36780
rect 27028 36768 27034 36780
rect 27157 36771 27215 36777
rect 27157 36768 27169 36771
rect 27028 36740 27169 36768
rect 27028 36728 27034 36740
rect 27157 36737 27169 36740
rect 27203 36737 27215 36771
rect 27157 36731 27215 36737
rect 16025 36703 16083 36709
rect 16025 36700 16037 36703
rect 12406 36672 16037 36700
rect 4396 36660 4402 36672
rect 16025 36669 16037 36672
rect 16071 36669 16083 36703
rect 16206 36700 16212 36712
rect 16167 36672 16212 36700
rect 16025 36663 16083 36669
rect 16206 36660 16212 36672
rect 16264 36660 16270 36712
rect 20346 36709 20352 36712
rect 20331 36703 20352 36709
rect 20331 36669 20343 36703
rect 20331 36663 20352 36669
rect 20346 36660 20352 36663
rect 20404 36660 20410 36712
rect 20442 36703 20500 36709
rect 20442 36669 20454 36703
rect 20488 36700 20500 36703
rect 20714 36700 20720 36712
rect 20488 36672 20720 36700
rect 20488 36669 20500 36672
rect 20442 36663 20500 36669
rect 20714 36660 20720 36672
rect 20772 36660 20778 36712
rect 4154 36632 4160 36644
rect 1872 36604 4160 36632
rect 4154 36592 4160 36604
rect 4212 36592 4218 36644
rect 20533 36635 20591 36641
rect 20533 36601 20545 36635
rect 20579 36632 20591 36635
rect 20806 36632 20812 36644
rect 20579 36604 20812 36632
rect 20579 36601 20591 36604
rect 20533 36595 20591 36601
rect 20806 36592 20812 36604
rect 20864 36592 20870 36644
rect 1762 36564 1768 36576
rect 1723 36536 1768 36564
rect 1762 36524 1768 36536
rect 1820 36524 1826 36576
rect 15565 36567 15623 36573
rect 15565 36533 15577 36567
rect 15611 36564 15623 36567
rect 15746 36564 15752 36576
rect 15611 36536 15752 36564
rect 15611 36533 15623 36536
rect 15565 36527 15623 36533
rect 15746 36524 15752 36536
rect 15804 36524 15810 36576
rect 19245 36567 19303 36573
rect 19245 36533 19257 36567
rect 19291 36564 19303 36567
rect 19518 36564 19524 36576
rect 19291 36536 19524 36564
rect 19291 36533 19303 36536
rect 19245 36527 19303 36533
rect 19518 36524 19524 36536
rect 19576 36524 19582 36576
rect 27890 36564 27896 36576
rect 27851 36536 27896 36564
rect 27890 36524 27896 36536
rect 27948 36524 27954 36576
rect 1104 36474 28888 36496
rect 1104 36422 4423 36474
rect 4475 36422 4487 36474
rect 4539 36422 4551 36474
rect 4603 36422 4615 36474
rect 4667 36422 4679 36474
rect 4731 36422 11369 36474
rect 11421 36422 11433 36474
rect 11485 36422 11497 36474
rect 11549 36422 11561 36474
rect 11613 36422 11625 36474
rect 11677 36422 18315 36474
rect 18367 36422 18379 36474
rect 18431 36422 18443 36474
rect 18495 36422 18507 36474
rect 18559 36422 18571 36474
rect 18623 36422 25261 36474
rect 25313 36422 25325 36474
rect 25377 36422 25389 36474
rect 25441 36422 25453 36474
rect 25505 36422 25517 36474
rect 25569 36422 28888 36474
rect 1104 36400 28888 36422
rect 4982 36320 4988 36372
rect 5040 36360 5046 36372
rect 5040 36332 6914 36360
rect 5040 36320 5046 36332
rect 1670 36292 1676 36304
rect 1596 36264 1676 36292
rect 1596 36233 1624 36264
rect 1670 36252 1676 36264
rect 1728 36252 1734 36304
rect 6886 36292 6914 36332
rect 19610 36320 19616 36372
rect 19668 36360 19674 36372
rect 19797 36363 19855 36369
rect 19797 36360 19809 36363
rect 19668 36332 19809 36360
rect 19668 36320 19674 36332
rect 19797 36329 19809 36332
rect 19843 36329 19855 36363
rect 20806 36360 20812 36372
rect 20767 36332 20812 36360
rect 19797 36323 19855 36329
rect 20806 36320 20812 36332
rect 20864 36320 20870 36372
rect 27798 36292 27804 36304
rect 6886 36264 27804 36292
rect 27798 36252 27804 36264
rect 27856 36252 27862 36304
rect 1581 36227 1639 36233
rect 1581 36193 1593 36227
rect 1627 36193 1639 36227
rect 1762 36224 1768 36236
rect 1723 36196 1768 36224
rect 1581 36187 1639 36193
rect 1762 36184 1768 36196
rect 1820 36184 1826 36236
rect 2774 36224 2780 36236
rect 2735 36196 2780 36224
rect 2774 36184 2780 36196
rect 2832 36184 2838 36236
rect 18138 36224 18144 36236
rect 16960 36196 18144 36224
rect 4246 36156 4252 36168
rect 4207 36128 4252 36156
rect 4246 36116 4252 36128
rect 4304 36116 4310 36168
rect 16960 36165 16988 36196
rect 18138 36184 18144 36196
rect 18196 36224 18202 36236
rect 19058 36224 19064 36236
rect 18196 36196 19064 36224
rect 18196 36184 18202 36196
rect 19058 36184 19064 36196
rect 19116 36184 19122 36236
rect 20162 36224 20168 36236
rect 19996 36196 20168 36224
rect 16945 36159 17003 36165
rect 16945 36125 16957 36159
rect 16991 36125 17003 36159
rect 16945 36119 17003 36125
rect 17034 36116 17040 36168
rect 17092 36156 17098 36168
rect 19996 36165 20024 36196
rect 20162 36184 20168 36196
rect 20220 36224 20226 36236
rect 23934 36224 23940 36236
rect 20220 36196 23940 36224
rect 20220 36184 20226 36196
rect 23934 36184 23940 36196
rect 23992 36184 23998 36236
rect 26513 36227 26571 36233
rect 26513 36193 26525 36227
rect 26559 36224 26571 36227
rect 27890 36224 27896 36236
rect 26559 36196 27896 36224
rect 26559 36193 26571 36196
rect 26513 36187 26571 36193
rect 27890 36184 27896 36196
rect 27948 36184 27954 36236
rect 17129 36159 17187 36165
rect 17129 36156 17141 36159
rect 17092 36128 17141 36156
rect 17092 36116 17098 36128
rect 17129 36125 17141 36128
rect 17175 36125 17187 36159
rect 17129 36119 17187 36125
rect 19981 36159 20039 36165
rect 19981 36125 19993 36159
rect 20027 36125 20039 36159
rect 19981 36119 20039 36125
rect 20073 36159 20131 36165
rect 20073 36125 20085 36159
rect 20119 36156 20131 36159
rect 20119 36128 20300 36156
rect 20119 36125 20131 36128
rect 20073 36119 20131 36125
rect 4890 36088 4896 36100
rect 4803 36060 4896 36088
rect 4890 36048 4896 36060
rect 4948 36088 4954 36100
rect 12066 36088 12072 36100
rect 4948 36060 12072 36088
rect 4948 36048 4954 36060
rect 12066 36048 12072 36060
rect 12124 36048 12130 36100
rect 19794 36048 19800 36100
rect 19852 36088 19858 36100
rect 20165 36091 20223 36097
rect 20165 36088 20177 36091
rect 19852 36060 20177 36088
rect 19852 36048 19858 36060
rect 20165 36057 20177 36060
rect 20211 36057 20223 36091
rect 20272 36088 20300 36128
rect 20346 36116 20352 36168
rect 20404 36156 20410 36168
rect 20806 36156 20812 36168
rect 20404 36128 20449 36156
rect 20767 36128 20812 36156
rect 20404 36116 20410 36128
rect 20806 36116 20812 36128
rect 20864 36116 20870 36168
rect 20993 36159 21051 36165
rect 20993 36125 21005 36159
rect 21039 36156 21051 36159
rect 21266 36156 21272 36168
rect 21039 36128 21272 36156
rect 21039 36125 21051 36128
rect 20993 36119 21051 36125
rect 21266 36116 21272 36128
rect 21324 36116 21330 36168
rect 22738 36156 22744 36168
rect 22699 36128 22744 36156
rect 22738 36116 22744 36128
rect 22796 36116 22802 36168
rect 28350 36156 28356 36168
rect 28311 36128 28356 36156
rect 28350 36116 28356 36128
rect 28408 36116 28414 36168
rect 20438 36088 20444 36100
rect 20272 36060 20444 36088
rect 20165 36051 20223 36057
rect 20438 36048 20444 36060
rect 20496 36048 20502 36100
rect 22925 36091 22983 36097
rect 22925 36057 22937 36091
rect 22971 36088 22983 36091
rect 23474 36088 23480 36100
rect 22971 36060 23480 36088
rect 22971 36057 22983 36060
rect 22925 36051 22983 36057
rect 23474 36048 23480 36060
rect 23532 36088 23538 36100
rect 24118 36088 24124 36100
rect 23532 36060 24124 36088
rect 23532 36048 23538 36060
rect 24118 36048 24124 36060
rect 24176 36048 24182 36100
rect 26694 36088 26700 36100
rect 26655 36060 26700 36088
rect 26694 36048 26700 36060
rect 26752 36048 26758 36100
rect 17037 36023 17095 36029
rect 17037 35989 17049 36023
rect 17083 36020 17095 36023
rect 17310 36020 17316 36032
rect 17083 35992 17316 36020
rect 17083 35989 17095 35992
rect 17037 35983 17095 35989
rect 17310 35980 17316 35992
rect 17368 35980 17374 36032
rect 23014 35980 23020 36032
rect 23072 36020 23078 36032
rect 23109 36023 23167 36029
rect 23109 36020 23121 36023
rect 23072 35992 23121 36020
rect 23072 35980 23078 35992
rect 23109 35989 23121 35992
rect 23155 35989 23167 36023
rect 23109 35983 23167 35989
rect 1104 35930 29048 35952
rect 1104 35878 7896 35930
rect 7948 35878 7960 35930
rect 8012 35878 8024 35930
rect 8076 35878 8088 35930
rect 8140 35878 8152 35930
rect 8204 35878 14842 35930
rect 14894 35878 14906 35930
rect 14958 35878 14970 35930
rect 15022 35878 15034 35930
rect 15086 35878 15098 35930
rect 15150 35878 21788 35930
rect 21840 35878 21852 35930
rect 21904 35878 21916 35930
rect 21968 35878 21980 35930
rect 22032 35878 22044 35930
rect 22096 35878 28734 35930
rect 28786 35878 28798 35930
rect 28850 35878 28862 35930
rect 28914 35878 28926 35930
rect 28978 35878 28990 35930
rect 29042 35878 29048 35930
rect 1104 35856 29048 35878
rect 12066 35816 12072 35828
rect 11979 35788 12072 35816
rect 2314 35748 2320 35760
rect 2275 35720 2320 35748
rect 2314 35708 2320 35720
rect 2372 35708 2378 35760
rect 2590 35640 2596 35692
rect 2648 35680 2654 35692
rect 3145 35683 3203 35689
rect 3145 35680 3157 35683
rect 2648 35652 3157 35680
rect 2648 35640 2654 35652
rect 3145 35649 3157 35652
rect 3191 35680 3203 35683
rect 3789 35683 3847 35689
rect 3789 35680 3801 35683
rect 3191 35652 3801 35680
rect 3191 35649 3203 35652
rect 3145 35643 3203 35649
rect 3789 35649 3801 35652
rect 3835 35680 3847 35683
rect 4246 35680 4252 35692
rect 3835 35652 4252 35680
rect 3835 35649 3847 35652
rect 3789 35643 3847 35649
rect 4246 35640 4252 35652
rect 4304 35680 4310 35692
rect 11992 35689 12020 35788
rect 12066 35776 12072 35788
rect 12124 35816 12130 35828
rect 12124 35788 26234 35816
rect 12124 35776 12130 35788
rect 12710 35748 12716 35760
rect 12671 35720 12716 35748
rect 12710 35708 12716 35720
rect 12768 35708 12774 35760
rect 18782 35748 18788 35760
rect 18156 35720 18788 35748
rect 5169 35683 5227 35689
rect 5169 35680 5181 35683
rect 4304 35652 5181 35680
rect 4304 35640 4310 35652
rect 5169 35649 5181 35652
rect 5215 35649 5227 35683
rect 5169 35643 5227 35649
rect 11977 35683 12035 35689
rect 11977 35649 11989 35683
rect 12023 35649 12035 35683
rect 15746 35680 15752 35692
rect 15707 35652 15752 35680
rect 11977 35643 12035 35649
rect 15746 35640 15752 35652
rect 15804 35640 15810 35692
rect 18156 35689 18184 35720
rect 18782 35708 18788 35720
rect 18840 35708 18846 35760
rect 26206 35748 26234 35788
rect 26694 35776 26700 35828
rect 26752 35816 26758 35828
rect 27249 35819 27307 35825
rect 27249 35816 27261 35819
rect 26752 35788 27261 35816
rect 26752 35776 26758 35788
rect 27249 35785 27261 35788
rect 27295 35785 27307 35819
rect 27249 35779 27307 35785
rect 26878 35748 26884 35760
rect 26206 35720 26884 35748
rect 26878 35708 26884 35720
rect 26936 35708 26942 35760
rect 15933 35683 15991 35689
rect 15933 35649 15945 35683
rect 15979 35680 15991 35683
rect 16853 35683 16911 35689
rect 16853 35680 16865 35683
rect 15979 35652 16865 35680
rect 15979 35649 15991 35652
rect 15933 35643 15991 35649
rect 16853 35649 16865 35652
rect 16899 35649 16911 35683
rect 16853 35643 16911 35649
rect 18141 35683 18199 35689
rect 18141 35649 18153 35683
rect 18187 35649 18199 35683
rect 18141 35643 18199 35649
rect 18230 35640 18236 35692
rect 18288 35680 18294 35692
rect 18397 35683 18455 35689
rect 18397 35680 18409 35683
rect 18288 35652 18409 35680
rect 18288 35640 18294 35652
rect 18397 35649 18409 35652
rect 18443 35649 18455 35683
rect 23014 35680 23020 35692
rect 22975 35652 23020 35680
rect 18397 35643 18455 35649
rect 23014 35640 23020 35652
rect 23072 35640 23078 35692
rect 26421 35683 26479 35689
rect 26421 35649 26433 35683
rect 26467 35680 26479 35683
rect 27246 35680 27252 35692
rect 26467 35652 27252 35680
rect 26467 35649 26479 35652
rect 26421 35643 26479 35649
rect 27246 35640 27252 35652
rect 27304 35640 27310 35692
rect 27341 35683 27399 35689
rect 27341 35649 27353 35683
rect 27387 35680 27399 35683
rect 28442 35680 28448 35692
rect 27387 35652 28448 35680
rect 27387 35649 27399 35652
rect 27341 35643 27399 35649
rect 28442 35640 28448 35652
rect 28500 35640 28506 35692
rect 4154 35572 4160 35624
rect 4212 35612 4218 35624
rect 4433 35615 4491 35621
rect 4433 35612 4445 35615
rect 4212 35584 4445 35612
rect 4212 35572 4218 35584
rect 4433 35581 4445 35584
rect 4479 35612 4491 35615
rect 4798 35612 4804 35624
rect 4479 35584 4804 35612
rect 4479 35581 4491 35584
rect 4433 35575 4491 35581
rect 4798 35572 4804 35584
rect 4856 35572 4862 35624
rect 5718 35612 5724 35624
rect 5679 35584 5724 35612
rect 5718 35572 5724 35584
rect 5776 35572 5782 35624
rect 15562 35612 15568 35624
rect 15523 35584 15568 35612
rect 15562 35572 15568 35584
rect 15620 35572 15626 35624
rect 25682 35612 25688 35624
rect 25643 35584 25688 35612
rect 25682 35572 25688 35584
rect 25740 35572 25746 35624
rect 19150 35504 19156 35556
rect 19208 35544 19214 35556
rect 19521 35547 19579 35553
rect 19521 35544 19533 35547
rect 19208 35516 19533 35544
rect 19208 35504 19214 35516
rect 19521 35513 19533 35516
rect 19567 35513 19579 35547
rect 19521 35507 19579 35513
rect 17037 35479 17095 35485
rect 17037 35445 17049 35479
rect 17083 35476 17095 35479
rect 17126 35476 17132 35488
rect 17083 35448 17132 35476
rect 17083 35445 17095 35448
rect 17037 35439 17095 35445
rect 17126 35436 17132 35448
rect 17184 35436 17190 35488
rect 22830 35476 22836 35488
rect 22791 35448 22836 35476
rect 22830 35436 22836 35448
rect 22888 35436 22894 35488
rect 24946 35436 24952 35488
rect 25004 35476 25010 35488
rect 25133 35479 25191 35485
rect 25133 35476 25145 35479
rect 25004 35448 25145 35476
rect 25004 35436 25010 35448
rect 25133 35445 25145 35448
rect 25179 35445 25191 35479
rect 25133 35439 25191 35445
rect 26234 35436 26240 35488
rect 26292 35476 26298 35488
rect 27982 35476 27988 35488
rect 26292 35448 26337 35476
rect 27943 35448 27988 35476
rect 26292 35436 26298 35448
rect 27982 35436 27988 35448
rect 28040 35436 28046 35488
rect 1104 35386 28888 35408
rect 1104 35334 4423 35386
rect 4475 35334 4487 35386
rect 4539 35334 4551 35386
rect 4603 35334 4615 35386
rect 4667 35334 4679 35386
rect 4731 35334 11369 35386
rect 11421 35334 11433 35386
rect 11485 35334 11497 35386
rect 11549 35334 11561 35386
rect 11613 35334 11625 35386
rect 11677 35334 18315 35386
rect 18367 35334 18379 35386
rect 18431 35334 18443 35386
rect 18495 35334 18507 35386
rect 18559 35334 18571 35386
rect 18623 35334 25261 35386
rect 25313 35334 25325 35386
rect 25377 35334 25389 35386
rect 25441 35334 25453 35386
rect 25505 35334 25517 35386
rect 25569 35334 28888 35386
rect 1104 35312 28888 35334
rect 12710 35232 12716 35284
rect 12768 35272 12774 35284
rect 12768 35244 17908 35272
rect 12768 35232 12774 35244
rect 17880 35204 17908 35244
rect 17954 35232 17960 35284
rect 18012 35272 18018 35284
rect 18233 35275 18291 35281
rect 18233 35272 18245 35275
rect 18012 35244 18245 35272
rect 18012 35232 18018 35244
rect 18233 35241 18245 35244
rect 18279 35241 18291 35275
rect 20809 35275 20867 35281
rect 18233 35235 18291 35241
rect 18340 35244 20760 35272
rect 18340 35204 18368 35244
rect 17880 35176 18368 35204
rect 20732 35204 20760 35244
rect 20809 35241 20821 35275
rect 20855 35272 20867 35275
rect 20898 35272 20904 35284
rect 20855 35244 20904 35272
rect 20855 35241 20867 35244
rect 20809 35235 20867 35241
rect 20898 35232 20904 35244
rect 20956 35232 20962 35284
rect 21266 35272 21272 35284
rect 21227 35244 21272 35272
rect 21266 35232 21272 35244
rect 21324 35232 21330 35284
rect 28074 35272 28080 35284
rect 21376 35244 28080 35272
rect 21376 35204 21404 35244
rect 28074 35232 28080 35244
rect 28132 35232 28138 35284
rect 20732 35176 21404 35204
rect 2866 35136 2872 35148
rect 2827 35108 2872 35136
rect 2866 35096 2872 35108
rect 2924 35096 2930 35148
rect 4338 35136 4344 35148
rect 4299 35108 4344 35136
rect 4338 35096 4344 35108
rect 4396 35096 4402 35148
rect 1670 35068 1676 35080
rect 1631 35040 1676 35068
rect 1670 35028 1676 35040
rect 1728 35028 1734 35080
rect 2593 35071 2651 35077
rect 2593 35037 2605 35071
rect 2639 35068 2651 35071
rect 4157 35071 4215 35077
rect 4157 35068 4169 35071
rect 2639 35040 4169 35068
rect 2639 35037 2651 35040
rect 2593 35031 2651 35037
rect 4157 35037 4169 35040
rect 4203 35068 4215 35071
rect 4246 35068 4252 35080
rect 4203 35040 4252 35068
rect 4203 35037 4215 35040
rect 4157 35031 4215 35037
rect 4246 35028 4252 35040
rect 4304 35028 4310 35080
rect 17126 35077 17132 35080
rect 16853 35071 16911 35077
rect 16853 35037 16865 35071
rect 16899 35037 16911 35071
rect 17120 35068 17132 35077
rect 17087 35040 17132 35068
rect 16853 35031 16911 35037
rect 17120 35031 17132 35040
rect 4338 34960 4344 35012
rect 4396 35000 4402 35012
rect 14366 35000 14372 35012
rect 4396 34972 14372 35000
rect 4396 34960 4402 34972
rect 14366 34960 14372 34972
rect 14424 34960 14430 35012
rect 16868 35000 16896 35031
rect 17126 35028 17132 35031
rect 17184 35028 17190 35080
rect 18782 35028 18788 35080
rect 18840 35068 18846 35080
rect 19429 35071 19487 35077
rect 19429 35068 19441 35071
rect 18840 35040 19441 35068
rect 18840 35028 18846 35040
rect 19429 35037 19441 35040
rect 19475 35037 19487 35071
rect 19429 35031 19487 35037
rect 19518 35028 19524 35080
rect 19576 35068 19582 35080
rect 19685 35071 19743 35077
rect 19685 35068 19697 35071
rect 19576 35040 19697 35068
rect 19576 35028 19582 35040
rect 19685 35037 19697 35040
rect 19731 35037 19743 35071
rect 22370 35068 22376 35080
rect 22428 35077 22434 35080
rect 22340 35040 22376 35068
rect 19685 35031 19743 35037
rect 22370 35028 22376 35040
rect 22428 35031 22440 35077
rect 22649 35071 22707 35077
rect 22649 35037 22661 35071
rect 22695 35068 22707 35071
rect 26421 35071 26479 35077
rect 22695 35040 23428 35068
rect 22695 35037 22707 35040
rect 22649 35031 22707 35037
rect 22428 35028 22434 35031
rect 17034 35000 17040 35012
rect 16868 34972 17040 35000
rect 17034 34960 17040 34972
rect 17092 35000 17098 35012
rect 18800 35000 18828 35028
rect 23400 35012 23428 35040
rect 26421 35037 26433 35071
rect 26467 35068 26479 35071
rect 28261 35071 28319 35077
rect 28261 35068 28273 35071
rect 26467 35040 28273 35068
rect 26467 35037 26479 35040
rect 26421 35031 26479 35037
rect 28261 35037 28273 35040
rect 28307 35037 28319 35071
rect 28261 35031 28319 35037
rect 17092 34972 18828 35000
rect 17092 34960 17098 34972
rect 20530 34960 20536 35012
rect 20588 35000 20594 35012
rect 20588 34972 22094 35000
rect 20588 34960 20594 34972
rect 22066 34932 22094 34972
rect 23382 34960 23388 35012
rect 23440 35000 23446 35012
rect 26234 35009 26240 35012
rect 26176 35003 26240 35009
rect 26176 35000 26188 35003
rect 23440 34972 25176 35000
rect 26147 34972 26188 35000
rect 23440 34960 23446 34972
rect 25038 34932 25044 34944
rect 22066 34904 25044 34932
rect 25038 34892 25044 34904
rect 25096 34892 25102 34944
rect 25148 34932 25176 34972
rect 26176 34969 26188 34972
rect 26222 34969 26240 35003
rect 26176 34963 26240 34969
rect 26234 34960 26240 34963
rect 26292 34960 26298 35012
rect 26436 34932 26464 35031
rect 28016 35003 28074 35009
rect 28016 34969 28028 35003
rect 28062 35000 28074 35003
rect 28166 35000 28172 35012
rect 28062 34972 28172 35000
rect 28062 34969 28074 34972
rect 28016 34963 28074 34969
rect 28166 34960 28172 34972
rect 28224 34960 28230 35012
rect 26602 34932 26608 34944
rect 25148 34904 26608 34932
rect 26602 34892 26608 34904
rect 26660 34892 26666 34944
rect 26881 34935 26939 34941
rect 26881 34901 26893 34935
rect 26927 34932 26939 34935
rect 27706 34932 27712 34944
rect 26927 34904 27712 34932
rect 26927 34901 26939 34904
rect 26881 34895 26939 34901
rect 27706 34892 27712 34904
rect 27764 34892 27770 34944
rect 1104 34842 29048 34864
rect 1104 34790 7896 34842
rect 7948 34790 7960 34842
rect 8012 34790 8024 34842
rect 8076 34790 8088 34842
rect 8140 34790 8152 34842
rect 8204 34790 14842 34842
rect 14894 34790 14906 34842
rect 14958 34790 14970 34842
rect 15022 34790 15034 34842
rect 15086 34790 15098 34842
rect 15150 34790 21788 34842
rect 21840 34790 21852 34842
rect 21904 34790 21916 34842
rect 21968 34790 21980 34842
rect 22032 34790 22044 34842
rect 22096 34790 28734 34842
rect 28786 34790 28798 34842
rect 28850 34790 28862 34842
rect 28914 34790 28926 34842
rect 28978 34790 28990 34842
rect 29042 34790 29048 34842
rect 1104 34768 29048 34790
rect 15562 34688 15568 34740
rect 15620 34728 15626 34740
rect 15620 34700 17448 34728
rect 15620 34688 15626 34700
rect 7742 34660 7748 34672
rect 5184 34632 7748 34660
rect 1670 34592 1676 34604
rect 1631 34564 1676 34592
rect 1670 34552 1676 34564
rect 1728 34552 1734 34604
rect 4157 34595 4215 34601
rect 4157 34561 4169 34595
rect 4203 34592 4215 34595
rect 4246 34592 4252 34604
rect 4203 34564 4252 34592
rect 4203 34561 4215 34564
rect 4157 34555 4215 34561
rect 4246 34552 4252 34564
rect 4304 34552 4310 34604
rect 5184 34536 5212 34632
rect 7742 34620 7748 34632
rect 7800 34620 7806 34672
rect 15672 34660 15700 34700
rect 15580 34632 15700 34660
rect 15580 34601 15608 34632
rect 15565 34595 15623 34601
rect 15565 34561 15577 34595
rect 15611 34561 15623 34595
rect 15565 34555 15623 34561
rect 15657 34595 15715 34601
rect 15657 34561 15669 34595
rect 15703 34592 15715 34595
rect 16022 34592 16028 34604
rect 15703 34564 16028 34592
rect 15703 34561 15715 34564
rect 15657 34555 15715 34561
rect 16022 34552 16028 34564
rect 16080 34552 16086 34604
rect 17034 34592 17040 34604
rect 16995 34564 17040 34592
rect 17034 34552 17040 34564
rect 17092 34552 17098 34604
rect 17310 34601 17316 34604
rect 17304 34592 17316 34601
rect 17271 34564 17316 34592
rect 17304 34555 17316 34564
rect 17310 34552 17316 34555
rect 17368 34552 17374 34604
rect 17420 34592 17448 34700
rect 17862 34688 17868 34740
rect 17920 34728 17926 34740
rect 18417 34731 18475 34737
rect 18417 34728 18429 34731
rect 17920 34700 18429 34728
rect 17920 34688 17926 34700
rect 18417 34697 18429 34700
rect 18463 34697 18475 34731
rect 18417 34691 18475 34697
rect 20517 34731 20575 34737
rect 20517 34697 20529 34731
rect 20563 34728 20575 34731
rect 21174 34728 21180 34740
rect 20563 34700 21180 34728
rect 20563 34697 20575 34700
rect 20517 34691 20575 34697
rect 21174 34688 21180 34700
rect 21232 34688 21238 34740
rect 23934 34728 23940 34740
rect 23895 34700 23940 34728
rect 23934 34688 23940 34700
rect 23992 34688 23998 34740
rect 24854 34688 24860 34740
rect 24912 34728 24918 34740
rect 25225 34731 25283 34737
rect 25225 34728 25237 34731
rect 24912 34700 25237 34728
rect 24912 34688 24918 34700
rect 25225 34697 25237 34700
rect 25271 34728 25283 34731
rect 25682 34728 25688 34740
rect 25271 34700 25688 34728
rect 25271 34697 25283 34700
rect 25225 34691 25283 34697
rect 25682 34688 25688 34700
rect 25740 34688 25746 34740
rect 20717 34663 20775 34669
rect 20717 34629 20729 34663
rect 20763 34660 20775 34663
rect 21266 34660 21272 34672
rect 20763 34632 21272 34660
rect 20763 34629 20775 34632
rect 20717 34623 20775 34629
rect 21266 34620 21272 34632
rect 21324 34620 21330 34672
rect 22830 34669 22836 34672
rect 22824 34660 22836 34669
rect 22791 34632 22836 34660
rect 22824 34623 22836 34632
rect 22830 34620 22836 34623
rect 22888 34620 22894 34672
rect 26360 34663 26418 34669
rect 26360 34629 26372 34663
rect 26406 34660 26418 34663
rect 27157 34663 27215 34669
rect 27157 34660 27169 34663
rect 26406 34632 27169 34660
rect 26406 34629 26418 34632
rect 26360 34623 26418 34629
rect 27157 34629 27169 34632
rect 27203 34629 27215 34663
rect 27157 34623 27215 34629
rect 20070 34592 20076 34604
rect 17420 34564 20076 34592
rect 20070 34552 20076 34564
rect 20128 34552 20134 34604
rect 26602 34592 26608 34604
rect 26563 34564 26608 34592
rect 26602 34552 26608 34564
rect 26660 34552 26666 34604
rect 27706 34592 27712 34604
rect 27667 34564 27712 34592
rect 27706 34552 27712 34564
rect 27764 34552 27770 34604
rect 1854 34524 1860 34536
rect 1815 34496 1860 34524
rect 1854 34484 1860 34496
rect 1912 34484 1918 34536
rect 2774 34524 2780 34536
rect 2735 34496 2780 34524
rect 2774 34484 2780 34496
rect 2832 34484 2838 34536
rect 4801 34527 4859 34533
rect 4801 34493 4813 34527
rect 4847 34524 4859 34527
rect 5166 34524 5172 34536
rect 4847 34496 5172 34524
rect 4847 34493 4859 34496
rect 4801 34487 4859 34493
rect 5166 34484 5172 34496
rect 5224 34484 5230 34536
rect 5718 34484 5724 34536
rect 5776 34524 5782 34536
rect 8386 34524 8392 34536
rect 5776 34496 8392 34524
rect 5776 34484 5782 34496
rect 8386 34484 8392 34496
rect 8444 34524 8450 34536
rect 12802 34524 12808 34536
rect 8444 34496 12808 34524
rect 8444 34484 8450 34496
rect 12802 34484 12808 34496
rect 12860 34484 12866 34536
rect 20714 34524 20720 34536
rect 20364 34496 20720 34524
rect 20364 34465 20392 34496
rect 20714 34484 20720 34496
rect 20772 34484 20778 34536
rect 22554 34524 22560 34536
rect 22515 34496 22560 34524
rect 22554 34484 22560 34496
rect 22612 34484 22618 34536
rect 27798 34484 27804 34536
rect 27856 34524 27862 34536
rect 28074 34524 28080 34536
rect 27856 34496 28080 34524
rect 27856 34484 27862 34496
rect 28074 34484 28080 34496
rect 28132 34484 28138 34536
rect 20349 34459 20407 34465
rect 20349 34425 20361 34459
rect 20395 34425 20407 34459
rect 20349 34419 20407 34425
rect 15841 34391 15899 34397
rect 15841 34357 15853 34391
rect 15887 34388 15899 34391
rect 16022 34388 16028 34400
rect 15887 34360 16028 34388
rect 15887 34357 15899 34360
rect 15841 34351 15899 34357
rect 16022 34348 16028 34360
rect 16080 34348 16086 34400
rect 20533 34391 20591 34397
rect 20533 34357 20545 34391
rect 20579 34388 20591 34391
rect 20714 34388 20720 34400
rect 20579 34360 20720 34388
rect 20579 34357 20591 34360
rect 20533 34351 20591 34357
rect 20714 34348 20720 34360
rect 20772 34348 20778 34400
rect 1104 34298 28888 34320
rect 1104 34246 4423 34298
rect 4475 34246 4487 34298
rect 4539 34246 4551 34298
rect 4603 34246 4615 34298
rect 4667 34246 4679 34298
rect 4731 34246 11369 34298
rect 11421 34246 11433 34298
rect 11485 34246 11497 34298
rect 11549 34246 11561 34298
rect 11613 34246 11625 34298
rect 11677 34246 18315 34298
rect 18367 34246 18379 34298
rect 18431 34246 18443 34298
rect 18495 34246 18507 34298
rect 18559 34246 18571 34298
rect 18623 34246 25261 34298
rect 25313 34246 25325 34298
rect 25377 34246 25389 34298
rect 25441 34246 25453 34298
rect 25505 34246 25517 34298
rect 25569 34246 28888 34298
rect 1104 34224 28888 34246
rect 1854 34144 1860 34196
rect 1912 34184 1918 34196
rect 2133 34187 2191 34193
rect 2133 34184 2145 34187
rect 1912 34156 2145 34184
rect 1912 34144 1918 34156
rect 2133 34153 2145 34156
rect 2179 34153 2191 34187
rect 2133 34147 2191 34153
rect 20346 34144 20352 34196
rect 20404 34184 20410 34196
rect 20533 34187 20591 34193
rect 20533 34184 20545 34187
rect 20404 34156 20545 34184
rect 20404 34144 20410 34156
rect 20533 34153 20545 34156
rect 20579 34153 20591 34187
rect 20533 34147 20591 34153
rect 23382 34008 23388 34060
rect 23440 34048 23446 34060
rect 24673 34051 24731 34057
rect 24673 34048 24685 34051
rect 23440 34020 24685 34048
rect 23440 34008 23446 34020
rect 24673 34017 24685 34020
rect 24719 34017 24731 34051
rect 27522 34048 27528 34060
rect 27483 34020 27528 34048
rect 24673 34011 24731 34017
rect 27522 34008 27528 34020
rect 27580 34008 27586 34060
rect 27982 34008 27988 34060
rect 28040 34048 28046 34060
rect 28353 34051 28411 34057
rect 28353 34048 28365 34051
rect 28040 34020 28365 34048
rect 28040 34008 28046 34020
rect 28353 34017 28365 34020
rect 28399 34017 28411 34051
rect 28353 34011 28411 34017
rect 2225 33983 2283 33989
rect 2225 33949 2237 33983
rect 2271 33980 2283 33983
rect 2314 33980 2320 33992
rect 2271 33952 2320 33980
rect 2271 33949 2283 33952
rect 2225 33943 2283 33949
rect 2314 33940 2320 33952
rect 2372 33980 2378 33992
rect 2866 33980 2872 33992
rect 2372 33952 2872 33980
rect 2372 33940 2378 33952
rect 2866 33940 2872 33952
rect 2924 33940 2930 33992
rect 4246 33940 4252 33992
rect 4304 33980 4310 33992
rect 4801 33983 4859 33989
rect 4801 33980 4813 33983
rect 4304 33952 4813 33980
rect 4304 33940 4310 33952
rect 4801 33949 4813 33952
rect 4847 33949 4859 33983
rect 16022 33980 16028 33992
rect 15983 33952 16028 33980
rect 4801 33943 4859 33949
rect 16022 33940 16028 33952
rect 16080 33940 16086 33992
rect 20625 33983 20683 33989
rect 20625 33949 20637 33983
rect 20671 33980 20683 33983
rect 20714 33980 20720 33992
rect 20671 33952 20720 33980
rect 20671 33949 20683 33952
rect 20625 33943 20683 33949
rect 20714 33940 20720 33952
rect 20772 33940 20778 33992
rect 21266 33980 21272 33992
rect 21227 33952 21272 33980
rect 21266 33940 21272 33952
rect 21324 33940 21330 33992
rect 23658 33980 23664 33992
rect 23619 33952 23664 33980
rect 23658 33940 23664 33952
rect 23716 33940 23722 33992
rect 23750 33940 23756 33992
rect 23808 33980 23814 33992
rect 23937 33983 23995 33989
rect 23808 33952 23853 33980
rect 23808 33940 23814 33952
rect 23937 33949 23949 33983
rect 23983 33949 23995 33983
rect 23937 33943 23995 33949
rect 24029 33983 24087 33989
rect 24029 33949 24041 33983
rect 24075 33980 24087 33983
rect 24118 33980 24124 33992
rect 24075 33952 24124 33980
rect 24075 33949 24087 33952
rect 24029 33943 24087 33949
rect 4154 33912 4160 33924
rect 4115 33884 4160 33912
rect 4154 33872 4160 33884
rect 4212 33912 4218 33924
rect 5074 33912 5080 33924
rect 4212 33884 5080 33912
rect 4212 33872 4218 33884
rect 5074 33872 5080 33884
rect 5132 33872 5138 33924
rect 21358 33872 21364 33924
rect 21416 33912 21422 33924
rect 21514 33915 21572 33921
rect 21514 33912 21526 33915
rect 21416 33884 21526 33912
rect 21416 33872 21422 33884
rect 21514 33881 21526 33884
rect 21560 33881 21572 33915
rect 23952 33912 23980 33943
rect 24118 33940 24124 33952
rect 24176 33940 24182 33992
rect 24946 33989 24952 33992
rect 24940 33980 24952 33989
rect 24907 33952 24952 33980
rect 24940 33943 24952 33952
rect 24946 33940 24952 33943
rect 25004 33940 25010 33992
rect 25130 33912 25136 33924
rect 21514 33875 21572 33881
rect 22664 33884 23888 33912
rect 23952 33884 25136 33912
rect 16206 33844 16212 33856
rect 16167 33816 16212 33844
rect 16206 33804 16212 33816
rect 16264 33804 16270 33856
rect 20898 33804 20904 33856
rect 20956 33844 20962 33856
rect 22664 33853 22692 33884
rect 22649 33847 22707 33853
rect 22649 33844 22661 33847
rect 20956 33816 22661 33844
rect 20956 33804 20962 33816
rect 22649 33813 22661 33816
rect 22695 33813 22707 33847
rect 22649 33807 22707 33813
rect 23477 33847 23535 33853
rect 23477 33813 23489 33847
rect 23523 33844 23535 33847
rect 23566 33844 23572 33856
rect 23523 33816 23572 33844
rect 23523 33813 23535 33816
rect 23477 33807 23535 33813
rect 23566 33804 23572 33816
rect 23624 33804 23630 33856
rect 23860 33844 23888 33884
rect 25130 33872 25136 33884
rect 25188 33872 25194 33924
rect 28074 33872 28080 33924
rect 28132 33912 28138 33924
rect 28169 33915 28227 33921
rect 28169 33912 28181 33915
rect 28132 33884 28181 33912
rect 28132 33872 28138 33884
rect 28169 33881 28181 33884
rect 28215 33881 28227 33915
rect 28169 33875 28227 33881
rect 25774 33844 25780 33856
rect 23860 33816 25780 33844
rect 25774 33804 25780 33816
rect 25832 33804 25838 33856
rect 25866 33804 25872 33856
rect 25924 33844 25930 33856
rect 26053 33847 26111 33853
rect 26053 33844 26065 33847
rect 25924 33816 26065 33844
rect 25924 33804 25930 33816
rect 26053 33813 26065 33816
rect 26099 33813 26111 33847
rect 26053 33807 26111 33813
rect 1104 33754 29048 33776
rect 1104 33702 7896 33754
rect 7948 33702 7960 33754
rect 8012 33702 8024 33754
rect 8076 33702 8088 33754
rect 8140 33702 8152 33754
rect 8204 33702 14842 33754
rect 14894 33702 14906 33754
rect 14958 33702 14970 33754
rect 15022 33702 15034 33754
rect 15086 33702 15098 33754
rect 15150 33702 21788 33754
rect 21840 33702 21852 33754
rect 21904 33702 21916 33754
rect 21968 33702 21980 33754
rect 22032 33702 22044 33754
rect 22096 33702 28734 33754
rect 28786 33702 28798 33754
rect 28850 33702 28862 33754
rect 28914 33702 28926 33754
rect 28978 33702 28990 33754
rect 29042 33702 29048 33754
rect 1104 33680 29048 33702
rect 16301 33643 16359 33649
rect 16301 33609 16313 33643
rect 16347 33640 16359 33643
rect 16574 33640 16580 33652
rect 16347 33612 16580 33640
rect 16347 33609 16359 33612
rect 16301 33603 16359 33609
rect 16574 33600 16580 33612
rect 16632 33600 16638 33652
rect 21269 33643 21327 33649
rect 21269 33609 21281 33643
rect 21315 33640 21327 33643
rect 21358 33640 21364 33652
rect 21315 33612 21364 33640
rect 21315 33609 21327 33612
rect 21269 33603 21327 33609
rect 21358 33600 21364 33612
rect 21416 33600 21422 33652
rect 25038 33600 25044 33652
rect 25096 33640 25102 33652
rect 26237 33643 26295 33649
rect 26237 33640 26249 33643
rect 25096 33612 26249 33640
rect 25096 33600 25102 33612
rect 26237 33609 26249 33612
rect 26283 33609 26295 33643
rect 26237 33603 26295 33609
rect 26605 33643 26663 33649
rect 26605 33609 26617 33643
rect 26651 33640 26663 33643
rect 26651 33612 27200 33640
rect 26651 33609 26663 33612
rect 26605 33603 26663 33609
rect 16206 33532 16212 33584
rect 16264 33572 16270 33584
rect 18150 33575 18208 33581
rect 18150 33572 18162 33575
rect 16264 33544 18162 33572
rect 16264 33532 16270 33544
rect 18150 33541 18162 33544
rect 18196 33541 18208 33575
rect 18150 33535 18208 33541
rect 24118 33532 24124 33584
rect 24176 33572 24182 33584
rect 27172 33581 27200 33612
rect 27246 33600 27252 33652
rect 27304 33640 27310 33652
rect 27525 33643 27583 33649
rect 27525 33640 27537 33643
rect 27304 33612 27537 33640
rect 27304 33600 27310 33612
rect 27525 33609 27537 33612
rect 27571 33609 27583 33643
rect 28074 33640 28080 33652
rect 28035 33612 28080 33640
rect 27525 33603 27583 33609
rect 28074 33600 28080 33612
rect 28132 33600 28138 33652
rect 27157 33575 27215 33581
rect 24176 33544 26832 33572
rect 24176 33532 24182 33544
rect 15746 33504 15752 33516
rect 15707 33476 15752 33504
rect 15746 33464 15752 33476
rect 15804 33464 15810 33516
rect 15838 33464 15844 33516
rect 15896 33504 15902 33516
rect 16025 33507 16083 33513
rect 16025 33504 16037 33507
rect 15896 33476 16037 33504
rect 15896 33464 15902 33476
rect 16025 33473 16037 33476
rect 16071 33473 16083 33507
rect 16025 33467 16083 33473
rect 16114 33464 16120 33516
rect 16172 33504 16178 33516
rect 16172 33476 17080 33504
rect 16172 33464 16178 33476
rect 17052 33377 17080 33476
rect 20898 33464 20904 33516
rect 20956 33504 20962 33516
rect 21177 33507 21235 33513
rect 21177 33504 21189 33507
rect 20956 33476 21189 33504
rect 20956 33464 20962 33476
rect 21177 33473 21189 33476
rect 21223 33473 21235 33507
rect 21177 33467 21235 33473
rect 21361 33507 21419 33513
rect 21361 33473 21373 33507
rect 21407 33504 21419 33507
rect 21450 33504 21456 33516
rect 21407 33476 21456 33504
rect 21407 33473 21419 33476
rect 21361 33467 21419 33473
rect 21450 33464 21456 33476
rect 21508 33464 21514 33516
rect 23474 33464 23480 33516
rect 23532 33504 23538 33516
rect 23825 33507 23883 33513
rect 23825 33504 23837 33507
rect 23532 33476 23837 33504
rect 23532 33464 23538 33476
rect 23825 33473 23837 33476
rect 23871 33473 23883 33507
rect 26326 33504 26332 33516
rect 23825 33467 23883 33473
rect 26068 33476 26332 33504
rect 18417 33439 18475 33445
rect 18417 33405 18429 33439
rect 18463 33436 18475 33439
rect 18782 33436 18788 33448
rect 18463 33408 18788 33436
rect 18463 33405 18475 33408
rect 18417 33399 18475 33405
rect 18782 33396 18788 33408
rect 18840 33396 18846 33448
rect 21266 33396 21272 33448
rect 21324 33436 21330 33448
rect 22554 33436 22560 33448
rect 21324 33408 22560 33436
rect 21324 33396 21330 33408
rect 22554 33396 22560 33408
rect 22612 33436 22618 33448
rect 23382 33436 23388 33448
rect 22612 33408 23388 33436
rect 22612 33396 22618 33408
rect 23382 33396 23388 33408
rect 23440 33436 23446 33448
rect 26068 33445 26096 33476
rect 26326 33464 26332 33476
rect 26384 33464 26390 33516
rect 26804 33504 26832 33544
rect 27157 33541 27169 33575
rect 27203 33541 27215 33575
rect 27157 33535 27215 33541
rect 27341 33507 27399 33513
rect 27341 33504 27353 33507
rect 26804 33476 27353 33504
rect 27341 33473 27353 33476
rect 27387 33473 27399 33507
rect 27341 33467 27399 33473
rect 27985 33507 28043 33513
rect 27985 33473 27997 33507
rect 28031 33504 28043 33507
rect 28534 33504 28540 33516
rect 28031 33476 28540 33504
rect 28031 33473 28043 33476
rect 27985 33467 28043 33473
rect 28534 33464 28540 33476
rect 28592 33464 28598 33516
rect 23569 33439 23627 33445
rect 23569 33436 23581 33439
rect 23440 33408 23581 33436
rect 23440 33396 23446 33408
rect 23569 33405 23581 33408
rect 23615 33405 23627 33439
rect 23569 33399 23627 33405
rect 26053 33439 26111 33445
rect 26053 33405 26065 33439
rect 26099 33405 26111 33439
rect 26053 33399 26111 33405
rect 26145 33439 26203 33445
rect 26145 33405 26157 33439
rect 26191 33436 26203 33439
rect 28074 33436 28080 33448
rect 26191 33408 28080 33436
rect 26191 33405 26203 33408
rect 26145 33399 26203 33405
rect 28074 33396 28080 33408
rect 28132 33396 28138 33448
rect 17037 33371 17095 33377
rect 17037 33337 17049 33371
rect 17083 33337 17095 33371
rect 17037 33331 17095 33337
rect 3510 33260 3516 33312
rect 3568 33300 3574 33312
rect 13814 33300 13820 33312
rect 3568 33272 13820 33300
rect 3568 33260 3574 33272
rect 13814 33260 13820 33272
rect 13872 33260 13878 33312
rect 15841 33303 15899 33309
rect 15841 33269 15853 33303
rect 15887 33300 15899 33303
rect 16022 33300 16028 33312
rect 15887 33272 16028 33300
rect 15887 33269 15899 33272
rect 15841 33263 15899 33269
rect 16022 33260 16028 33272
rect 16080 33260 16086 33312
rect 23750 33260 23756 33312
rect 23808 33300 23814 33312
rect 24949 33303 25007 33309
rect 24949 33300 24961 33303
rect 23808 33272 24961 33300
rect 23808 33260 23814 33272
rect 24949 33269 24961 33272
rect 24995 33269 25007 33303
rect 24949 33263 25007 33269
rect 1104 33210 28888 33232
rect 1104 33158 4423 33210
rect 4475 33158 4487 33210
rect 4539 33158 4551 33210
rect 4603 33158 4615 33210
rect 4667 33158 4679 33210
rect 4731 33158 11369 33210
rect 11421 33158 11433 33210
rect 11485 33158 11497 33210
rect 11549 33158 11561 33210
rect 11613 33158 11625 33210
rect 11677 33158 18315 33210
rect 18367 33158 18379 33210
rect 18431 33158 18443 33210
rect 18495 33158 18507 33210
rect 18559 33158 18571 33210
rect 18623 33158 25261 33210
rect 25313 33158 25325 33210
rect 25377 33158 25389 33210
rect 25441 33158 25453 33210
rect 25505 33158 25517 33210
rect 25569 33158 28888 33210
rect 1104 33136 28888 33158
rect 16301 33099 16359 33105
rect 16301 33065 16313 33099
rect 16347 33096 16359 33099
rect 16758 33096 16764 33108
rect 16347 33068 16764 33096
rect 16347 33065 16359 33068
rect 16301 33059 16359 33065
rect 16758 33056 16764 33068
rect 16816 33056 16822 33108
rect 23385 33099 23443 33105
rect 23385 33065 23397 33099
rect 23431 33096 23443 33099
rect 23474 33096 23480 33108
rect 23431 33068 23480 33096
rect 23431 33065 23443 33068
rect 23385 33059 23443 33065
rect 23474 33056 23480 33068
rect 23532 33056 23538 33108
rect 24854 33096 24860 33108
rect 24815 33068 24860 33096
rect 24854 33056 24860 33068
rect 24912 33056 24918 33108
rect 15746 32988 15752 33040
rect 15804 33028 15810 33040
rect 16482 33028 16488 33040
rect 15804 33000 16488 33028
rect 15804 32988 15810 33000
rect 16482 32988 16488 33000
rect 16540 33028 16546 33040
rect 17037 33031 17095 33037
rect 17037 33028 17049 33031
rect 16540 33000 17049 33028
rect 16540 32988 16546 33000
rect 17037 32997 17049 33000
rect 17083 32997 17095 33031
rect 17037 32991 17095 32997
rect 20257 32963 20315 32969
rect 20257 32929 20269 32963
rect 20303 32960 20315 32963
rect 20806 32960 20812 32972
rect 20303 32932 20812 32960
rect 20303 32929 20315 32932
rect 20257 32923 20315 32929
rect 20806 32920 20812 32932
rect 20864 32920 20870 32972
rect 23474 32920 23480 32972
rect 23532 32960 23538 32972
rect 23750 32960 23756 32972
rect 23532 32932 23756 32960
rect 23532 32920 23538 32932
rect 23750 32920 23756 32932
rect 23808 32960 23814 32972
rect 27522 32960 27528 32972
rect 23808 32932 24072 32960
rect 27483 32932 27528 32960
rect 23808 32920 23814 32932
rect 16022 32892 16028 32904
rect 15983 32864 16028 32892
rect 16022 32852 16028 32864
rect 16080 32852 16086 32904
rect 16758 32852 16764 32904
rect 16816 32892 16822 32904
rect 17129 32895 17187 32901
rect 17129 32892 17141 32895
rect 16816 32864 17141 32892
rect 16816 32852 16822 32864
rect 17129 32861 17141 32864
rect 17175 32861 17187 32895
rect 17129 32855 17187 32861
rect 20073 32895 20131 32901
rect 20073 32861 20085 32895
rect 20119 32861 20131 32895
rect 20073 32855 20131 32861
rect 17034 32784 17040 32836
rect 17092 32824 17098 32836
rect 19978 32824 19984 32836
rect 17092 32796 19984 32824
rect 17092 32784 17098 32796
rect 19978 32784 19984 32796
rect 20036 32824 20042 32836
rect 20088 32824 20116 32855
rect 20162 32852 20168 32904
rect 20220 32892 20226 32904
rect 20220 32864 20265 32892
rect 20220 32852 20226 32864
rect 20346 32852 20352 32904
rect 20404 32892 20410 32904
rect 20533 32895 20591 32901
rect 20404 32864 20449 32892
rect 20404 32852 20410 32864
rect 20533 32861 20545 32895
rect 20579 32861 20591 32895
rect 23566 32892 23572 32904
rect 23527 32864 23572 32892
rect 20533 32855 20591 32861
rect 20036 32796 20116 32824
rect 20036 32784 20042 32796
rect 20254 32784 20260 32836
rect 20312 32824 20318 32836
rect 20548 32824 20576 32855
rect 23566 32852 23572 32864
rect 23624 32852 23630 32904
rect 23658 32852 23664 32904
rect 23716 32892 23722 32904
rect 24044 32901 24072 32932
rect 27522 32920 27528 32932
rect 27580 32920 27586 32972
rect 23845 32895 23903 32901
rect 23845 32892 23857 32895
rect 23716 32864 23857 32892
rect 23716 32852 23722 32864
rect 23845 32861 23857 32864
rect 23891 32861 23903 32895
rect 23845 32855 23903 32861
rect 24029 32895 24087 32901
rect 24029 32861 24041 32895
rect 24075 32861 24087 32895
rect 25866 32892 25872 32904
rect 25827 32864 25872 32892
rect 24029 32855 24087 32861
rect 20312 32796 20576 32824
rect 20312 32784 20318 32796
rect 16390 32716 16396 32768
rect 16448 32756 16454 32768
rect 16485 32759 16543 32765
rect 16485 32756 16497 32759
rect 16448 32728 16497 32756
rect 16448 32716 16454 32728
rect 16485 32725 16497 32728
rect 16531 32725 16543 32759
rect 16485 32719 16543 32725
rect 18874 32716 18880 32768
rect 18932 32756 18938 32768
rect 19889 32759 19947 32765
rect 19889 32756 19901 32759
rect 18932 32728 19901 32756
rect 18932 32716 18938 32728
rect 19889 32725 19901 32728
rect 19935 32725 19947 32759
rect 23860 32756 23888 32855
rect 25866 32852 25872 32864
rect 25924 32852 25930 32904
rect 28350 32852 28356 32904
rect 28408 32892 28414 32904
rect 28408 32864 28453 32892
rect 28408 32852 28414 32864
rect 25038 32824 25044 32836
rect 24999 32796 25044 32824
rect 25038 32784 25044 32796
rect 25096 32784 25102 32836
rect 28166 32824 28172 32836
rect 28127 32796 28172 32824
rect 28166 32784 28172 32796
rect 28224 32784 28230 32836
rect 24210 32756 24216 32768
rect 23860 32728 24216 32756
rect 19889 32719 19947 32725
rect 24210 32716 24216 32728
rect 24268 32756 24274 32768
rect 24673 32759 24731 32765
rect 24673 32756 24685 32759
rect 24268 32728 24685 32756
rect 24268 32716 24274 32728
rect 24673 32725 24685 32728
rect 24719 32725 24731 32759
rect 24673 32719 24731 32725
rect 24841 32759 24899 32765
rect 24841 32725 24853 32759
rect 24887 32756 24899 32759
rect 25685 32759 25743 32765
rect 25685 32756 25697 32759
rect 24887 32728 25697 32756
rect 24887 32725 24899 32728
rect 24841 32719 24899 32725
rect 25685 32725 25697 32728
rect 25731 32725 25743 32759
rect 25685 32719 25743 32725
rect 1104 32666 29048 32688
rect 1104 32614 7896 32666
rect 7948 32614 7960 32666
rect 8012 32614 8024 32666
rect 8076 32614 8088 32666
rect 8140 32614 8152 32666
rect 8204 32614 14842 32666
rect 14894 32614 14906 32666
rect 14958 32614 14970 32666
rect 15022 32614 15034 32666
rect 15086 32614 15098 32666
rect 15150 32614 21788 32666
rect 21840 32614 21852 32666
rect 21904 32614 21916 32666
rect 21968 32614 21980 32666
rect 22032 32614 22044 32666
rect 22096 32614 28734 32666
rect 28786 32614 28798 32666
rect 28850 32614 28862 32666
rect 28914 32614 28926 32666
rect 28978 32614 28990 32666
rect 29042 32614 29048 32666
rect 1104 32592 29048 32614
rect 18708 32524 19748 32552
rect 17586 32376 17592 32428
rect 17644 32416 17650 32428
rect 18708 32425 18736 32524
rect 18785 32487 18843 32493
rect 18785 32453 18797 32487
rect 18831 32484 18843 32487
rect 19582 32487 19640 32493
rect 19582 32484 19594 32487
rect 18831 32456 19594 32484
rect 18831 32453 18843 32456
rect 18785 32447 18843 32453
rect 19582 32453 19594 32456
rect 19628 32453 19640 32487
rect 19720 32484 19748 32524
rect 20162 32512 20168 32564
rect 20220 32552 20226 32564
rect 21269 32555 21327 32561
rect 21269 32552 21281 32555
rect 20220 32524 21281 32552
rect 20220 32512 20226 32524
rect 21269 32521 21281 32524
rect 21315 32521 21327 32555
rect 21269 32515 21327 32521
rect 21450 32484 21456 32496
rect 19720 32456 21456 32484
rect 19582 32447 19640 32453
rect 21450 32444 21456 32456
rect 21508 32444 21514 32496
rect 18693 32419 18751 32425
rect 18693 32416 18705 32419
rect 17644 32388 18705 32416
rect 17644 32376 17650 32388
rect 18693 32385 18705 32388
rect 18739 32385 18751 32419
rect 18874 32416 18880 32428
rect 18835 32388 18880 32416
rect 18693 32379 18751 32385
rect 18874 32376 18880 32388
rect 18932 32376 18938 32428
rect 21174 32416 21180 32428
rect 21135 32388 21180 32416
rect 21174 32376 21180 32388
rect 21232 32376 21238 32428
rect 21361 32419 21419 32425
rect 21361 32385 21373 32419
rect 21407 32385 21419 32419
rect 23106 32416 23112 32428
rect 23067 32388 23112 32416
rect 21361 32379 21419 32385
rect 12713 32351 12771 32357
rect 12713 32317 12725 32351
rect 12759 32317 12771 32351
rect 12894 32348 12900 32360
rect 12855 32320 12900 32348
rect 12713 32311 12771 32317
rect 12728 32280 12756 32311
rect 12894 32308 12900 32320
rect 12952 32308 12958 32360
rect 13814 32348 13820 32360
rect 13775 32320 13820 32348
rect 13814 32308 13820 32320
rect 13872 32308 13878 32360
rect 19337 32351 19395 32357
rect 19337 32348 19349 32351
rect 18892 32320 19349 32348
rect 18892 32292 18920 32320
rect 19337 32317 19349 32320
rect 19383 32317 19395 32351
rect 21376 32348 21404 32379
rect 23106 32376 23112 32388
rect 23164 32376 23170 32428
rect 25866 32416 25872 32428
rect 25827 32388 25872 32416
rect 25866 32376 25872 32388
rect 25924 32376 25930 32428
rect 27433 32419 27491 32425
rect 27433 32385 27445 32419
rect 27479 32416 27491 32419
rect 28350 32416 28356 32428
rect 27479 32388 28356 32416
rect 27479 32385 27491 32388
rect 27433 32379 27491 32385
rect 28350 32376 28356 32388
rect 28408 32376 28414 32428
rect 19337 32311 19395 32317
rect 20732 32320 21404 32348
rect 20732 32292 20760 32320
rect 13262 32280 13268 32292
rect 12728 32252 13268 32280
rect 13262 32240 13268 32252
rect 13320 32240 13326 32292
rect 18874 32240 18880 32292
rect 18932 32240 18938 32292
rect 20714 32280 20720 32292
rect 20675 32252 20720 32280
rect 20714 32240 20720 32252
rect 20772 32240 20778 32292
rect 23293 32215 23351 32221
rect 23293 32181 23305 32215
rect 23339 32212 23351 32215
rect 23658 32212 23664 32224
rect 23339 32184 23664 32212
rect 23339 32181 23351 32184
rect 23293 32175 23351 32181
rect 23658 32172 23664 32184
rect 23716 32172 23722 32224
rect 25958 32212 25964 32224
rect 25919 32184 25964 32212
rect 25958 32172 25964 32184
rect 26016 32172 26022 32224
rect 26602 32172 26608 32224
rect 26660 32212 26666 32224
rect 27893 32215 27951 32221
rect 27893 32212 27905 32215
rect 26660 32184 27905 32212
rect 26660 32172 26666 32184
rect 27893 32181 27905 32184
rect 27939 32181 27951 32215
rect 27893 32175 27951 32181
rect 1104 32122 28888 32144
rect 1104 32070 4423 32122
rect 4475 32070 4487 32122
rect 4539 32070 4551 32122
rect 4603 32070 4615 32122
rect 4667 32070 4679 32122
rect 4731 32070 11369 32122
rect 11421 32070 11433 32122
rect 11485 32070 11497 32122
rect 11549 32070 11561 32122
rect 11613 32070 11625 32122
rect 11677 32070 18315 32122
rect 18367 32070 18379 32122
rect 18431 32070 18443 32122
rect 18495 32070 18507 32122
rect 18559 32070 18571 32122
rect 18623 32070 25261 32122
rect 25313 32070 25325 32122
rect 25377 32070 25389 32122
rect 25441 32070 25453 32122
rect 25505 32070 25517 32122
rect 25569 32070 28888 32122
rect 1104 32048 28888 32070
rect 12894 32008 12900 32020
rect 12855 31980 12900 32008
rect 12894 31968 12900 31980
rect 12952 31968 12958 32020
rect 16574 31968 16580 32020
rect 16632 32008 16638 32020
rect 19426 32008 19432 32020
rect 16632 31980 16712 32008
rect 19387 31980 19432 32008
rect 16632 31968 16638 31980
rect 12802 31940 12808 31952
rect 12715 31912 12808 31940
rect 12802 31900 12808 31912
rect 12860 31940 12866 31952
rect 16684 31949 16712 31980
rect 19426 31968 19432 31980
rect 19484 31968 19490 32020
rect 20717 32011 20775 32017
rect 19536 31980 20484 32008
rect 16669 31943 16727 31949
rect 12860 31912 16620 31940
rect 12860 31900 12866 31912
rect 12820 31813 12848 31900
rect 16482 31872 16488 31884
rect 16443 31844 16488 31872
rect 16482 31832 16488 31844
rect 16540 31832 16546 31884
rect 16592 31872 16620 31912
rect 16669 31909 16681 31943
rect 16715 31909 16727 31943
rect 19536 31940 19564 31980
rect 20346 31940 20352 31952
rect 16669 31903 16727 31909
rect 16776 31912 19564 31940
rect 19812 31912 20352 31940
rect 16776 31872 16804 31912
rect 16592 31844 16804 31872
rect 16945 31875 17003 31881
rect 16945 31841 16957 31875
rect 16991 31872 17003 31875
rect 17497 31875 17555 31881
rect 16991 31844 17448 31872
rect 16991 31841 17003 31844
rect 16945 31835 17003 31841
rect 12805 31807 12863 31813
rect 12805 31773 12817 31807
rect 12851 31773 12863 31807
rect 12805 31767 12863 31773
rect 16301 31807 16359 31813
rect 16301 31773 16313 31807
rect 16347 31804 16359 31807
rect 16574 31804 16580 31816
rect 16347 31776 16436 31804
rect 16535 31776 16580 31804
rect 16347 31773 16359 31776
rect 16301 31767 16359 31773
rect 16408 31736 16436 31776
rect 16574 31764 16580 31776
rect 16632 31764 16638 31816
rect 16761 31807 16819 31813
rect 16761 31773 16773 31807
rect 16807 31804 16819 31807
rect 17034 31804 17040 31816
rect 16807 31776 17040 31804
rect 16807 31773 16819 31776
rect 16761 31767 16819 31773
rect 17034 31764 17040 31776
rect 17092 31764 17098 31816
rect 17420 31813 17448 31844
rect 17497 31841 17509 31875
rect 17543 31872 17555 31875
rect 18598 31872 18604 31884
rect 17543 31844 18604 31872
rect 17543 31841 17555 31844
rect 17497 31835 17555 31841
rect 18598 31832 18604 31844
rect 18656 31832 18662 31884
rect 19812 31872 19840 31912
rect 20346 31900 20352 31912
rect 20404 31900 20410 31952
rect 20456 31940 20484 31980
rect 20717 31977 20729 32011
rect 20763 32008 20775 32011
rect 20806 32008 20812 32020
rect 20763 31980 20812 32008
rect 20763 31977 20775 31980
rect 20717 31971 20775 31977
rect 20806 31968 20812 31980
rect 20864 31968 20870 32020
rect 22557 32011 22615 32017
rect 20916 31980 22508 32008
rect 20916 31940 20944 31980
rect 20456 31912 20944 31940
rect 22480 31940 22508 31980
rect 22557 31977 22569 32011
rect 22603 32008 22615 32011
rect 22922 32008 22928 32020
rect 22603 31980 22928 32008
rect 22603 31977 22615 31980
rect 22557 31971 22615 31977
rect 22922 31968 22928 31980
rect 22980 32008 22986 32020
rect 23106 32008 23112 32020
rect 22980 31980 23112 32008
rect 22980 31968 22986 31980
rect 23106 31968 23112 31980
rect 23164 31968 23170 32020
rect 25866 32008 25872 32020
rect 23308 31980 25872 32008
rect 23308 31940 23336 31980
rect 25866 31968 25872 31980
rect 25924 32008 25930 32020
rect 27062 32008 27068 32020
rect 25924 31980 27068 32008
rect 25924 31968 25930 31980
rect 27062 31968 27068 31980
rect 27120 31968 27126 32020
rect 28166 32008 28172 32020
rect 28127 31980 28172 32008
rect 28166 31968 28172 31980
rect 28224 31968 28230 32020
rect 24302 31940 24308 31952
rect 22480 31912 23336 31940
rect 23400 31912 24308 31940
rect 19720 31844 19840 31872
rect 20088 31844 20760 31872
rect 17405 31807 17463 31813
rect 17405 31773 17417 31807
rect 17451 31773 17463 31807
rect 17586 31804 17592 31816
rect 17547 31776 17592 31804
rect 17405 31767 17463 31773
rect 17586 31764 17592 31776
rect 17644 31764 17650 31816
rect 19720 31813 19748 31844
rect 20088 31816 20116 31844
rect 19705 31807 19763 31813
rect 19705 31773 19717 31807
rect 19751 31773 19763 31807
rect 19705 31767 19763 31773
rect 19797 31807 19855 31813
rect 19797 31773 19809 31807
rect 19843 31773 19855 31807
rect 19797 31767 19855 31773
rect 16850 31736 16856 31748
rect 16408 31708 16856 31736
rect 16850 31696 16856 31708
rect 16908 31696 16914 31748
rect 19610 31696 19616 31748
rect 19668 31736 19674 31748
rect 19812 31736 19840 31767
rect 19886 31764 19892 31816
rect 19944 31804 19950 31816
rect 19944 31776 19989 31804
rect 19944 31764 19950 31776
rect 20070 31764 20076 31816
rect 20128 31804 20134 31816
rect 20128 31776 20173 31804
rect 20128 31764 20134 31776
rect 20346 31764 20352 31816
rect 20404 31804 20410 31816
rect 20732 31813 20760 31844
rect 20533 31807 20591 31813
rect 20533 31804 20545 31807
rect 20404 31776 20545 31804
rect 20404 31764 20410 31776
rect 20533 31773 20545 31776
rect 20579 31773 20591 31807
rect 20533 31767 20591 31773
rect 20717 31807 20775 31813
rect 20717 31773 20729 31807
rect 20763 31773 20775 31807
rect 20717 31767 20775 31773
rect 21177 31807 21235 31813
rect 21177 31773 21189 31807
rect 21223 31804 21235 31807
rect 21266 31804 21272 31816
rect 21223 31776 21272 31804
rect 21223 31773 21235 31776
rect 21177 31767 21235 31773
rect 21266 31764 21272 31776
rect 21324 31764 21330 31816
rect 21444 31807 21502 31813
rect 21444 31773 21456 31807
rect 21490 31804 21502 31807
rect 22186 31804 22192 31816
rect 21490 31776 22192 31804
rect 21490 31773 21502 31776
rect 21444 31767 21502 31773
rect 22186 31764 22192 31776
rect 22244 31764 22250 31816
rect 23198 31807 23256 31813
rect 23198 31773 23210 31807
rect 23244 31804 23256 31807
rect 23400 31804 23428 31912
rect 24302 31900 24308 31912
rect 24360 31900 24366 31952
rect 23658 31872 23664 31884
rect 23619 31844 23664 31872
rect 23658 31832 23664 31844
rect 23716 31832 23722 31884
rect 25774 31872 25780 31884
rect 25735 31844 25780 31872
rect 25774 31832 25780 31844
rect 25832 31832 25838 31884
rect 25958 31872 25964 31884
rect 25919 31844 25964 31872
rect 25958 31832 25964 31844
rect 26016 31832 26022 31884
rect 27522 31872 27528 31884
rect 27483 31844 27528 31872
rect 27522 31832 27528 31844
rect 27580 31832 27586 31884
rect 23566 31804 23572 31816
rect 23244 31776 23428 31804
rect 23527 31776 23572 31804
rect 23244 31773 23256 31776
rect 23198 31767 23256 31773
rect 23566 31764 23572 31776
rect 23624 31764 23630 31816
rect 27890 31764 27896 31816
rect 27948 31804 27954 31816
rect 28077 31807 28135 31813
rect 28077 31804 28089 31807
rect 27948 31776 28089 31804
rect 27948 31764 27954 31776
rect 28077 31773 28089 31776
rect 28123 31804 28135 31807
rect 28166 31804 28172 31816
rect 28123 31776 28172 31804
rect 28123 31773 28135 31776
rect 28077 31767 28135 31773
rect 28166 31764 28172 31776
rect 28224 31764 28230 31816
rect 19668 31708 19840 31736
rect 19668 31696 19674 31708
rect 23934 31696 23940 31748
rect 23992 31736 23998 31748
rect 24765 31739 24823 31745
rect 24765 31736 24777 31739
rect 23992 31708 24777 31736
rect 23992 31696 23998 31708
rect 24765 31705 24777 31708
rect 24811 31705 24823 31739
rect 24946 31736 24952 31748
rect 24907 31708 24952 31736
rect 24765 31699 24823 31705
rect 24946 31696 24952 31708
rect 25004 31696 25010 31748
rect 22554 31628 22560 31680
rect 22612 31668 22618 31680
rect 23017 31671 23075 31677
rect 23017 31668 23029 31671
rect 22612 31640 23029 31668
rect 22612 31628 22618 31640
rect 23017 31637 23029 31640
rect 23063 31637 23075 31671
rect 23198 31668 23204 31680
rect 23159 31640 23204 31668
rect 23017 31631 23075 31637
rect 23198 31628 23204 31640
rect 23256 31628 23262 31680
rect 1104 31578 29048 31600
rect 1104 31526 7896 31578
rect 7948 31526 7960 31578
rect 8012 31526 8024 31578
rect 8076 31526 8088 31578
rect 8140 31526 8152 31578
rect 8204 31526 14842 31578
rect 14894 31526 14906 31578
rect 14958 31526 14970 31578
rect 15022 31526 15034 31578
rect 15086 31526 15098 31578
rect 15150 31526 21788 31578
rect 21840 31526 21852 31578
rect 21904 31526 21916 31578
rect 21968 31526 21980 31578
rect 22032 31526 22044 31578
rect 22096 31526 28734 31578
rect 28786 31526 28798 31578
rect 28850 31526 28862 31578
rect 28914 31526 28926 31578
rect 28978 31526 28990 31578
rect 29042 31526 29048 31578
rect 1104 31504 29048 31526
rect 16101 31467 16159 31473
rect 16101 31433 16113 31467
rect 16147 31464 16159 31467
rect 16206 31464 16212 31476
rect 16147 31436 16212 31464
rect 16147 31433 16159 31436
rect 16101 31427 16159 31433
rect 16206 31424 16212 31436
rect 16264 31424 16270 31476
rect 16666 31424 16672 31476
rect 16724 31464 16730 31476
rect 16945 31467 17003 31473
rect 16945 31464 16957 31467
rect 16724 31436 16957 31464
rect 16724 31424 16730 31436
rect 16945 31433 16957 31436
rect 16991 31433 17003 31467
rect 16945 31427 17003 31433
rect 22097 31467 22155 31473
rect 22097 31433 22109 31467
rect 22143 31464 22155 31467
rect 22186 31464 22192 31476
rect 22143 31436 22192 31464
rect 22143 31433 22155 31436
rect 22097 31427 22155 31433
rect 22186 31424 22192 31436
rect 22244 31424 22250 31476
rect 23198 31464 23204 31476
rect 23159 31436 23204 31464
rect 23198 31424 23204 31436
rect 23256 31424 23262 31476
rect 23566 31424 23572 31476
rect 23624 31464 23630 31476
rect 23845 31467 23903 31473
rect 23845 31464 23857 31467
rect 23624 31436 23857 31464
rect 23624 31424 23630 31436
rect 23845 31433 23857 31436
rect 23891 31433 23903 31467
rect 23845 31427 23903 31433
rect 16301 31399 16359 31405
rect 16301 31365 16313 31399
rect 16347 31365 16359 31399
rect 16301 31359 16359 31365
rect 16316 31328 16344 31359
rect 18598 31356 18604 31408
rect 18656 31405 18662 31408
rect 18656 31396 18668 31405
rect 18656 31368 18701 31396
rect 18656 31359 18668 31368
rect 18656 31356 18662 31359
rect 22462 31356 22468 31408
rect 22520 31396 22526 31408
rect 22922 31396 22928 31408
rect 22520 31368 22928 31396
rect 22520 31356 22526 31368
rect 22922 31356 22928 31368
rect 22980 31356 22986 31408
rect 24210 31396 24216 31408
rect 24171 31368 24216 31396
rect 24210 31356 24216 31368
rect 24268 31356 24274 31408
rect 16758 31328 16764 31340
rect 16316 31300 16764 31328
rect 16758 31288 16764 31300
rect 16816 31328 16822 31340
rect 16853 31331 16911 31337
rect 16853 31328 16865 31331
rect 16816 31300 16865 31328
rect 16816 31288 16822 31300
rect 16853 31297 16865 31300
rect 16899 31297 16911 31331
rect 16853 31291 16911 31297
rect 17037 31331 17095 31337
rect 17037 31297 17049 31331
rect 17083 31328 17095 31331
rect 17218 31328 17224 31340
rect 17083 31300 17224 31328
rect 17083 31297 17095 31300
rect 17037 31291 17095 31297
rect 16868 31260 16896 31291
rect 17218 31288 17224 31300
rect 17276 31288 17282 31340
rect 20165 31331 20223 31337
rect 20165 31297 20177 31331
rect 20211 31328 20223 31331
rect 21082 31328 21088 31340
rect 20211 31300 21088 31328
rect 20211 31297 20223 31300
rect 20165 31291 20223 31297
rect 21082 31288 21088 31300
rect 21140 31288 21146 31340
rect 21634 31288 21640 31340
rect 21692 31328 21698 31340
rect 22005 31331 22063 31337
rect 22005 31328 22017 31331
rect 21692 31300 22017 31328
rect 21692 31288 21698 31300
rect 22005 31297 22017 31300
rect 22051 31297 22063 31331
rect 22005 31291 22063 31297
rect 22189 31331 22247 31337
rect 22189 31297 22201 31331
rect 22235 31328 22247 31331
rect 22554 31328 22560 31340
rect 22235 31300 22560 31328
rect 22235 31297 22247 31300
rect 22189 31291 22247 31297
rect 22554 31288 22560 31300
rect 22612 31288 22618 31340
rect 22649 31331 22707 31337
rect 22649 31297 22661 31331
rect 22695 31297 22707 31331
rect 22830 31328 22836 31340
rect 22791 31300 22836 31328
rect 22649 31291 22707 31297
rect 18874 31260 18880 31272
rect 16868 31232 17540 31260
rect 18835 31232 18880 31260
rect 15933 31195 15991 31201
rect 15933 31161 15945 31195
rect 15979 31192 15991 31195
rect 16574 31192 16580 31204
rect 15979 31164 16580 31192
rect 15979 31161 15991 31164
rect 15933 31155 15991 31161
rect 16574 31152 16580 31164
rect 16632 31152 16638 31204
rect 17512 31201 17540 31232
rect 18874 31220 18880 31232
rect 18932 31220 18938 31272
rect 22664 31260 22692 31291
rect 22830 31288 22836 31300
rect 22888 31288 22894 31340
rect 23017 31331 23075 31337
rect 23017 31297 23029 31331
rect 23063 31328 23075 31331
rect 23106 31328 23112 31340
rect 23063 31300 23112 31328
rect 23063 31297 23075 31300
rect 23017 31291 23075 31297
rect 23106 31288 23112 31300
rect 23164 31288 23170 31340
rect 23934 31288 23940 31340
rect 23992 31328 23998 31340
rect 24029 31331 24087 31337
rect 24029 31328 24041 31331
rect 23992 31300 24041 31328
rect 23992 31288 23998 31300
rect 24029 31297 24041 31300
rect 24075 31297 24087 31331
rect 24029 31291 24087 31297
rect 26602 31288 26608 31340
rect 26660 31328 26666 31340
rect 26660 31300 26705 31328
rect 26660 31288 26666 31300
rect 27614 31288 27620 31340
rect 27672 31328 27678 31340
rect 27709 31331 27767 31337
rect 27709 31328 27721 31331
rect 27672 31300 27721 31328
rect 27672 31288 27678 31300
rect 27709 31297 27721 31300
rect 27755 31297 27767 31331
rect 27709 31291 27767 31297
rect 23382 31260 23388 31272
rect 22664 31232 23388 31260
rect 23382 31220 23388 31232
rect 23440 31220 23446 31272
rect 26142 31260 26148 31272
rect 26103 31232 26148 31260
rect 26142 31220 26148 31232
rect 26200 31220 26206 31272
rect 26421 31263 26479 31269
rect 26421 31229 26433 31263
rect 26467 31260 26479 31263
rect 27801 31263 27859 31269
rect 27801 31260 27813 31263
rect 26467 31232 27813 31260
rect 26467 31229 26479 31232
rect 26421 31223 26479 31229
rect 27801 31229 27813 31232
rect 27847 31229 27859 31263
rect 27801 31223 27859 31229
rect 17497 31195 17555 31201
rect 17497 31161 17509 31195
rect 17543 31161 17555 31195
rect 17497 31155 17555 31161
rect 16117 31127 16175 31133
rect 16117 31093 16129 31127
rect 16163 31124 16175 31127
rect 16666 31124 16672 31136
rect 16163 31096 16672 31124
rect 16163 31093 16175 31096
rect 16117 31087 16175 31093
rect 16666 31084 16672 31096
rect 16724 31084 16730 31136
rect 19886 31084 19892 31136
rect 19944 31124 19950 31136
rect 20070 31124 20076 31136
rect 19944 31096 20076 31124
rect 19944 31084 19950 31096
rect 20070 31084 20076 31096
rect 20128 31124 20134 31136
rect 20257 31127 20315 31133
rect 20257 31124 20269 31127
rect 20128 31096 20269 31124
rect 20128 31084 20134 31096
rect 20257 31093 20269 31096
rect 20303 31093 20315 31127
rect 20257 31087 20315 31093
rect 1104 31034 28888 31056
rect 1104 30982 4423 31034
rect 4475 30982 4487 31034
rect 4539 30982 4551 31034
rect 4603 30982 4615 31034
rect 4667 30982 4679 31034
rect 4731 30982 11369 31034
rect 11421 30982 11433 31034
rect 11485 30982 11497 31034
rect 11549 30982 11561 31034
rect 11613 30982 11625 31034
rect 11677 30982 18315 31034
rect 18367 30982 18379 31034
rect 18431 30982 18443 31034
rect 18495 30982 18507 31034
rect 18559 30982 18571 31034
rect 18623 30982 25261 31034
rect 25313 30982 25325 31034
rect 25377 30982 25389 31034
rect 25441 30982 25453 31034
rect 25505 30982 25517 31034
rect 25569 30982 28888 31034
rect 1104 30960 28888 30982
rect 15838 30880 15844 30932
rect 15896 30920 15902 30932
rect 16025 30923 16083 30929
rect 16025 30920 16037 30923
rect 15896 30892 16037 30920
rect 15896 30880 15902 30892
rect 16025 30889 16037 30892
rect 16071 30889 16083 30923
rect 16025 30883 16083 30889
rect 22649 30923 22707 30929
rect 22649 30889 22661 30923
rect 22695 30920 22707 30923
rect 22830 30920 22836 30932
rect 22695 30892 22836 30920
rect 22695 30889 22707 30892
rect 22649 30883 22707 30889
rect 22830 30880 22836 30892
rect 22888 30880 22894 30932
rect 23106 30920 23112 30932
rect 23067 30892 23112 30920
rect 23106 30880 23112 30892
rect 23164 30880 23170 30932
rect 24946 30880 24952 30932
rect 25004 30920 25010 30932
rect 25777 30923 25835 30929
rect 25777 30920 25789 30923
rect 25004 30892 25789 30920
rect 25004 30880 25010 30892
rect 25777 30889 25789 30892
rect 25823 30889 25835 30923
rect 25777 30883 25835 30889
rect 16298 30744 16304 30796
rect 16356 30784 16362 30796
rect 23293 30787 23351 30793
rect 23293 30784 23305 30787
rect 16356 30756 16804 30784
rect 16356 30744 16362 30756
rect 16117 30719 16175 30725
rect 16117 30685 16129 30719
rect 16163 30716 16175 30719
rect 16666 30716 16672 30728
rect 16163 30688 16672 30716
rect 16163 30685 16175 30688
rect 16117 30679 16175 30685
rect 16666 30676 16672 30688
rect 16724 30676 16730 30728
rect 16776 30725 16804 30756
rect 22664 30756 23305 30784
rect 16761 30719 16819 30725
rect 16761 30685 16773 30719
rect 16807 30685 16819 30719
rect 16761 30679 16819 30685
rect 18325 30719 18383 30725
rect 18325 30685 18337 30719
rect 18371 30716 18383 30719
rect 19334 30716 19340 30728
rect 18371 30688 19340 30716
rect 18371 30685 18383 30688
rect 18325 30679 18383 30685
rect 19334 30676 19340 30688
rect 19392 30676 19398 30728
rect 22462 30716 22468 30728
rect 22423 30688 22468 30716
rect 22462 30676 22468 30688
rect 22520 30676 22526 30728
rect 22664 30725 22692 30756
rect 23293 30753 23305 30756
rect 23339 30784 23351 30787
rect 23934 30784 23940 30796
rect 23339 30756 23940 30784
rect 23339 30753 23351 30756
rect 23293 30747 23351 30753
rect 23934 30744 23940 30756
rect 23992 30744 23998 30796
rect 28258 30784 28264 30796
rect 28219 30756 28264 30784
rect 28258 30744 28264 30756
rect 28316 30744 28322 30796
rect 22649 30719 22707 30725
rect 22649 30685 22661 30719
rect 22695 30685 22707 30719
rect 22649 30679 22707 30685
rect 23382 30676 23388 30728
rect 23440 30716 23446 30728
rect 23440 30688 23485 30716
rect 23440 30676 23446 30688
rect 23566 30676 23572 30728
rect 23624 30716 23630 30728
rect 24765 30719 24823 30725
rect 24765 30716 24777 30719
rect 23624 30688 24777 30716
rect 23624 30676 23630 30688
rect 24765 30685 24777 30688
rect 24811 30685 24823 30719
rect 24765 30679 24823 30685
rect 24854 30676 24860 30728
rect 24912 30716 24918 30728
rect 24912 30688 24957 30716
rect 24912 30676 24918 30688
rect 26326 30676 26332 30728
rect 26384 30716 26390 30728
rect 26421 30719 26479 30725
rect 26421 30716 26433 30719
rect 26384 30688 26433 30716
rect 26384 30676 26390 30688
rect 26421 30685 26433 30688
rect 26467 30685 26479 30719
rect 26421 30679 26479 30685
rect 18693 30651 18751 30657
rect 18693 30617 18705 30651
rect 18739 30648 18751 30651
rect 21634 30648 21640 30660
rect 18739 30620 21640 30648
rect 18739 30617 18751 30620
rect 18693 30611 18751 30617
rect 21634 30608 21640 30620
rect 21692 30608 21698 30660
rect 23658 30648 23664 30660
rect 23619 30620 23664 30648
rect 23658 30608 23664 30620
rect 23716 30608 23722 30660
rect 23750 30608 23756 30660
rect 23808 30648 23814 30660
rect 25130 30648 25136 30660
rect 23808 30620 23853 30648
rect 23952 30620 25136 30648
rect 23808 30608 23814 30620
rect 16945 30583 17003 30589
rect 16945 30549 16957 30583
rect 16991 30580 17003 30583
rect 17218 30580 17224 30592
rect 16991 30552 17224 30580
rect 16991 30549 17003 30552
rect 16945 30543 17003 30549
rect 17218 30540 17224 30552
rect 17276 30540 17282 30592
rect 23106 30540 23112 30592
rect 23164 30580 23170 30592
rect 23952 30580 23980 30620
rect 25130 30608 25136 30620
rect 25188 30648 25194 30660
rect 25409 30651 25467 30657
rect 25409 30648 25421 30651
rect 25188 30620 25421 30648
rect 25188 30608 25194 30620
rect 25409 30617 25421 30620
rect 25455 30617 25467 30651
rect 25409 30611 25467 30617
rect 25593 30651 25651 30657
rect 25593 30617 25605 30651
rect 25639 30617 25651 30651
rect 26602 30648 26608 30660
rect 26563 30620 26608 30648
rect 25593 30611 25651 30617
rect 24578 30580 24584 30592
rect 23164 30552 23980 30580
rect 24539 30552 24584 30580
rect 23164 30540 23170 30552
rect 24578 30540 24584 30552
rect 24636 30540 24642 30592
rect 24762 30540 24768 30592
rect 24820 30580 24826 30592
rect 25608 30580 25636 30611
rect 26602 30608 26608 30620
rect 26660 30608 26666 30660
rect 24820 30552 25636 30580
rect 24820 30540 24826 30552
rect 1104 30490 29048 30512
rect 1104 30438 7896 30490
rect 7948 30438 7960 30490
rect 8012 30438 8024 30490
rect 8076 30438 8088 30490
rect 8140 30438 8152 30490
rect 8204 30438 14842 30490
rect 14894 30438 14906 30490
rect 14958 30438 14970 30490
rect 15022 30438 15034 30490
rect 15086 30438 15098 30490
rect 15150 30438 21788 30490
rect 21840 30438 21852 30490
rect 21904 30438 21916 30490
rect 21968 30438 21980 30490
rect 22032 30438 22044 30490
rect 22096 30438 28734 30490
rect 28786 30438 28798 30490
rect 28850 30438 28862 30490
rect 28914 30438 28926 30490
rect 28978 30438 28990 30490
rect 29042 30438 29048 30490
rect 1104 30416 29048 30438
rect 19334 30336 19340 30388
rect 19392 30376 19398 30388
rect 20165 30379 20223 30385
rect 19392 30348 20024 30376
rect 19392 30336 19398 30348
rect 16666 30308 16672 30320
rect 16132 30280 16672 30308
rect 16132 30249 16160 30280
rect 16666 30268 16672 30280
rect 16724 30268 16730 30320
rect 16850 30268 16856 30320
rect 16908 30308 16914 30320
rect 19153 30311 19211 30317
rect 16908 30280 17540 30308
rect 16908 30268 16914 30280
rect 17512 30252 17540 30280
rect 19153 30277 19165 30311
rect 19199 30308 19211 30311
rect 19886 30308 19892 30320
rect 19199 30280 19892 30308
rect 19199 30277 19211 30280
rect 19153 30271 19211 30277
rect 19886 30268 19892 30280
rect 19944 30268 19950 30320
rect 16117 30243 16175 30249
rect 16117 30209 16129 30243
rect 16163 30209 16175 30243
rect 16298 30240 16304 30252
rect 16259 30212 16304 30240
rect 16117 30203 16175 30209
rect 16298 30200 16304 30212
rect 16356 30200 16362 30252
rect 17034 30240 17040 30252
rect 16995 30212 17040 30240
rect 17034 30200 17040 30212
rect 17092 30200 17098 30252
rect 17218 30240 17224 30252
rect 17179 30212 17224 30240
rect 17218 30200 17224 30212
rect 17276 30200 17282 30252
rect 17494 30240 17500 30252
rect 17455 30212 17500 30240
rect 17494 30200 17500 30212
rect 17552 30200 17558 30252
rect 19996 30249 20024 30348
rect 20165 30345 20177 30379
rect 20211 30376 20223 30379
rect 21082 30376 21088 30388
rect 20211 30348 21088 30376
rect 20211 30345 20223 30348
rect 20165 30339 20223 30345
rect 21082 30336 21088 30348
rect 21140 30336 21146 30388
rect 24210 30336 24216 30388
rect 24268 30376 24274 30388
rect 24268 30348 26372 30376
rect 24268 30336 24274 30348
rect 21634 30268 21640 30320
rect 21692 30308 21698 30320
rect 22005 30311 22063 30317
rect 22005 30308 22017 30311
rect 21692 30280 22017 30308
rect 21692 30268 21698 30280
rect 22005 30277 22017 30280
rect 22051 30277 22063 30311
rect 22005 30271 22063 30277
rect 23290 30268 23296 30320
rect 23348 30308 23354 30320
rect 24854 30308 24860 30320
rect 23348 30280 24860 30308
rect 23348 30268 23354 30280
rect 24854 30268 24860 30280
rect 24912 30268 24918 30320
rect 19061 30243 19119 30249
rect 19061 30209 19073 30243
rect 19107 30240 19119 30243
rect 19337 30243 19395 30249
rect 19107 30212 19288 30240
rect 19107 30209 19119 30212
rect 19061 30203 19119 30209
rect 1578 30172 1584 30184
rect 1539 30144 1584 30172
rect 1578 30132 1584 30144
rect 1636 30132 1642 30184
rect 1854 30172 1860 30184
rect 1815 30144 1860 30172
rect 1854 30132 1860 30144
rect 1912 30132 1918 30184
rect 15838 30132 15844 30184
rect 15896 30172 15902 30184
rect 17313 30175 17371 30181
rect 17313 30172 17325 30175
rect 15896 30144 17325 30172
rect 15896 30132 15902 30144
rect 17313 30141 17325 30144
rect 17359 30141 17371 30175
rect 17313 30135 17371 30141
rect 16301 30107 16359 30113
rect 16301 30073 16313 30107
rect 16347 30104 16359 30107
rect 17129 30107 17187 30113
rect 17129 30104 17141 30107
rect 16347 30076 17141 30104
rect 16347 30073 16359 30076
rect 16301 30067 16359 30073
rect 17129 30073 17141 30076
rect 17175 30073 17187 30107
rect 19260 30104 19288 30212
rect 19337 30209 19349 30243
rect 19383 30240 19395 30243
rect 19797 30243 19855 30249
rect 19797 30240 19809 30243
rect 19383 30212 19809 30240
rect 19383 30209 19395 30212
rect 19337 30203 19395 30209
rect 19797 30209 19809 30212
rect 19843 30209 19855 30243
rect 19797 30203 19855 30209
rect 19981 30243 20039 30249
rect 19981 30209 19993 30243
rect 20027 30209 20039 30243
rect 19981 30203 20039 30209
rect 20070 30200 20076 30252
rect 20128 30240 20134 30252
rect 20257 30243 20315 30249
rect 20257 30240 20269 30243
rect 20128 30212 20269 30240
rect 20128 30200 20134 30212
rect 20257 30209 20269 30212
rect 20303 30209 20315 30243
rect 20257 30203 20315 30209
rect 22189 30243 22247 30249
rect 22189 30209 22201 30243
rect 22235 30209 22247 30243
rect 22189 30203 22247 30209
rect 22204 30172 22232 30203
rect 22278 30200 22284 30252
rect 22336 30240 22342 30252
rect 22336 30212 22381 30240
rect 22336 30200 22342 30212
rect 22462 30200 22468 30252
rect 22520 30240 22526 30252
rect 23477 30243 23535 30249
rect 23477 30240 23489 30243
rect 22520 30212 23489 30240
rect 22520 30200 22526 30212
rect 23477 30209 23489 30212
rect 23523 30209 23535 30243
rect 23477 30203 23535 30209
rect 23661 30243 23719 30249
rect 23661 30209 23673 30243
rect 23707 30240 23719 30243
rect 24210 30240 24216 30252
rect 23707 30212 24216 30240
rect 23707 30209 23719 30212
rect 23661 30203 23719 30209
rect 24210 30200 24216 30212
rect 24268 30200 24274 30252
rect 24489 30243 24547 30249
rect 24489 30209 24501 30243
rect 24535 30240 24547 30243
rect 24578 30240 24584 30252
rect 24535 30212 24584 30240
rect 24535 30209 24547 30212
rect 24489 30203 24547 30209
rect 24578 30200 24584 30212
rect 24636 30200 24642 30252
rect 25958 30200 25964 30252
rect 26016 30240 26022 30252
rect 26053 30243 26111 30249
rect 26053 30240 26065 30243
rect 26016 30212 26065 30240
rect 26016 30200 26022 30212
rect 26053 30209 26065 30212
rect 26099 30209 26111 30243
rect 26053 30203 26111 30209
rect 26142 30200 26148 30252
rect 26200 30240 26206 30252
rect 26344 30249 26372 30348
rect 26602 30336 26608 30388
rect 26660 30376 26666 30388
rect 27249 30379 27307 30385
rect 27249 30376 27261 30379
rect 26660 30348 27261 30376
rect 26660 30336 26666 30348
rect 27249 30345 27261 30348
rect 27295 30345 27307 30379
rect 27249 30339 27307 30345
rect 26329 30243 26387 30249
rect 26200 30212 26245 30240
rect 26200 30200 26206 30212
rect 26329 30209 26341 30243
rect 26375 30240 26387 30243
rect 26970 30240 26976 30252
rect 26375 30212 26976 30240
rect 26375 30209 26387 30212
rect 26329 30203 26387 30209
rect 26970 30200 26976 30212
rect 27028 30200 27034 30252
rect 27154 30200 27160 30252
rect 27212 30240 27218 30252
rect 27341 30243 27399 30249
rect 27341 30240 27353 30243
rect 27212 30212 27353 30240
rect 27212 30200 27218 30212
rect 27341 30209 27353 30212
rect 27387 30209 27399 30243
rect 28350 30240 28356 30252
rect 28311 30212 28356 30240
rect 27341 30203 27399 30209
rect 28350 30200 28356 30212
rect 28408 30200 28414 30252
rect 23198 30172 23204 30184
rect 22204 30144 23204 30172
rect 23198 30132 23204 30144
rect 23256 30132 23262 30184
rect 24762 30172 24768 30184
rect 24675 30144 24768 30172
rect 22738 30104 22744 30116
rect 19260 30076 22744 30104
rect 17129 30067 17187 30073
rect 22738 30064 22744 30076
rect 22796 30064 22802 30116
rect 23658 30064 23664 30116
rect 23716 30104 23722 30116
rect 24302 30104 24308 30116
rect 23716 30076 24164 30104
rect 24263 30076 24308 30104
rect 23716 30064 23722 30076
rect 16850 30036 16856 30048
rect 16811 30008 16856 30036
rect 16850 29996 16856 30008
rect 16908 29996 16914 30048
rect 19337 30039 19395 30045
rect 19337 30005 19349 30039
rect 19383 30036 19395 30039
rect 19518 30036 19524 30048
rect 19383 30008 19524 30036
rect 19383 30005 19395 30008
rect 19337 29999 19395 30005
rect 19518 29996 19524 30008
rect 19576 29996 19582 30048
rect 22002 30036 22008 30048
rect 21963 30008 22008 30036
rect 22002 29996 22008 30008
rect 22060 29996 22066 30048
rect 23290 30036 23296 30048
rect 23251 30008 23296 30036
rect 23290 29996 23296 30008
rect 23348 29996 23354 30048
rect 23569 30039 23627 30045
rect 23569 30005 23581 30039
rect 23615 30036 23627 30039
rect 23750 30036 23756 30048
rect 23615 30008 23756 30036
rect 23615 30005 23627 30008
rect 23569 29999 23627 30005
rect 23750 29996 23756 30008
rect 23808 29996 23814 30048
rect 24136 30036 24164 30076
rect 24302 30064 24308 30076
rect 24360 30064 24366 30116
rect 24688 30036 24716 30144
rect 24762 30132 24768 30144
rect 24820 30172 24826 30184
rect 25133 30175 25191 30181
rect 25133 30172 25145 30175
rect 24820 30144 25145 30172
rect 24820 30132 24826 30144
rect 25133 30141 25145 30144
rect 25179 30141 25191 30175
rect 25133 30135 25191 30141
rect 25225 30175 25283 30181
rect 25225 30141 25237 30175
rect 25271 30141 25283 30175
rect 25225 30135 25283 30141
rect 25593 30175 25651 30181
rect 25593 30141 25605 30175
rect 25639 30172 25651 30175
rect 26510 30172 26516 30184
rect 25639 30144 26516 30172
rect 25639 30141 25651 30144
rect 25593 30135 25651 30141
rect 25240 30104 25268 30135
rect 26510 30132 26516 30144
rect 26568 30132 26574 30184
rect 26050 30104 26056 30116
rect 25240 30076 26056 30104
rect 26050 30064 26056 30076
rect 26108 30064 26114 30116
rect 28074 30064 28080 30116
rect 28132 30104 28138 30116
rect 28169 30107 28227 30113
rect 28169 30104 28181 30107
rect 28132 30076 28181 30104
rect 28132 30064 28138 30076
rect 28169 30073 28181 30076
rect 28215 30073 28227 30107
rect 28169 30067 28227 30073
rect 24946 30036 24952 30048
rect 24136 30008 24716 30036
rect 24907 30008 24952 30036
rect 24946 29996 24952 30008
rect 25004 29996 25010 30048
rect 26234 29996 26240 30048
rect 26292 30036 26298 30048
rect 26513 30039 26571 30045
rect 26513 30036 26525 30039
rect 26292 30008 26525 30036
rect 26292 29996 26298 30008
rect 26513 30005 26525 30008
rect 26559 30005 26571 30039
rect 26513 29999 26571 30005
rect 1104 29946 28888 29968
rect 1104 29894 4423 29946
rect 4475 29894 4487 29946
rect 4539 29894 4551 29946
rect 4603 29894 4615 29946
rect 4667 29894 4679 29946
rect 4731 29894 11369 29946
rect 11421 29894 11433 29946
rect 11485 29894 11497 29946
rect 11549 29894 11561 29946
rect 11613 29894 11625 29946
rect 11677 29894 18315 29946
rect 18367 29894 18379 29946
rect 18431 29894 18443 29946
rect 18495 29894 18507 29946
rect 18559 29894 18571 29946
rect 18623 29894 25261 29946
rect 25313 29894 25325 29946
rect 25377 29894 25389 29946
rect 25441 29894 25453 29946
rect 25505 29894 25517 29946
rect 25569 29894 28888 29946
rect 1104 29872 28888 29894
rect 16666 29792 16672 29844
rect 16724 29832 16730 29844
rect 17313 29835 17371 29841
rect 17313 29832 17325 29835
rect 16724 29804 17325 29832
rect 16724 29792 16730 29804
rect 17313 29801 17325 29804
rect 17359 29801 17371 29835
rect 17313 29795 17371 29801
rect 17494 29792 17500 29844
rect 17552 29832 17558 29844
rect 17770 29832 17776 29844
rect 17552 29804 17776 29832
rect 17552 29792 17558 29804
rect 17770 29792 17776 29804
rect 17828 29832 17834 29844
rect 20346 29832 20352 29844
rect 17828 29804 20352 29832
rect 17828 29792 17834 29804
rect 20346 29792 20352 29804
rect 20404 29792 20410 29844
rect 20809 29835 20867 29841
rect 20809 29801 20821 29835
rect 20855 29832 20867 29835
rect 21082 29832 21088 29844
rect 20855 29804 21088 29832
rect 20855 29801 20867 29804
rect 20809 29795 20867 29801
rect 21082 29792 21088 29804
rect 21140 29792 21146 29844
rect 24946 29832 24952 29844
rect 24907 29804 24952 29832
rect 24946 29792 24952 29804
rect 25004 29792 25010 29844
rect 26053 29835 26111 29841
rect 26053 29801 26065 29835
rect 26099 29832 26111 29835
rect 26510 29832 26516 29844
rect 26099 29804 26516 29832
rect 26099 29801 26111 29804
rect 26053 29795 26111 29801
rect 26510 29792 26516 29804
rect 26568 29792 26574 29844
rect 23750 29724 23756 29776
rect 23808 29764 23814 29776
rect 25685 29767 25743 29773
rect 25685 29764 25697 29767
rect 23808 29736 25697 29764
rect 23808 29724 23814 29736
rect 25685 29733 25697 29736
rect 25731 29764 25743 29767
rect 26142 29764 26148 29776
rect 25731 29736 26148 29764
rect 25731 29733 25743 29736
rect 25685 29727 25743 29733
rect 26142 29724 26148 29736
rect 26200 29724 26206 29776
rect 17586 29696 17592 29708
rect 16684 29668 17592 29696
rect 16684 29637 16712 29668
rect 17586 29656 17592 29668
rect 17644 29656 17650 29708
rect 24026 29656 24032 29708
rect 24084 29696 24090 29708
rect 24857 29699 24915 29705
rect 24857 29696 24869 29699
rect 24084 29668 24869 29696
rect 24084 29656 24090 29668
rect 24857 29665 24869 29668
rect 24903 29665 24915 29699
rect 27522 29696 27528 29708
rect 27483 29668 27528 29696
rect 24857 29659 24915 29665
rect 27522 29656 27528 29668
rect 27580 29656 27586 29708
rect 16669 29631 16727 29637
rect 16669 29597 16681 29631
rect 16715 29597 16727 29631
rect 16850 29628 16856 29640
rect 16811 29600 16856 29628
rect 16669 29591 16727 29597
rect 16850 29588 16856 29600
rect 16908 29588 16914 29640
rect 18693 29631 18751 29637
rect 18693 29597 18705 29631
rect 18739 29628 18751 29631
rect 18874 29628 18880 29640
rect 18739 29600 18880 29628
rect 18739 29597 18751 29600
rect 18693 29591 18751 29597
rect 18874 29588 18880 29600
rect 18932 29628 18938 29640
rect 19429 29631 19487 29637
rect 19429 29628 19441 29631
rect 18932 29600 19441 29628
rect 18932 29588 18938 29600
rect 19429 29597 19441 29600
rect 19475 29597 19487 29631
rect 19429 29591 19487 29597
rect 19518 29588 19524 29640
rect 19576 29628 19582 29640
rect 19685 29631 19743 29637
rect 19685 29628 19697 29631
rect 19576 29600 19697 29628
rect 19576 29588 19582 29600
rect 19685 29597 19697 29600
rect 19731 29597 19743 29631
rect 19685 29591 19743 29597
rect 21174 29588 21180 29640
rect 21232 29628 21238 29640
rect 22646 29628 22652 29640
rect 21232 29600 22652 29628
rect 21232 29588 21238 29600
rect 22646 29588 22652 29600
rect 22704 29588 22710 29640
rect 24578 29628 24584 29640
rect 24539 29600 24584 29628
rect 24578 29588 24584 29600
rect 24636 29588 24642 29640
rect 25866 29628 25872 29640
rect 25827 29600 25872 29628
rect 25866 29588 25872 29600
rect 25924 29588 25930 29640
rect 26050 29588 26056 29640
rect 26108 29628 26114 29640
rect 26510 29628 26516 29640
rect 26108 29600 26153 29628
rect 26471 29600 26516 29628
rect 26108 29588 26114 29600
rect 26510 29588 26516 29600
rect 26568 29588 26574 29640
rect 16761 29563 16819 29569
rect 16761 29529 16773 29563
rect 16807 29560 16819 29563
rect 18426 29563 18484 29569
rect 18426 29560 18438 29563
rect 16807 29532 18438 29560
rect 16807 29529 16819 29532
rect 16761 29523 16819 29529
rect 18426 29529 18438 29532
rect 18472 29529 18484 29563
rect 18426 29523 18484 29529
rect 22002 29520 22008 29572
rect 22060 29560 22066 29572
rect 22382 29563 22440 29569
rect 22382 29560 22394 29563
rect 22060 29532 22394 29560
rect 22060 29520 22066 29532
rect 22382 29529 22394 29532
rect 22428 29529 22440 29563
rect 26697 29563 26755 29569
rect 22382 29523 22440 29529
rect 22480 29532 25268 29560
rect 21266 29492 21272 29504
rect 21227 29464 21272 29492
rect 21266 29452 21272 29464
rect 21324 29452 21330 29504
rect 22186 29452 22192 29504
rect 22244 29492 22250 29504
rect 22480 29492 22508 29532
rect 22244 29464 22508 29492
rect 22244 29452 22250 29464
rect 25038 29452 25044 29504
rect 25096 29492 25102 29504
rect 25133 29495 25191 29501
rect 25133 29492 25145 29495
rect 25096 29464 25145 29492
rect 25096 29452 25102 29464
rect 25133 29461 25145 29464
rect 25179 29461 25191 29495
rect 25240 29492 25268 29532
rect 26697 29529 26709 29563
rect 26743 29560 26755 29563
rect 27338 29560 27344 29572
rect 26743 29532 27344 29560
rect 26743 29529 26755 29532
rect 26697 29523 26755 29529
rect 27338 29520 27344 29532
rect 27396 29520 27402 29572
rect 27062 29492 27068 29504
rect 25240 29464 27068 29492
rect 25133 29455 25191 29461
rect 27062 29452 27068 29464
rect 27120 29452 27126 29504
rect 1104 29402 29048 29424
rect 1104 29350 7896 29402
rect 7948 29350 7960 29402
rect 8012 29350 8024 29402
rect 8076 29350 8088 29402
rect 8140 29350 8152 29402
rect 8204 29350 14842 29402
rect 14894 29350 14906 29402
rect 14958 29350 14970 29402
rect 15022 29350 15034 29402
rect 15086 29350 15098 29402
rect 15150 29350 21788 29402
rect 21840 29350 21852 29402
rect 21904 29350 21916 29402
rect 21968 29350 21980 29402
rect 22032 29350 22044 29402
rect 22096 29350 28734 29402
rect 28786 29350 28798 29402
rect 28850 29350 28862 29402
rect 28914 29350 28926 29402
rect 28978 29350 28990 29402
rect 29042 29350 29048 29402
rect 1104 29328 29048 29350
rect 20254 29248 20260 29300
rect 20312 29288 20318 29300
rect 20625 29291 20683 29297
rect 20625 29288 20637 29291
rect 20312 29260 20637 29288
rect 20312 29248 20318 29260
rect 20625 29257 20637 29260
rect 20671 29257 20683 29291
rect 20625 29251 20683 29257
rect 22278 29248 22284 29300
rect 22336 29288 22342 29300
rect 22649 29291 22707 29297
rect 22649 29288 22661 29291
rect 22336 29260 22661 29288
rect 22336 29248 22342 29260
rect 22649 29257 22661 29260
rect 22695 29257 22707 29291
rect 23198 29288 23204 29300
rect 23159 29260 23204 29288
rect 22649 29251 22707 29257
rect 23198 29248 23204 29260
rect 23256 29248 23262 29300
rect 23658 29248 23664 29300
rect 23716 29288 23722 29300
rect 23845 29291 23903 29297
rect 23845 29288 23857 29291
rect 23716 29260 23857 29288
rect 23716 29248 23722 29260
rect 23845 29257 23857 29260
rect 23891 29257 23903 29291
rect 25958 29288 25964 29300
rect 25919 29260 25964 29288
rect 23845 29251 23903 29257
rect 25958 29248 25964 29260
rect 26016 29248 26022 29300
rect 27338 29288 27344 29300
rect 27299 29260 27344 29288
rect 27338 29248 27344 29260
rect 27396 29248 27402 29300
rect 4798 29180 4804 29232
rect 4856 29220 4862 29232
rect 19981 29223 20039 29229
rect 4856 29192 6914 29220
rect 4856 29180 4862 29192
rect 6886 29016 6914 29192
rect 19981 29189 19993 29223
rect 20027 29220 20039 29223
rect 20806 29220 20812 29232
rect 20027 29192 20812 29220
rect 20027 29189 20039 29192
rect 19981 29183 20039 29189
rect 20806 29180 20812 29192
rect 20864 29180 20870 29232
rect 22388 29192 23980 29220
rect 20070 29112 20076 29164
rect 20128 29152 20134 29164
rect 20533 29155 20591 29161
rect 20533 29152 20545 29155
rect 20128 29124 20545 29152
rect 20128 29112 20134 29124
rect 20533 29121 20545 29124
rect 20579 29121 20591 29155
rect 22186 29152 22192 29164
rect 20533 29115 20591 29121
rect 22112 29124 22192 29152
rect 21266 29044 21272 29096
rect 21324 29084 21330 29096
rect 22005 29087 22063 29093
rect 22005 29084 22017 29087
rect 21324 29056 22017 29084
rect 21324 29044 21330 29056
rect 22005 29053 22017 29056
rect 22051 29053 22063 29087
rect 22005 29047 22063 29053
rect 22112 29016 22140 29124
rect 22186 29112 22192 29124
rect 22244 29112 22250 29164
rect 22278 29112 22284 29164
rect 22336 29152 22342 29164
rect 22388 29161 22416 29192
rect 22373 29155 22431 29161
rect 22373 29152 22385 29155
rect 22336 29124 22385 29152
rect 22336 29112 22342 29124
rect 22373 29121 22385 29124
rect 22419 29121 22431 29155
rect 22373 29115 22431 29121
rect 23109 29155 23167 29161
rect 23109 29121 23121 29155
rect 23155 29152 23167 29155
rect 23198 29152 23204 29164
rect 23155 29124 23204 29152
rect 23155 29121 23167 29124
rect 23109 29115 23167 29121
rect 23198 29112 23204 29124
rect 23256 29112 23262 29164
rect 23293 29155 23351 29161
rect 23293 29121 23305 29155
rect 23339 29152 23351 29155
rect 23474 29152 23480 29164
rect 23339 29124 23480 29152
rect 23339 29121 23351 29124
rect 23293 29115 23351 29121
rect 23474 29112 23480 29124
rect 23532 29112 23538 29164
rect 23952 29161 23980 29192
rect 23753 29155 23811 29161
rect 23753 29121 23765 29155
rect 23799 29121 23811 29155
rect 23753 29115 23811 29121
rect 23937 29155 23995 29161
rect 23937 29121 23949 29155
rect 23983 29152 23995 29155
rect 24946 29152 24952 29164
rect 23983 29124 24952 29152
rect 23983 29121 23995 29124
rect 23937 29115 23995 29121
rect 22465 29087 22523 29093
rect 22465 29053 22477 29087
rect 22511 29084 22523 29087
rect 22738 29084 22744 29096
rect 22511 29056 22744 29084
rect 22511 29053 22523 29056
rect 22465 29047 22523 29053
rect 22738 29044 22744 29056
rect 22796 29044 22802 29096
rect 6886 28988 22140 29016
rect 22186 28976 22192 29028
rect 22244 29016 22250 29028
rect 23768 29016 23796 29115
rect 24946 29112 24952 29124
rect 25004 29112 25010 29164
rect 25685 29155 25743 29161
rect 25685 29121 25697 29155
rect 25731 29152 25743 29155
rect 26602 29152 26608 29164
rect 25731 29124 26608 29152
rect 25731 29121 25743 29124
rect 25685 29115 25743 29121
rect 26602 29112 26608 29124
rect 26660 29112 26666 29164
rect 27062 29112 27068 29164
rect 27120 29152 27126 29164
rect 27433 29155 27491 29161
rect 27433 29152 27445 29155
rect 27120 29124 27445 29152
rect 27120 29112 27126 29124
rect 27433 29121 27445 29124
rect 27479 29121 27491 29155
rect 27433 29115 27491 29121
rect 25866 29084 25872 29096
rect 22244 28988 23796 29016
rect 24964 29056 25872 29084
rect 22244 28976 22250 28988
rect 18693 28951 18751 28957
rect 18693 28917 18705 28951
rect 18739 28948 18751 28951
rect 18874 28948 18880 28960
rect 18739 28920 18880 28948
rect 18739 28917 18751 28920
rect 18693 28911 18751 28917
rect 18874 28908 18880 28920
rect 18932 28908 18938 28960
rect 23750 28908 23756 28960
rect 23808 28948 23814 28960
rect 24964 28948 24992 29056
rect 25866 29044 25872 29056
rect 25924 29084 25930 29096
rect 25961 29087 26019 29093
rect 25961 29084 25973 29087
rect 25924 29056 25973 29084
rect 25924 29044 25930 29056
rect 25961 29053 25973 29056
rect 26007 29053 26019 29087
rect 25961 29047 26019 29053
rect 25777 29019 25835 29025
rect 25777 28985 25789 29019
rect 25823 29016 25835 29019
rect 26050 29016 26056 29028
rect 25823 28988 26056 29016
rect 25823 28985 25835 28988
rect 25777 28979 25835 28985
rect 26050 28976 26056 28988
rect 26108 28976 26114 29028
rect 26510 28976 26516 29028
rect 26568 29016 26574 29028
rect 27893 29019 27951 29025
rect 27893 29016 27905 29019
rect 26568 28988 27905 29016
rect 26568 28976 26574 28988
rect 27893 28985 27905 28988
rect 27939 28985 27951 29019
rect 27893 28979 27951 28985
rect 23808 28920 24992 28948
rect 23808 28908 23814 28920
rect 1104 28858 28888 28880
rect 1104 28806 4423 28858
rect 4475 28806 4487 28858
rect 4539 28806 4551 28858
rect 4603 28806 4615 28858
rect 4667 28806 4679 28858
rect 4731 28806 11369 28858
rect 11421 28806 11433 28858
rect 11485 28806 11497 28858
rect 11549 28806 11561 28858
rect 11613 28806 11625 28858
rect 11677 28806 18315 28858
rect 18367 28806 18379 28858
rect 18431 28806 18443 28858
rect 18495 28806 18507 28858
rect 18559 28806 18571 28858
rect 18623 28806 25261 28858
rect 25313 28806 25325 28858
rect 25377 28806 25389 28858
rect 25441 28806 25453 28858
rect 25505 28806 25517 28858
rect 25569 28806 28888 28858
rect 1104 28784 28888 28806
rect 16022 28704 16028 28756
rect 16080 28744 16086 28756
rect 16853 28747 16911 28753
rect 16853 28744 16865 28747
rect 16080 28716 16865 28744
rect 16080 28704 16086 28716
rect 16853 28713 16865 28716
rect 16899 28713 16911 28747
rect 24670 28744 24676 28756
rect 24631 28716 24676 28744
rect 16853 28707 16911 28713
rect 24670 28704 24676 28716
rect 24728 28704 24734 28756
rect 22465 28611 22523 28617
rect 22465 28577 22477 28611
rect 22511 28608 22523 28611
rect 22646 28608 22652 28620
rect 22511 28580 22652 28608
rect 22511 28577 22523 28580
rect 22465 28571 22523 28577
rect 22646 28568 22652 28580
rect 22704 28608 22710 28620
rect 25130 28608 25136 28620
rect 22704 28580 25136 28608
rect 22704 28568 22710 28580
rect 25130 28568 25136 28580
rect 25188 28568 25194 28620
rect 26510 28608 26516 28620
rect 26471 28580 26516 28608
rect 26510 28568 26516 28580
rect 26568 28568 26574 28620
rect 27430 28608 27436 28620
rect 27391 28580 27436 28608
rect 27430 28568 27436 28580
rect 27488 28568 27494 28620
rect 18233 28543 18291 28549
rect 18233 28509 18245 28543
rect 18279 28540 18291 28543
rect 18874 28540 18880 28552
rect 18279 28512 18880 28540
rect 18279 28509 18291 28512
rect 18233 28503 18291 28509
rect 18874 28500 18880 28512
rect 18932 28500 18938 28552
rect 20806 28540 20812 28552
rect 20767 28512 20812 28540
rect 20806 28500 20812 28512
rect 20864 28540 20870 28552
rect 22554 28540 22560 28552
rect 20864 28512 22560 28540
rect 20864 28500 20870 28512
rect 22554 28500 22560 28512
rect 22612 28500 22618 28552
rect 23382 28500 23388 28552
rect 23440 28540 23446 28552
rect 24581 28543 24639 28549
rect 24581 28540 24593 28543
rect 23440 28512 24593 28540
rect 23440 28500 23446 28512
rect 24581 28509 24593 28512
rect 24627 28509 24639 28543
rect 24581 28503 24639 28509
rect 24673 28543 24731 28549
rect 24673 28509 24685 28543
rect 24719 28509 24731 28543
rect 24673 28503 24731 28509
rect 15654 28472 15660 28484
rect 15615 28444 15660 28472
rect 15654 28432 15660 28444
rect 15712 28432 15718 28484
rect 15746 28432 15752 28484
rect 15804 28472 15810 28484
rect 15841 28475 15899 28481
rect 15841 28472 15853 28475
rect 15804 28444 15853 28472
rect 15804 28432 15810 28444
rect 15841 28441 15853 28444
rect 15887 28472 15899 28475
rect 15887 28444 16988 28472
rect 15887 28441 15899 28444
rect 15841 28435 15899 28441
rect 16025 28407 16083 28413
rect 16025 28373 16037 28407
rect 16071 28404 16083 28407
rect 16758 28404 16764 28416
rect 16071 28376 16764 28404
rect 16071 28373 16083 28376
rect 16025 28367 16083 28373
rect 16758 28364 16764 28376
rect 16816 28364 16822 28416
rect 16960 28404 16988 28444
rect 17034 28432 17040 28484
rect 17092 28472 17098 28484
rect 17966 28475 18024 28481
rect 17966 28472 17978 28475
rect 17092 28444 17978 28472
rect 17092 28432 17098 28444
rect 17966 28441 17978 28444
rect 18012 28441 18024 28475
rect 17966 28435 18024 28441
rect 22462 28432 22468 28484
rect 22520 28472 22526 28484
rect 23109 28475 23167 28481
rect 23109 28472 23121 28475
rect 22520 28444 23121 28472
rect 22520 28432 22526 28444
rect 23109 28441 23121 28444
rect 23155 28441 23167 28475
rect 23109 28435 23167 28441
rect 23934 28432 23940 28484
rect 23992 28472 23998 28484
rect 24688 28472 24716 28503
rect 23992 28444 24716 28472
rect 26697 28475 26755 28481
rect 23992 28432 23998 28444
rect 26697 28441 26709 28475
rect 26743 28472 26755 28475
rect 27338 28472 27344 28484
rect 26743 28444 27344 28472
rect 26743 28441 26755 28444
rect 26697 28435 26755 28441
rect 27338 28432 27344 28444
rect 27396 28432 27402 28484
rect 19334 28404 19340 28416
rect 16960 28376 19340 28404
rect 19334 28364 19340 28376
rect 19392 28364 19398 28416
rect 22646 28364 22652 28416
rect 22704 28404 22710 28416
rect 23198 28404 23204 28416
rect 22704 28376 23204 28404
rect 22704 28364 22710 28376
rect 23198 28364 23204 28376
rect 23256 28364 23262 28416
rect 24486 28364 24492 28416
rect 24544 28404 24550 28416
rect 24949 28407 25007 28413
rect 24949 28404 24961 28407
rect 24544 28376 24961 28404
rect 24544 28364 24550 28376
rect 24949 28373 24961 28376
rect 24995 28373 25007 28407
rect 24949 28367 25007 28373
rect 1104 28314 29048 28336
rect 1104 28262 7896 28314
rect 7948 28262 7960 28314
rect 8012 28262 8024 28314
rect 8076 28262 8088 28314
rect 8140 28262 8152 28314
rect 8204 28262 14842 28314
rect 14894 28262 14906 28314
rect 14958 28262 14970 28314
rect 15022 28262 15034 28314
rect 15086 28262 15098 28314
rect 15150 28262 21788 28314
rect 21840 28262 21852 28314
rect 21904 28262 21916 28314
rect 21968 28262 21980 28314
rect 22032 28262 22044 28314
rect 22096 28262 28734 28314
rect 28786 28262 28798 28314
rect 28850 28262 28862 28314
rect 28914 28262 28926 28314
rect 28978 28262 28990 28314
rect 29042 28262 29048 28314
rect 1104 28240 29048 28262
rect 17034 28200 17040 28212
rect 16995 28172 17040 28200
rect 17034 28160 17040 28172
rect 17092 28160 17098 28212
rect 22462 28200 22468 28212
rect 22423 28172 22468 28200
rect 22462 28160 22468 28172
rect 22520 28160 22526 28212
rect 23382 28200 23388 28212
rect 23343 28172 23388 28200
rect 23382 28160 23388 28172
rect 23440 28160 23446 28212
rect 27338 28200 27344 28212
rect 27299 28172 27344 28200
rect 27338 28160 27344 28172
rect 27396 28160 27402 28212
rect 23553 28135 23611 28141
rect 23553 28101 23565 28135
rect 23599 28132 23611 28135
rect 23658 28132 23664 28144
rect 23599 28104 23664 28132
rect 23599 28101 23611 28104
rect 23553 28095 23611 28101
rect 23658 28092 23664 28104
rect 23716 28092 23722 28144
rect 23750 28092 23756 28144
rect 23808 28132 23814 28144
rect 26234 28132 26240 28144
rect 23808 28104 23853 28132
rect 24596 28104 26240 28132
rect 23808 28092 23814 28104
rect 1578 28064 1584 28076
rect 1539 28036 1584 28064
rect 1578 28024 1584 28036
rect 1636 28024 1642 28076
rect 16758 28024 16764 28076
rect 16816 28064 16822 28076
rect 16853 28067 16911 28073
rect 16853 28064 16865 28067
rect 16816 28036 16865 28064
rect 16816 28024 16822 28036
rect 16853 28033 16865 28036
rect 16899 28033 16911 28067
rect 16853 28027 16911 28033
rect 19334 28024 19340 28076
rect 19392 28064 19398 28076
rect 22186 28064 22192 28076
rect 19392 28036 20392 28064
rect 22147 28036 22192 28064
rect 19392 28024 19398 28036
rect 2958 27956 2964 28008
rect 3016 27996 3022 28008
rect 14277 27999 14335 28005
rect 14277 27996 14289 27999
rect 3016 27968 14289 27996
rect 3016 27956 3022 27968
rect 14277 27965 14289 27968
rect 14323 27965 14335 27999
rect 14277 27959 14335 27965
rect 15194 27956 15200 28008
rect 15252 27996 15258 28008
rect 15933 27999 15991 28005
rect 15933 27996 15945 27999
rect 15252 27968 15945 27996
rect 15252 27956 15258 27968
rect 15933 27965 15945 27968
rect 15979 27965 15991 27999
rect 15933 27959 15991 27965
rect 16117 27999 16175 28005
rect 16117 27965 16129 27999
rect 16163 27996 16175 27999
rect 20254 27996 20260 28008
rect 16163 27968 20260 27996
rect 16163 27965 16175 27968
rect 16117 27959 16175 27965
rect 20254 27956 20260 27968
rect 20312 27956 20318 28008
rect 20364 27996 20392 28036
rect 22186 28024 22192 28036
rect 22244 28024 22250 28076
rect 22278 28024 22284 28076
rect 22336 28064 22342 28076
rect 22336 28036 22381 28064
rect 22336 28024 22342 28036
rect 24118 28024 24124 28076
rect 24176 28064 24182 28076
rect 24305 28067 24363 28073
rect 24305 28064 24317 28067
rect 24176 28036 24317 28064
rect 24176 28024 24182 28036
rect 24305 28033 24317 28036
rect 24351 28033 24363 28067
rect 24486 28064 24492 28076
rect 24447 28036 24492 28064
rect 24305 28027 24363 28033
rect 24486 28024 24492 28036
rect 24544 28024 24550 28076
rect 24596 28073 24624 28104
rect 26234 28092 26240 28104
rect 26292 28092 26298 28144
rect 24581 28067 24639 28073
rect 24581 28033 24593 28067
rect 24627 28033 24639 28067
rect 24581 28027 24639 28033
rect 25492 28067 25550 28073
rect 25492 28033 25504 28067
rect 25538 28064 25550 28067
rect 25774 28064 25780 28076
rect 25538 28036 25780 28064
rect 25538 28033 25550 28036
rect 25492 28027 25550 28033
rect 25774 28024 25780 28036
rect 25832 28024 25838 28076
rect 27246 28024 27252 28076
rect 27304 28064 27310 28076
rect 27433 28067 27491 28073
rect 27433 28064 27445 28067
rect 27304 28036 27445 28064
rect 27304 28024 27310 28036
rect 27433 28033 27445 28036
rect 27479 28064 27491 28067
rect 27982 28064 27988 28076
rect 27479 28036 27988 28064
rect 27479 28033 27491 28036
rect 27433 28027 27491 28033
rect 27982 28024 27988 28036
rect 28040 28024 28046 28076
rect 20364 27968 22094 27996
rect 22066 27928 22094 27968
rect 24136 27928 24164 28024
rect 24394 27996 24400 28008
rect 24355 27968 24400 27996
rect 24394 27956 24400 27968
rect 24452 27956 24458 28008
rect 25130 27956 25136 28008
rect 25188 27996 25194 28008
rect 25225 27999 25283 28005
rect 25225 27996 25237 27999
rect 25188 27968 25237 27996
rect 25188 27956 25194 27968
rect 25225 27965 25237 27968
rect 25271 27965 25283 27999
rect 25225 27959 25283 27965
rect 22066 27900 24164 27928
rect 24412 27928 24440 27956
rect 24412 27900 25268 27928
rect 1762 27860 1768 27872
rect 1723 27832 1768 27860
rect 1762 27820 1768 27832
rect 1820 27820 1826 27872
rect 23569 27863 23627 27869
rect 23569 27829 23581 27863
rect 23615 27860 23627 27863
rect 24486 27860 24492 27872
rect 23615 27832 24492 27860
rect 23615 27829 23627 27832
rect 23569 27823 23627 27829
rect 24486 27820 24492 27832
rect 24544 27820 24550 27872
rect 24762 27860 24768 27872
rect 24723 27832 24768 27860
rect 24762 27820 24768 27832
rect 24820 27820 24826 27872
rect 25240 27860 25268 27900
rect 25590 27860 25596 27872
rect 25240 27832 25596 27860
rect 25590 27820 25596 27832
rect 25648 27820 25654 27872
rect 26602 27860 26608 27872
rect 26563 27832 26608 27860
rect 26602 27820 26608 27832
rect 26660 27820 26666 27872
rect 28074 27860 28080 27872
rect 28035 27832 28080 27860
rect 28074 27820 28080 27832
rect 28132 27820 28138 27872
rect 1104 27770 28888 27792
rect 1104 27718 4423 27770
rect 4475 27718 4487 27770
rect 4539 27718 4551 27770
rect 4603 27718 4615 27770
rect 4667 27718 4679 27770
rect 4731 27718 11369 27770
rect 11421 27718 11433 27770
rect 11485 27718 11497 27770
rect 11549 27718 11561 27770
rect 11613 27718 11625 27770
rect 11677 27718 18315 27770
rect 18367 27718 18379 27770
rect 18431 27718 18443 27770
rect 18495 27718 18507 27770
rect 18559 27718 18571 27770
rect 18623 27718 25261 27770
rect 25313 27718 25325 27770
rect 25377 27718 25389 27770
rect 25441 27718 25453 27770
rect 25505 27718 25517 27770
rect 25569 27718 28888 27770
rect 1104 27696 28888 27718
rect 15654 27616 15660 27668
rect 15712 27656 15718 27668
rect 15933 27659 15991 27665
rect 15933 27656 15945 27659
rect 15712 27628 15945 27656
rect 15712 27616 15718 27628
rect 15933 27625 15945 27628
rect 15979 27625 15991 27659
rect 15933 27619 15991 27625
rect 24486 27616 24492 27668
rect 24544 27656 24550 27668
rect 25774 27656 25780 27668
rect 24544 27628 25452 27656
rect 25735 27628 25780 27656
rect 24544 27616 24550 27628
rect 2590 27548 2596 27600
rect 2648 27588 2654 27600
rect 4982 27588 4988 27600
rect 2648 27560 4988 27588
rect 2648 27548 2654 27560
rect 4982 27548 4988 27560
rect 5040 27548 5046 27600
rect 14461 27591 14519 27597
rect 14461 27557 14473 27591
rect 14507 27588 14519 27591
rect 15194 27588 15200 27600
rect 14507 27560 15200 27588
rect 14507 27557 14519 27560
rect 14461 27551 14519 27557
rect 15194 27548 15200 27560
rect 15252 27548 15258 27600
rect 21450 27548 21456 27600
rect 21508 27588 21514 27600
rect 22186 27588 22192 27600
rect 21508 27560 22192 27588
rect 21508 27548 21514 27560
rect 22186 27548 22192 27560
rect 22244 27548 22250 27600
rect 25130 27548 25136 27600
rect 25188 27548 25194 27600
rect 25424 27588 25452 27628
rect 25774 27616 25780 27628
rect 25832 27616 25838 27668
rect 26602 27656 26608 27668
rect 26160 27628 26608 27656
rect 26160 27588 26188 27628
rect 26602 27616 26608 27628
rect 26660 27616 26666 27668
rect 25424 27560 26188 27588
rect 15381 27523 15439 27529
rect 15381 27489 15393 27523
rect 15427 27520 15439 27523
rect 15838 27520 15844 27532
rect 15427 27492 15844 27520
rect 15427 27489 15439 27492
rect 15381 27483 15439 27489
rect 15838 27480 15844 27492
rect 15896 27480 15902 27532
rect 23937 27523 23995 27529
rect 23937 27489 23949 27523
rect 23983 27520 23995 27523
rect 25148 27520 25176 27548
rect 23983 27492 25176 27520
rect 25424 27520 25452 27560
rect 27522 27520 27528 27532
rect 25424 27492 25544 27520
rect 27483 27492 27528 27520
rect 23983 27489 23995 27492
rect 23937 27483 23995 27489
rect 14366 27452 14372 27464
rect 14327 27424 14372 27452
rect 14366 27412 14372 27424
rect 14424 27412 14430 27464
rect 15565 27455 15623 27461
rect 15565 27421 15577 27455
rect 15611 27452 15623 27455
rect 16022 27452 16028 27464
rect 15611 27424 16028 27452
rect 15611 27421 15623 27424
rect 15565 27415 15623 27421
rect 16022 27412 16028 27424
rect 16080 27412 16086 27464
rect 16298 27412 16304 27464
rect 16356 27452 16362 27464
rect 16485 27455 16543 27461
rect 16485 27452 16497 27455
rect 16356 27424 16497 27452
rect 16356 27412 16362 27424
rect 16485 27421 16497 27424
rect 16531 27421 16543 27455
rect 16485 27415 16543 27421
rect 18874 27412 18880 27464
rect 18932 27452 18938 27464
rect 19429 27455 19487 27461
rect 19429 27452 19441 27455
rect 18932 27424 19441 27452
rect 18932 27412 18938 27424
rect 19429 27421 19441 27424
rect 19475 27421 19487 27455
rect 19429 27415 19487 27421
rect 24946 27412 24952 27464
rect 25004 27452 25010 27464
rect 25516 27461 25544 27492
rect 27522 27480 27528 27492
rect 27580 27480 27586 27532
rect 28074 27480 28080 27532
rect 28132 27520 28138 27532
rect 28353 27523 28411 27529
rect 28353 27520 28365 27523
rect 28132 27492 28365 27520
rect 28132 27480 28138 27492
rect 28353 27489 28365 27492
rect 28399 27489 28411 27523
rect 28353 27483 28411 27489
rect 25133 27455 25191 27461
rect 25133 27452 25145 27455
rect 25004 27424 25145 27452
rect 25004 27412 25010 27424
rect 25133 27421 25145 27424
rect 25179 27421 25191 27455
rect 25133 27415 25191 27421
rect 25317 27455 25375 27461
rect 25317 27421 25329 27455
rect 25363 27421 25375 27455
rect 25317 27415 25375 27421
rect 25409 27455 25467 27461
rect 25409 27421 25421 27455
rect 25455 27421 25467 27455
rect 25409 27415 25467 27421
rect 25501 27455 25559 27461
rect 25501 27421 25513 27455
rect 25547 27421 25559 27455
rect 25501 27415 25559 27421
rect 1762 27344 1768 27396
rect 1820 27384 1826 27396
rect 15473 27387 15531 27393
rect 15473 27384 15485 27387
rect 1820 27356 15485 27384
rect 1820 27344 1826 27356
rect 15473 27353 15485 27356
rect 15519 27353 15531 27387
rect 15473 27347 15531 27353
rect 19696 27387 19754 27393
rect 19696 27353 19708 27387
rect 19742 27384 19754 27387
rect 19794 27384 19800 27396
rect 19742 27356 19800 27384
rect 19742 27353 19754 27356
rect 19696 27347 19754 27353
rect 19794 27344 19800 27356
rect 19852 27344 19858 27396
rect 23198 27344 23204 27396
rect 23256 27384 23262 27396
rect 23670 27387 23728 27393
rect 23670 27384 23682 27387
rect 23256 27356 23682 27384
rect 23256 27344 23262 27356
rect 23670 27353 23682 27356
rect 23716 27353 23728 27387
rect 23670 27347 23728 27353
rect 25038 27344 25044 27396
rect 25096 27384 25102 27396
rect 25332 27384 25360 27415
rect 25096 27356 25360 27384
rect 25424 27384 25452 27415
rect 25590 27384 25596 27396
rect 25424 27356 25596 27384
rect 25096 27344 25102 27356
rect 25590 27344 25596 27356
rect 25648 27344 25654 27396
rect 27798 27344 27804 27396
rect 27856 27384 27862 27396
rect 28169 27387 28227 27393
rect 28169 27384 28181 27387
rect 27856 27356 28181 27384
rect 27856 27344 27862 27356
rect 28169 27353 28181 27356
rect 28215 27353 28227 27387
rect 28169 27347 28227 27353
rect 16669 27319 16727 27325
rect 16669 27285 16681 27319
rect 16715 27316 16727 27319
rect 17126 27316 17132 27328
rect 16715 27288 17132 27316
rect 16715 27285 16727 27288
rect 16669 27279 16727 27285
rect 17126 27276 17132 27288
rect 17184 27276 17190 27328
rect 20809 27319 20867 27325
rect 20809 27285 20821 27319
rect 20855 27316 20867 27319
rect 21082 27316 21088 27328
rect 20855 27288 21088 27316
rect 20855 27285 20867 27288
rect 20809 27279 20867 27285
rect 21082 27276 21088 27288
rect 21140 27276 21146 27328
rect 22278 27276 22284 27328
rect 22336 27316 22342 27328
rect 22557 27319 22615 27325
rect 22557 27316 22569 27319
rect 22336 27288 22569 27316
rect 22336 27276 22342 27288
rect 22557 27285 22569 27288
rect 22603 27285 22615 27319
rect 22557 27279 22615 27285
rect 1104 27226 29048 27248
rect 1104 27174 7896 27226
rect 7948 27174 7960 27226
rect 8012 27174 8024 27226
rect 8076 27174 8088 27226
rect 8140 27174 8152 27226
rect 8204 27174 14842 27226
rect 14894 27174 14906 27226
rect 14958 27174 14970 27226
rect 15022 27174 15034 27226
rect 15086 27174 15098 27226
rect 15150 27174 21788 27226
rect 21840 27174 21852 27226
rect 21904 27174 21916 27226
rect 21968 27174 21980 27226
rect 22032 27174 22044 27226
rect 22096 27174 28734 27226
rect 28786 27174 28798 27226
rect 28850 27174 28862 27226
rect 28914 27174 28926 27226
rect 28978 27174 28990 27226
rect 29042 27174 29048 27226
rect 1104 27152 29048 27174
rect 16298 27112 16304 27124
rect 16259 27084 16304 27112
rect 16298 27072 16304 27084
rect 16356 27072 16362 27124
rect 20254 27112 20260 27124
rect 20215 27084 20260 27112
rect 20254 27072 20260 27084
rect 20312 27072 20318 27124
rect 21634 27112 21640 27124
rect 21192 27084 21640 27112
rect 17052 27016 18644 27044
rect 15930 26976 15936 26988
rect 15891 26948 15936 26976
rect 15930 26936 15936 26948
rect 15988 26936 15994 26988
rect 16117 26979 16175 26985
rect 16117 26945 16129 26979
rect 16163 26976 16175 26979
rect 16163 26948 16804 26976
rect 16163 26945 16175 26948
rect 16117 26939 16175 26945
rect 16776 26920 16804 26948
rect 16758 26868 16764 26920
rect 16816 26868 16822 26920
rect 16850 26868 16856 26920
rect 16908 26908 16914 26920
rect 17052 26917 17080 27016
rect 17126 26936 17132 26988
rect 17184 26976 17190 26988
rect 17293 26979 17351 26985
rect 17293 26976 17305 26979
rect 17184 26948 17305 26976
rect 17184 26936 17190 26948
rect 17293 26945 17305 26948
rect 17339 26945 17351 26979
rect 18616 26976 18644 27016
rect 20714 27004 20720 27056
rect 20772 27044 20778 27056
rect 21192 27053 21220 27084
rect 21634 27072 21640 27084
rect 21692 27072 21698 27124
rect 23198 27112 23204 27124
rect 23159 27084 23204 27112
rect 23198 27072 23204 27084
rect 23256 27072 23262 27124
rect 24486 27112 24492 27124
rect 24447 27084 24492 27112
rect 24486 27072 24492 27084
rect 24544 27072 24550 27124
rect 27798 27112 27804 27124
rect 27759 27084 27804 27112
rect 27798 27072 27804 27084
rect 27856 27072 27862 27124
rect 21177 27047 21235 27053
rect 21177 27044 21189 27047
rect 20772 27016 21189 27044
rect 20772 27004 20778 27016
rect 21177 27013 21189 27016
rect 21223 27013 21235 27047
rect 21177 27007 21235 27013
rect 21361 27047 21419 27053
rect 21361 27013 21373 27047
rect 21407 27044 21419 27047
rect 22922 27044 22928 27056
rect 21407 27016 22928 27044
rect 21407 27013 21419 27016
rect 21361 27007 21419 27013
rect 22922 27004 22928 27016
rect 22980 27004 22986 27056
rect 23750 27004 23756 27056
rect 23808 27044 23814 27056
rect 23808 27016 24532 27044
rect 23808 27004 23814 27016
rect 24504 26988 24532 27016
rect 18874 26976 18880 26988
rect 18616 26948 18880 26976
rect 17293 26939 17351 26945
rect 18874 26936 18880 26948
rect 18932 26936 18938 26988
rect 18966 26936 18972 26988
rect 19024 26976 19030 26988
rect 19133 26979 19191 26985
rect 19133 26976 19145 26979
rect 19024 26948 19145 26976
rect 19024 26936 19030 26948
rect 19133 26945 19145 26948
rect 19179 26945 19191 26979
rect 19133 26939 19191 26945
rect 21453 26979 21511 26985
rect 21453 26945 21465 26979
rect 21499 26976 21511 26979
rect 22649 26979 22707 26985
rect 22649 26976 22661 26979
rect 21499 26948 22661 26976
rect 21499 26945 21511 26948
rect 21453 26939 21511 26945
rect 22649 26945 22661 26948
rect 22695 26945 22707 26979
rect 22649 26939 22707 26945
rect 23109 26979 23167 26985
rect 23109 26945 23121 26979
rect 23155 26945 23167 26979
rect 23290 26976 23296 26988
rect 23251 26948 23296 26976
rect 23109 26939 23167 26945
rect 17037 26911 17095 26917
rect 17037 26908 17049 26911
rect 16908 26880 17049 26908
rect 16908 26868 16914 26880
rect 17037 26877 17049 26880
rect 17083 26877 17095 26911
rect 22002 26908 22008 26920
rect 21963 26880 22008 26908
rect 17037 26871 17095 26877
rect 22002 26868 22008 26880
rect 22060 26868 22066 26920
rect 22370 26908 22376 26920
rect 22331 26880 22376 26908
rect 22370 26868 22376 26880
rect 22428 26868 22434 26920
rect 22465 26911 22523 26917
rect 22465 26877 22477 26911
rect 22511 26908 22523 26911
rect 22738 26908 22744 26920
rect 22511 26880 22744 26908
rect 22511 26877 22523 26880
rect 22465 26871 22523 26877
rect 22738 26868 22744 26880
rect 22796 26868 22802 26920
rect 22186 26800 22192 26852
rect 22244 26840 22250 26852
rect 23124 26840 23152 26939
rect 23290 26936 23296 26948
rect 23348 26936 23354 26988
rect 23658 26936 23664 26988
rect 23716 26976 23722 26988
rect 24118 26976 24124 26988
rect 23716 26948 24124 26976
rect 23716 26936 23722 26948
rect 24118 26936 24124 26948
rect 24176 26976 24182 26988
rect 24397 26979 24455 26985
rect 24397 26976 24409 26979
rect 24176 26948 24409 26976
rect 24176 26936 24182 26948
rect 24397 26945 24409 26948
rect 24443 26945 24455 26979
rect 24397 26939 24455 26945
rect 24486 26936 24492 26988
rect 24544 26976 24550 26988
rect 24673 26979 24731 26985
rect 24673 26976 24685 26979
rect 24544 26948 24685 26976
rect 24544 26936 24550 26948
rect 24673 26945 24685 26948
rect 24719 26945 24731 26979
rect 27706 26976 27712 26988
rect 27619 26948 27712 26976
rect 24673 26939 24731 26945
rect 27706 26936 27712 26948
rect 27764 26976 27770 26988
rect 28258 26976 28264 26988
rect 27764 26948 28264 26976
rect 27764 26936 27770 26948
rect 28258 26936 28264 26948
rect 28316 26936 28322 26988
rect 24670 26840 24676 26852
rect 22244 26812 23152 26840
rect 24631 26812 24676 26840
rect 22244 26800 22250 26812
rect 24670 26800 24676 26812
rect 24728 26800 24734 26852
rect 18230 26732 18236 26784
rect 18288 26772 18294 26784
rect 18417 26775 18475 26781
rect 18417 26772 18429 26775
rect 18288 26744 18429 26772
rect 18288 26732 18294 26744
rect 18417 26741 18429 26744
rect 18463 26772 18475 26775
rect 19610 26772 19616 26784
rect 18463 26744 19616 26772
rect 18463 26741 18475 26744
rect 18417 26735 18475 26741
rect 19610 26732 19616 26744
rect 19668 26732 19674 26784
rect 21174 26772 21180 26784
rect 21135 26744 21180 26772
rect 21174 26732 21180 26744
rect 21232 26732 21238 26784
rect 1104 26682 28888 26704
rect 1104 26630 4423 26682
rect 4475 26630 4487 26682
rect 4539 26630 4551 26682
rect 4603 26630 4615 26682
rect 4667 26630 4679 26682
rect 4731 26630 11369 26682
rect 11421 26630 11433 26682
rect 11485 26630 11497 26682
rect 11549 26630 11561 26682
rect 11613 26630 11625 26682
rect 11677 26630 18315 26682
rect 18367 26630 18379 26682
rect 18431 26630 18443 26682
rect 18495 26630 18507 26682
rect 18559 26630 18571 26682
rect 18623 26630 25261 26682
rect 25313 26630 25325 26682
rect 25377 26630 25389 26682
rect 25441 26630 25453 26682
rect 25505 26630 25517 26682
rect 25569 26630 28888 26682
rect 1104 26608 28888 26630
rect 15930 26528 15936 26580
rect 15988 26568 15994 26580
rect 16209 26571 16267 26577
rect 16209 26568 16221 26571
rect 15988 26540 16221 26568
rect 15988 26528 15994 26540
rect 16209 26537 16221 26540
rect 16255 26537 16267 26571
rect 19794 26568 19800 26580
rect 19755 26540 19800 26568
rect 16209 26531 16267 26537
rect 19794 26528 19800 26540
rect 19852 26528 19858 26580
rect 20898 26528 20904 26580
rect 20956 26568 20962 26580
rect 22002 26568 22008 26580
rect 20956 26540 22008 26568
rect 20956 26528 20962 26540
rect 22002 26528 22008 26540
rect 22060 26528 22066 26580
rect 24026 26568 24032 26580
rect 23987 26540 24032 26568
rect 24026 26528 24032 26540
rect 24084 26568 24090 26580
rect 24670 26568 24676 26580
rect 24084 26540 24676 26568
rect 24084 26528 24090 26540
rect 24670 26528 24676 26540
rect 24728 26528 24734 26580
rect 24118 26460 24124 26512
rect 24176 26500 24182 26512
rect 24857 26503 24915 26509
rect 24857 26500 24869 26503
rect 24176 26472 24869 26500
rect 24176 26460 24182 26472
rect 24857 26469 24869 26472
rect 24903 26469 24915 26503
rect 24857 26463 24915 26469
rect 15470 26392 15476 26444
rect 15528 26432 15534 26444
rect 15565 26435 15623 26441
rect 15565 26432 15577 26435
rect 15528 26404 15577 26432
rect 15528 26392 15534 26404
rect 15565 26401 15577 26404
rect 15611 26401 15623 26435
rect 15565 26395 15623 26401
rect 18874 26392 18880 26444
rect 18932 26432 18938 26444
rect 20625 26435 20683 26441
rect 20625 26432 20637 26435
rect 18932 26404 20637 26432
rect 18932 26392 18938 26404
rect 20625 26401 20637 26404
rect 20671 26401 20683 26435
rect 24581 26435 24639 26441
rect 24581 26432 24593 26435
rect 20625 26395 20683 26401
rect 23952 26404 24593 26432
rect 23952 26376 23980 26404
rect 24581 26401 24593 26404
rect 24627 26401 24639 26435
rect 24581 26395 24639 26401
rect 2225 26367 2283 26373
rect 2225 26333 2237 26367
rect 2271 26364 2283 26367
rect 2590 26364 2596 26376
rect 2271 26336 2596 26364
rect 2271 26333 2283 26336
rect 2225 26327 2283 26333
rect 2590 26324 2596 26336
rect 2648 26324 2654 26376
rect 15841 26367 15899 26373
rect 15841 26333 15853 26367
rect 15887 26364 15899 26367
rect 18230 26364 18236 26376
rect 15887 26336 18236 26364
rect 15887 26333 15899 26336
rect 15841 26327 15899 26333
rect 18230 26324 18236 26336
rect 18288 26324 18294 26376
rect 19978 26364 19984 26376
rect 19939 26336 19984 26364
rect 19978 26324 19984 26336
rect 20036 26324 20042 26376
rect 20892 26367 20950 26373
rect 20892 26333 20904 26367
rect 20938 26364 20950 26367
rect 21174 26364 21180 26376
rect 20938 26336 21180 26364
rect 20938 26333 20950 26336
rect 20892 26327 20950 26333
rect 21174 26324 21180 26336
rect 21232 26324 21238 26376
rect 23845 26367 23903 26373
rect 23845 26333 23857 26367
rect 23891 26364 23903 26367
rect 23934 26364 23940 26376
rect 23891 26336 23940 26364
rect 23891 26333 23903 26336
rect 23845 26327 23903 26333
rect 23934 26324 23940 26336
rect 23992 26324 23998 26376
rect 24029 26367 24087 26373
rect 24029 26333 24041 26367
rect 24075 26364 24087 26367
rect 24118 26364 24124 26376
rect 24075 26336 24124 26364
rect 24075 26333 24087 26336
rect 24029 26327 24087 26333
rect 24118 26324 24124 26336
rect 24176 26324 24182 26376
rect 25130 26324 25136 26376
rect 25188 26364 25194 26376
rect 27341 26367 27399 26373
rect 27341 26364 27353 26367
rect 25188 26336 27353 26364
rect 25188 26324 25194 26336
rect 27341 26333 27353 26336
rect 27387 26333 27399 26367
rect 27341 26327 27399 26333
rect 15746 26296 15752 26308
rect 15707 26268 15752 26296
rect 15746 26256 15752 26268
rect 15804 26256 15810 26308
rect 26234 26256 26240 26308
rect 26292 26296 26298 26308
rect 27074 26299 27132 26305
rect 27074 26296 27086 26299
rect 26292 26268 27086 26296
rect 26292 26256 26298 26268
rect 27074 26265 27086 26268
rect 27120 26265 27132 26299
rect 27074 26259 27132 26265
rect 1854 26188 1860 26240
rect 1912 26228 1918 26240
rect 2133 26231 2191 26237
rect 2133 26228 2145 26231
rect 1912 26200 2145 26228
rect 1912 26188 1918 26200
rect 2133 26197 2145 26200
rect 2179 26197 2191 26231
rect 2133 26191 2191 26197
rect 25041 26231 25099 26237
rect 25041 26197 25053 26231
rect 25087 26228 25099 26231
rect 25498 26228 25504 26240
rect 25087 26200 25504 26228
rect 25087 26197 25099 26200
rect 25041 26191 25099 26197
rect 25498 26188 25504 26200
rect 25556 26188 25562 26240
rect 25958 26228 25964 26240
rect 25919 26200 25964 26228
rect 25958 26188 25964 26200
rect 26016 26188 26022 26240
rect 1104 26138 29048 26160
rect 1104 26086 7896 26138
rect 7948 26086 7960 26138
rect 8012 26086 8024 26138
rect 8076 26086 8088 26138
rect 8140 26086 8152 26138
rect 8204 26086 14842 26138
rect 14894 26086 14906 26138
rect 14958 26086 14970 26138
rect 15022 26086 15034 26138
rect 15086 26086 15098 26138
rect 15150 26086 21788 26138
rect 21840 26086 21852 26138
rect 21904 26086 21916 26138
rect 21968 26086 21980 26138
rect 22032 26086 22044 26138
rect 22096 26086 28734 26138
rect 28786 26086 28798 26138
rect 28850 26086 28862 26138
rect 28914 26086 28926 26138
rect 28978 26086 28990 26138
rect 29042 26086 29048 26138
rect 1104 26064 29048 26086
rect 16301 26027 16359 26033
rect 16301 25993 16313 26027
rect 16347 25993 16359 26027
rect 16301 25987 16359 25993
rect 1854 25956 1860 25968
rect 1815 25928 1860 25956
rect 1854 25916 1860 25928
rect 1912 25916 1918 25968
rect 16316 25956 16344 25987
rect 16482 25984 16488 26036
rect 16540 26024 16546 26036
rect 18233 26027 18291 26033
rect 18233 26024 18245 26027
rect 16540 25996 18245 26024
rect 16540 25984 16546 25996
rect 18233 25993 18245 25996
rect 18279 26024 18291 26027
rect 19702 26024 19708 26036
rect 18279 25996 19708 26024
rect 18279 25993 18291 25996
rect 18233 25987 18291 25993
rect 19702 25984 19708 25996
rect 19760 25984 19766 26036
rect 19797 26027 19855 26033
rect 19797 25993 19809 26027
rect 19843 26024 19855 26027
rect 19978 26024 19984 26036
rect 19843 25996 19984 26024
rect 19843 25993 19855 25996
rect 19797 25987 19855 25993
rect 19978 25984 19984 25996
rect 20036 25984 20042 26036
rect 22922 26024 22928 26036
rect 22883 25996 22928 26024
rect 22922 25984 22928 25996
rect 22980 25984 22986 26036
rect 25133 26027 25191 26033
rect 25133 25993 25145 26027
rect 25179 26024 25191 26027
rect 25590 26024 25596 26036
rect 25179 25996 25596 26024
rect 25179 25993 25191 25996
rect 25133 25987 25191 25993
rect 25590 25984 25596 25996
rect 25648 25984 25654 26036
rect 27062 25984 27068 26036
rect 27120 26024 27126 26036
rect 27430 26024 27436 26036
rect 27120 25996 27436 26024
rect 27120 25984 27126 25996
rect 27430 25984 27436 25996
rect 27488 25984 27494 26036
rect 17098 25959 17156 25965
rect 17098 25956 17110 25959
rect 16316 25928 17110 25956
rect 17098 25925 17110 25928
rect 17144 25925 17156 25959
rect 17098 25919 17156 25925
rect 22848 25928 23520 25956
rect 16114 25888 16120 25900
rect 16075 25860 16120 25888
rect 16114 25848 16120 25860
rect 16172 25848 16178 25900
rect 19978 25888 19984 25900
rect 19939 25860 19984 25888
rect 19978 25848 19984 25860
rect 20036 25848 20042 25900
rect 20162 25888 20168 25900
rect 20123 25860 20168 25888
rect 20162 25848 20168 25860
rect 20220 25848 20226 25900
rect 22646 25848 22652 25900
rect 22704 25888 22710 25900
rect 22848 25897 22876 25928
rect 23492 25897 23520 25928
rect 23676 25928 26004 25956
rect 23676 25897 23704 25928
rect 25976 25900 26004 25928
rect 26050 25916 26056 25968
rect 26108 25956 26114 25968
rect 26605 25959 26663 25965
rect 26605 25956 26617 25959
rect 26108 25928 26617 25956
rect 26108 25916 26114 25928
rect 26605 25925 26617 25928
rect 26651 25956 26663 25959
rect 26651 25928 27384 25956
rect 26651 25925 26663 25928
rect 26605 25919 26663 25925
rect 22833 25891 22891 25897
rect 22833 25888 22845 25891
rect 22704 25860 22845 25888
rect 22704 25848 22710 25860
rect 22833 25857 22845 25860
rect 22879 25857 22891 25891
rect 22833 25851 22891 25857
rect 23017 25891 23075 25897
rect 23017 25857 23029 25891
rect 23063 25857 23075 25891
rect 23017 25851 23075 25857
rect 23477 25891 23535 25897
rect 23477 25857 23489 25891
rect 23523 25857 23535 25891
rect 23477 25851 23535 25857
rect 23661 25891 23719 25897
rect 23661 25857 23673 25891
rect 23707 25857 23719 25891
rect 23661 25851 23719 25857
rect 25317 25891 25375 25897
rect 25317 25857 25329 25891
rect 25363 25857 25375 25891
rect 25498 25888 25504 25900
rect 25459 25860 25504 25888
rect 25317 25851 25375 25857
rect 1670 25820 1676 25832
rect 1631 25792 1676 25820
rect 1670 25780 1676 25792
rect 1728 25780 1734 25832
rect 2774 25820 2780 25832
rect 2735 25792 2780 25820
rect 2774 25780 2780 25792
rect 2832 25780 2838 25832
rect 16850 25820 16856 25832
rect 16811 25792 16856 25820
rect 16850 25780 16856 25792
rect 16908 25780 16914 25832
rect 23032 25820 23060 25851
rect 25332 25820 25360 25851
rect 25498 25848 25504 25860
rect 25556 25848 25562 25900
rect 25958 25848 25964 25900
rect 26016 25888 26022 25900
rect 26421 25891 26479 25897
rect 26421 25888 26433 25891
rect 26016 25860 26433 25888
rect 26016 25848 26022 25860
rect 26421 25857 26433 25860
rect 26467 25857 26479 25891
rect 26421 25851 26479 25857
rect 26970 25848 26976 25900
rect 27028 25888 27034 25900
rect 27356 25897 27384 25928
rect 27157 25891 27215 25897
rect 27157 25888 27169 25891
rect 27028 25860 27169 25888
rect 27028 25848 27034 25860
rect 27157 25857 27169 25860
rect 27203 25857 27215 25891
rect 27157 25851 27215 25857
rect 27341 25891 27399 25897
rect 27341 25857 27353 25891
rect 27387 25857 27399 25891
rect 27341 25851 27399 25857
rect 25593 25823 25651 25829
rect 23032 25792 23704 25820
rect 25332 25792 25452 25820
rect 23676 25764 23704 25792
rect 23569 25755 23627 25761
rect 23569 25752 23581 25755
rect 22066 25724 23581 25752
rect 21726 25644 21732 25696
rect 21784 25684 21790 25696
rect 22066 25684 22094 25724
rect 23569 25721 23581 25724
rect 23615 25721 23627 25755
rect 23569 25715 23627 25721
rect 23658 25712 23664 25764
rect 23716 25712 23722 25764
rect 21784 25656 22094 25684
rect 25424 25684 25452 25792
rect 25593 25789 25605 25823
rect 25639 25789 25651 25823
rect 26142 25820 26148 25832
rect 26103 25792 26148 25820
rect 25593 25783 25651 25789
rect 25608 25752 25636 25783
rect 26142 25780 26148 25792
rect 26200 25780 26206 25832
rect 25866 25752 25872 25764
rect 25608 25724 25872 25752
rect 25866 25712 25872 25724
rect 25924 25752 25930 25764
rect 27157 25755 27215 25761
rect 27157 25752 27169 25755
rect 25924 25724 27169 25752
rect 25924 25712 25930 25724
rect 27157 25721 27169 25724
rect 27203 25721 27215 25755
rect 27157 25715 27215 25721
rect 25682 25684 25688 25696
rect 25424 25656 25688 25684
rect 21784 25644 21790 25656
rect 25682 25644 25688 25656
rect 25740 25644 25746 25696
rect 25774 25644 25780 25696
rect 25832 25684 25838 25696
rect 26237 25687 26295 25693
rect 26237 25684 26249 25687
rect 25832 25656 26249 25684
rect 25832 25644 25838 25656
rect 26237 25653 26249 25656
rect 26283 25653 26295 25687
rect 26237 25647 26295 25653
rect 1104 25594 28888 25616
rect 1104 25542 4423 25594
rect 4475 25542 4487 25594
rect 4539 25542 4551 25594
rect 4603 25542 4615 25594
rect 4667 25542 4679 25594
rect 4731 25542 11369 25594
rect 11421 25542 11433 25594
rect 11485 25542 11497 25594
rect 11549 25542 11561 25594
rect 11613 25542 11625 25594
rect 11677 25542 18315 25594
rect 18367 25542 18379 25594
rect 18431 25542 18443 25594
rect 18495 25542 18507 25594
rect 18559 25542 18571 25594
rect 18623 25542 25261 25594
rect 25313 25542 25325 25594
rect 25377 25542 25389 25594
rect 25441 25542 25453 25594
rect 25505 25542 25517 25594
rect 25569 25542 28888 25594
rect 1104 25520 28888 25542
rect 1670 25480 1676 25492
rect 1631 25452 1676 25480
rect 1670 25440 1676 25452
rect 1728 25440 1734 25492
rect 16114 25440 16120 25492
rect 16172 25480 16178 25492
rect 17037 25483 17095 25489
rect 17037 25480 17049 25483
rect 16172 25452 17049 25480
rect 16172 25440 16178 25452
rect 17037 25449 17049 25452
rect 17083 25449 17095 25483
rect 17037 25443 17095 25449
rect 18509 25483 18567 25489
rect 18509 25449 18521 25483
rect 18555 25480 18567 25483
rect 18966 25480 18972 25492
rect 18555 25452 18972 25480
rect 18555 25449 18567 25452
rect 18509 25443 18567 25449
rect 18966 25440 18972 25452
rect 19024 25440 19030 25492
rect 25777 25483 25835 25489
rect 25777 25449 25789 25483
rect 25823 25480 25835 25483
rect 26234 25480 26240 25492
rect 25823 25452 26240 25480
rect 25823 25449 25835 25452
rect 25777 25443 25835 25449
rect 26234 25440 26240 25452
rect 26292 25440 26298 25492
rect 21545 25415 21603 25421
rect 21545 25381 21557 25415
rect 21591 25412 21603 25415
rect 22370 25412 22376 25424
rect 21591 25384 22376 25412
rect 21591 25381 21603 25384
rect 21545 25375 21603 25381
rect 22370 25372 22376 25384
rect 22428 25372 22434 25424
rect 15470 25304 15476 25356
rect 15528 25344 15534 25356
rect 15565 25347 15623 25353
rect 15565 25344 15577 25347
rect 15528 25316 15577 25344
rect 15528 25304 15534 25316
rect 15565 25313 15577 25316
rect 15611 25313 15623 25347
rect 15565 25307 15623 25313
rect 24946 25304 24952 25356
rect 25004 25344 25010 25356
rect 25317 25347 25375 25353
rect 25317 25344 25329 25347
rect 25004 25316 25329 25344
rect 25004 25304 25010 25316
rect 25317 25313 25329 25316
rect 25363 25313 25375 25347
rect 25317 25307 25375 25313
rect 25409 25347 25467 25353
rect 25409 25313 25421 25347
rect 25455 25344 25467 25347
rect 25682 25344 25688 25356
rect 25455 25316 25688 25344
rect 25455 25313 25467 25316
rect 25409 25307 25467 25313
rect 25682 25304 25688 25316
rect 25740 25304 25746 25356
rect 26513 25347 26571 25353
rect 26513 25313 26525 25347
rect 26559 25344 26571 25347
rect 27706 25344 27712 25356
rect 26559 25316 27712 25344
rect 26559 25313 26571 25316
rect 26513 25307 26571 25313
rect 27706 25304 27712 25316
rect 27764 25304 27770 25356
rect 15841 25279 15899 25285
rect 15841 25245 15853 25279
rect 15887 25276 15899 25279
rect 16482 25276 16488 25288
rect 15887 25248 16488 25276
rect 15887 25245 15899 25248
rect 15841 25239 15899 25245
rect 16482 25236 16488 25248
rect 16540 25236 16546 25288
rect 18230 25236 18236 25288
rect 18288 25276 18294 25288
rect 18509 25279 18567 25285
rect 18509 25276 18521 25279
rect 18288 25248 18521 25276
rect 18288 25236 18294 25248
rect 18509 25245 18521 25248
rect 18555 25245 18567 25279
rect 18509 25239 18567 25245
rect 18693 25279 18751 25285
rect 18693 25245 18705 25279
rect 18739 25276 18751 25279
rect 20714 25276 20720 25288
rect 18739 25248 20720 25276
rect 18739 25245 18751 25248
rect 18693 25239 18751 25245
rect 16669 25211 16727 25217
rect 16669 25177 16681 25211
rect 16715 25177 16727 25211
rect 16669 25171 16727 25177
rect 9490 25100 9496 25152
rect 9548 25140 9554 25152
rect 15749 25143 15807 25149
rect 15749 25140 15761 25143
rect 9548 25112 15761 25140
rect 9548 25100 9554 25112
rect 15749 25109 15761 25112
rect 15795 25109 15807 25143
rect 15749 25103 15807 25109
rect 16209 25143 16267 25149
rect 16209 25109 16221 25143
rect 16255 25140 16267 25143
rect 16684 25140 16712 25171
rect 16758 25168 16764 25220
rect 16816 25208 16822 25220
rect 16853 25211 16911 25217
rect 16853 25208 16865 25211
rect 16816 25180 16865 25208
rect 16816 25168 16822 25180
rect 16853 25177 16865 25180
rect 16899 25208 16911 25211
rect 17126 25208 17132 25220
rect 16899 25180 17132 25208
rect 16899 25177 16911 25180
rect 16853 25171 16911 25177
rect 17126 25168 17132 25180
rect 17184 25208 17190 25220
rect 18708 25208 18736 25239
rect 20714 25236 20720 25248
rect 20772 25276 20778 25288
rect 21450 25276 21456 25288
rect 20772 25248 21456 25276
rect 20772 25236 20778 25248
rect 21450 25236 21456 25248
rect 21508 25276 21514 25288
rect 21545 25279 21603 25285
rect 21545 25276 21557 25279
rect 21508 25248 21557 25276
rect 21508 25236 21514 25248
rect 21545 25245 21557 25248
rect 21591 25245 21603 25279
rect 21726 25276 21732 25288
rect 21687 25248 21732 25276
rect 21545 25239 21603 25245
rect 21726 25236 21732 25248
rect 21784 25236 21790 25288
rect 21821 25279 21879 25285
rect 21821 25245 21833 25279
rect 21867 25276 21879 25279
rect 22830 25276 22836 25288
rect 21867 25248 22836 25276
rect 21867 25245 21879 25248
rect 21821 25239 21879 25245
rect 22830 25236 22836 25248
rect 22888 25236 22894 25288
rect 24029 25279 24087 25285
rect 24029 25245 24041 25279
rect 24075 25276 24087 25279
rect 24854 25276 24860 25288
rect 24075 25248 24860 25276
rect 24075 25245 24087 25248
rect 24029 25239 24087 25245
rect 24854 25236 24860 25248
rect 24912 25236 24918 25288
rect 25038 25276 25044 25288
rect 24951 25248 25044 25276
rect 25038 25236 25044 25248
rect 25096 25236 25102 25288
rect 25222 25276 25228 25288
rect 25183 25248 25228 25276
rect 25222 25236 25228 25248
rect 25280 25236 25286 25288
rect 25590 25236 25596 25288
rect 25648 25276 25654 25288
rect 25958 25276 25964 25288
rect 25648 25248 25964 25276
rect 25648 25236 25654 25248
rect 25958 25236 25964 25248
rect 26016 25236 26022 25288
rect 17184 25180 18736 25208
rect 17184 25168 17190 25180
rect 24210 25168 24216 25220
rect 24268 25208 24274 25220
rect 25056 25208 25084 25236
rect 26694 25208 26700 25220
rect 24268 25180 25084 25208
rect 26655 25180 26700 25208
rect 24268 25168 24274 25180
rect 26694 25168 26700 25180
rect 26752 25168 26758 25220
rect 28350 25208 28356 25220
rect 28311 25180 28356 25208
rect 28350 25168 28356 25180
rect 28408 25168 28414 25220
rect 22554 25140 22560 25152
rect 16255 25112 16712 25140
rect 22515 25112 22560 25140
rect 16255 25109 16267 25112
rect 16209 25103 16267 25109
rect 22554 25100 22560 25112
rect 22612 25100 22618 25152
rect 1104 25050 29048 25072
rect 1104 24998 7896 25050
rect 7948 24998 7960 25050
rect 8012 24998 8024 25050
rect 8076 24998 8088 25050
rect 8140 24998 8152 25050
rect 8204 24998 14842 25050
rect 14894 24998 14906 25050
rect 14958 24998 14970 25050
rect 15022 24998 15034 25050
rect 15086 24998 15098 25050
rect 15150 24998 21788 25050
rect 21840 24998 21852 25050
rect 21904 24998 21916 25050
rect 21968 24998 21980 25050
rect 22032 24998 22044 25050
rect 22096 24998 28734 25050
rect 28786 24998 28798 25050
rect 28850 24998 28862 25050
rect 28914 24998 28926 25050
rect 28978 24998 28990 25050
rect 29042 24998 29048 25050
rect 1104 24976 29048 24998
rect 19978 24896 19984 24948
rect 20036 24936 20042 24948
rect 20533 24939 20591 24945
rect 20533 24936 20545 24939
rect 20036 24908 20545 24936
rect 20036 24896 20042 24908
rect 20533 24905 20545 24908
rect 20579 24905 20591 24939
rect 20533 24899 20591 24905
rect 25222 24896 25228 24948
rect 25280 24936 25286 24948
rect 25409 24939 25467 24945
rect 25409 24936 25421 24939
rect 25280 24908 25421 24936
rect 25280 24896 25286 24908
rect 25409 24905 25421 24908
rect 25455 24905 25467 24939
rect 25409 24899 25467 24905
rect 26694 24896 26700 24948
rect 26752 24936 26758 24948
rect 27249 24939 27307 24945
rect 27249 24936 27261 24939
rect 26752 24908 27261 24936
rect 26752 24896 26758 24908
rect 27249 24905 27261 24908
rect 27295 24905 27307 24939
rect 27249 24899 27307 24905
rect 20901 24871 20959 24877
rect 20901 24837 20913 24871
rect 20947 24868 20959 24871
rect 21082 24868 21088 24880
rect 20947 24840 21088 24868
rect 20947 24837 20959 24840
rect 20901 24831 20959 24837
rect 21082 24828 21088 24840
rect 21140 24868 21146 24880
rect 21542 24868 21548 24880
rect 21140 24840 21548 24868
rect 21140 24828 21146 24840
rect 21542 24828 21548 24840
rect 21600 24828 21606 24880
rect 26142 24868 26148 24880
rect 23768 24840 24532 24868
rect 1578 24800 1584 24812
rect 1539 24772 1584 24800
rect 1578 24760 1584 24772
rect 1636 24760 1642 24812
rect 16850 24760 16856 24812
rect 16908 24800 16914 24812
rect 17405 24803 17463 24809
rect 17405 24800 17417 24803
rect 16908 24772 17417 24800
rect 16908 24760 16914 24772
rect 17405 24769 17417 24772
rect 17451 24769 17463 24803
rect 17405 24763 17463 24769
rect 17494 24760 17500 24812
rect 17552 24800 17558 24812
rect 17661 24803 17719 24809
rect 17661 24800 17673 24803
rect 17552 24772 17673 24800
rect 17552 24760 17558 24772
rect 17661 24769 17673 24772
rect 17707 24769 17719 24803
rect 17661 24763 17719 24769
rect 19889 24803 19947 24809
rect 19889 24769 19901 24803
rect 19935 24800 19947 24803
rect 20438 24800 20444 24812
rect 19935 24772 20444 24800
rect 19935 24769 19947 24772
rect 19889 24763 19947 24769
rect 20438 24760 20444 24772
rect 20496 24760 20502 24812
rect 20993 24803 21051 24809
rect 20993 24769 21005 24803
rect 21039 24800 21051 24803
rect 21634 24800 21640 24812
rect 21039 24772 21640 24800
rect 21039 24769 21051 24772
rect 20993 24763 21051 24769
rect 21634 24760 21640 24772
rect 21692 24800 21698 24812
rect 22189 24803 22247 24809
rect 22189 24800 22201 24803
rect 21692 24772 22201 24800
rect 21692 24760 21698 24772
rect 22189 24769 22201 24772
rect 22235 24769 22247 24803
rect 22189 24763 22247 24769
rect 22462 24760 22468 24812
rect 22520 24800 22526 24812
rect 22557 24803 22615 24809
rect 22557 24800 22569 24803
rect 22520 24772 22569 24800
rect 22520 24760 22526 24772
rect 22557 24769 22569 24772
rect 22603 24769 22615 24803
rect 22830 24800 22836 24812
rect 22791 24772 22836 24800
rect 22557 24763 22615 24769
rect 22830 24760 22836 24772
rect 22888 24760 22894 24812
rect 23768 24809 23796 24840
rect 23753 24803 23811 24809
rect 23753 24769 23765 24803
rect 23799 24769 23811 24803
rect 23753 24763 23811 24769
rect 23845 24803 23903 24809
rect 23845 24769 23857 24803
rect 23891 24800 23903 24803
rect 24026 24800 24032 24812
rect 23891 24772 24032 24800
rect 23891 24769 23903 24772
rect 23845 24763 23903 24769
rect 24026 24760 24032 24772
rect 24084 24760 24090 24812
rect 24504 24809 24532 24840
rect 25700 24840 26148 24868
rect 24489 24803 24547 24809
rect 24489 24769 24501 24803
rect 24535 24800 24547 24803
rect 25590 24800 25596 24812
rect 24535 24772 25596 24800
rect 24535 24769 24547 24772
rect 24489 24763 24547 24769
rect 25590 24760 25596 24772
rect 25648 24760 25654 24812
rect 25700 24809 25728 24840
rect 26142 24828 26148 24840
rect 26200 24828 26206 24880
rect 25685 24803 25743 24809
rect 25685 24769 25697 24803
rect 25731 24769 25743 24803
rect 25866 24800 25872 24812
rect 25827 24772 25872 24800
rect 25685 24763 25743 24769
rect 25866 24760 25872 24772
rect 25924 24760 25930 24812
rect 26878 24760 26884 24812
rect 26936 24800 26942 24812
rect 27062 24800 27068 24812
rect 26936 24772 27068 24800
rect 26936 24760 26942 24772
rect 27062 24760 27068 24772
rect 27120 24800 27126 24812
rect 27157 24803 27215 24809
rect 27157 24800 27169 24803
rect 27120 24772 27169 24800
rect 27120 24760 27126 24772
rect 27157 24769 27169 24772
rect 27203 24769 27215 24803
rect 27157 24763 27215 24769
rect 27706 24760 27712 24812
rect 27764 24800 27770 24812
rect 27801 24803 27859 24809
rect 27801 24800 27813 24803
rect 27764 24772 27813 24800
rect 27764 24760 27770 24772
rect 27801 24769 27813 24772
rect 27847 24769 27859 24803
rect 27801 24763 27859 24769
rect 20073 24735 20131 24741
rect 20073 24701 20085 24735
rect 20119 24732 20131 24735
rect 20162 24732 20168 24744
rect 20119 24704 20168 24732
rect 20119 24701 20131 24704
rect 20073 24695 20131 24701
rect 20162 24692 20168 24704
rect 20220 24692 20226 24744
rect 21174 24732 21180 24744
rect 21135 24704 21180 24732
rect 21174 24692 21180 24704
rect 21232 24692 21238 24744
rect 22649 24735 22707 24741
rect 22649 24701 22661 24735
rect 22695 24732 22707 24735
rect 22738 24732 22744 24744
rect 22695 24704 22744 24732
rect 22695 24701 22707 24704
rect 22649 24695 22707 24701
rect 22738 24692 22744 24704
rect 22796 24692 22802 24744
rect 24044 24732 24072 24760
rect 24581 24735 24639 24741
rect 24581 24732 24593 24735
rect 24044 24704 24593 24732
rect 24581 24701 24593 24704
rect 24627 24701 24639 24735
rect 24581 24695 24639 24701
rect 24670 24692 24676 24744
rect 24728 24732 24734 24744
rect 24765 24735 24823 24741
rect 24765 24732 24777 24735
rect 24728 24704 24777 24732
rect 24728 24692 24734 24704
rect 24765 24701 24777 24704
rect 24811 24701 24823 24735
rect 25774 24732 25780 24744
rect 25735 24704 25780 24732
rect 24765 24695 24823 24701
rect 25774 24692 25780 24704
rect 25832 24692 25838 24744
rect 18782 24664 18788 24676
rect 18743 24636 18788 24664
rect 18782 24624 18788 24636
rect 18840 24624 18846 24676
rect 24029 24667 24087 24673
rect 24029 24633 24041 24667
rect 24075 24664 24087 24667
rect 24118 24664 24124 24676
rect 24075 24636 24124 24664
rect 24075 24633 24087 24636
rect 24029 24627 24087 24633
rect 24118 24624 24124 24636
rect 24176 24624 24182 24676
rect 1765 24599 1823 24605
rect 1765 24565 1777 24599
rect 1811 24596 1823 24599
rect 15746 24596 15752 24608
rect 1811 24568 15752 24596
rect 1811 24565 1823 24568
rect 1765 24559 1823 24565
rect 15746 24556 15752 24568
rect 15804 24556 15810 24608
rect 19705 24599 19763 24605
rect 19705 24565 19717 24599
rect 19751 24596 19763 24599
rect 19886 24596 19892 24608
rect 19751 24568 19892 24596
rect 19751 24565 19763 24568
rect 19705 24559 19763 24565
rect 19886 24556 19892 24568
rect 19944 24556 19950 24608
rect 24670 24556 24676 24608
rect 24728 24596 24734 24608
rect 24728 24568 24773 24596
rect 24728 24556 24734 24568
rect 1104 24506 28888 24528
rect 1104 24454 4423 24506
rect 4475 24454 4487 24506
rect 4539 24454 4551 24506
rect 4603 24454 4615 24506
rect 4667 24454 4679 24506
rect 4731 24454 11369 24506
rect 11421 24454 11433 24506
rect 11485 24454 11497 24506
rect 11549 24454 11561 24506
rect 11613 24454 11625 24506
rect 11677 24454 18315 24506
rect 18367 24454 18379 24506
rect 18431 24454 18443 24506
rect 18495 24454 18507 24506
rect 18559 24454 18571 24506
rect 18623 24454 25261 24506
rect 25313 24454 25325 24506
rect 25377 24454 25389 24506
rect 25441 24454 25453 24506
rect 25505 24454 25517 24506
rect 25569 24454 28888 24506
rect 1104 24432 28888 24454
rect 17313 24395 17371 24401
rect 17313 24361 17325 24395
rect 17359 24392 17371 24395
rect 17494 24392 17500 24404
rect 17359 24364 17500 24392
rect 17359 24361 17371 24364
rect 17313 24355 17371 24361
rect 17494 24352 17500 24364
rect 17552 24352 17558 24404
rect 21634 24392 21640 24404
rect 21595 24364 21640 24392
rect 21634 24352 21640 24364
rect 21692 24352 21698 24404
rect 23661 24395 23719 24401
rect 23661 24361 23673 24395
rect 23707 24392 23719 24395
rect 23750 24392 23756 24404
rect 23707 24364 23756 24392
rect 23707 24361 23719 24364
rect 23661 24355 23719 24361
rect 23750 24352 23756 24364
rect 23808 24352 23814 24404
rect 24765 24395 24823 24401
rect 24765 24361 24777 24395
rect 24811 24392 24823 24395
rect 24946 24392 24952 24404
rect 24811 24364 24952 24392
rect 24811 24361 24823 24364
rect 24765 24355 24823 24361
rect 24946 24352 24952 24364
rect 25004 24352 25010 24404
rect 28350 24256 28356 24268
rect 28311 24228 28356 24256
rect 28350 24216 28356 24228
rect 28408 24216 28414 24268
rect 17126 24188 17132 24200
rect 17087 24160 17132 24188
rect 17126 24148 17132 24160
rect 17184 24148 17190 24200
rect 17310 24188 17316 24200
rect 17271 24160 17316 24188
rect 17310 24148 17316 24160
rect 17368 24148 17374 24200
rect 19426 24188 19432 24200
rect 19387 24160 19432 24188
rect 19426 24148 19432 24160
rect 19484 24148 19490 24200
rect 22370 24148 22376 24200
rect 22428 24188 22434 24200
rect 22750 24191 22808 24197
rect 22750 24188 22762 24191
rect 22428 24160 22762 24188
rect 22428 24148 22434 24160
rect 22750 24157 22762 24160
rect 22796 24157 22808 24191
rect 22750 24151 22808 24157
rect 23017 24191 23075 24197
rect 23017 24157 23029 24191
rect 23063 24188 23075 24191
rect 23382 24188 23388 24200
rect 23063 24160 23388 24188
rect 23063 24157 23075 24160
rect 23017 24151 23075 24157
rect 23382 24148 23388 24160
rect 23440 24148 23446 24200
rect 24670 24188 24676 24200
rect 24631 24160 24676 24188
rect 24670 24148 24676 24160
rect 24728 24148 24734 24200
rect 24854 24148 24860 24200
rect 24912 24188 24918 24200
rect 25682 24188 25688 24200
rect 24912 24160 25688 24188
rect 24912 24148 24918 24160
rect 25682 24148 25688 24160
rect 25740 24148 25746 24200
rect 26510 24188 26516 24200
rect 26471 24160 26516 24188
rect 26510 24148 26516 24160
rect 26568 24148 26574 24200
rect 19702 24129 19708 24132
rect 19696 24083 19708 24129
rect 19760 24120 19766 24132
rect 23474 24120 23480 24132
rect 19760 24092 19796 24120
rect 23435 24092 23480 24120
rect 19702 24080 19708 24083
rect 19760 24080 19766 24092
rect 23474 24080 23480 24092
rect 23532 24080 23538 24132
rect 23658 24080 23664 24132
rect 23716 24129 23722 24132
rect 23716 24123 23735 24129
rect 23723 24089 23735 24123
rect 23716 24083 23735 24089
rect 26697 24123 26755 24129
rect 26697 24089 26709 24123
rect 26743 24120 26755 24123
rect 27338 24120 27344 24132
rect 26743 24092 27344 24120
rect 26743 24089 26755 24092
rect 26697 24083 26755 24089
rect 23716 24080 23722 24083
rect 27338 24080 27344 24092
rect 27396 24080 27402 24132
rect 20809 24055 20867 24061
rect 20809 24021 20821 24055
rect 20855 24052 20867 24055
rect 20990 24052 20996 24064
rect 20855 24024 20996 24052
rect 20855 24021 20867 24024
rect 20809 24015 20867 24021
rect 20990 24012 20996 24024
rect 21048 24012 21054 24064
rect 23845 24055 23903 24061
rect 23845 24021 23857 24055
rect 23891 24052 23903 24055
rect 24026 24052 24032 24064
rect 23891 24024 24032 24052
rect 23891 24021 23903 24024
rect 23845 24015 23903 24021
rect 24026 24012 24032 24024
rect 24084 24012 24090 24064
rect 1104 23962 29048 23984
rect 1104 23910 7896 23962
rect 7948 23910 7960 23962
rect 8012 23910 8024 23962
rect 8076 23910 8088 23962
rect 8140 23910 8152 23962
rect 8204 23910 14842 23962
rect 14894 23910 14906 23962
rect 14958 23910 14970 23962
rect 15022 23910 15034 23962
rect 15086 23910 15098 23962
rect 15150 23910 21788 23962
rect 21840 23910 21852 23962
rect 21904 23910 21916 23962
rect 21968 23910 21980 23962
rect 22032 23910 22044 23962
rect 22096 23910 28734 23962
rect 28786 23910 28798 23962
rect 28850 23910 28862 23962
rect 28914 23910 28926 23962
rect 28978 23910 28990 23962
rect 29042 23910 29048 23962
rect 1104 23888 29048 23910
rect 19702 23848 19708 23860
rect 19663 23820 19708 23848
rect 19702 23808 19708 23820
rect 19760 23808 19766 23860
rect 20438 23848 20444 23860
rect 20399 23820 20444 23848
rect 20438 23808 20444 23820
rect 20496 23808 20502 23860
rect 20898 23848 20904 23860
rect 20859 23820 20904 23848
rect 20898 23808 20904 23820
rect 20956 23808 20962 23860
rect 27338 23848 27344 23860
rect 27299 23820 27344 23848
rect 27338 23808 27344 23820
rect 27396 23808 27402 23860
rect 16574 23740 16580 23792
rect 16632 23780 16638 23792
rect 17465 23783 17523 23789
rect 17465 23780 17477 23783
rect 16632 23752 17477 23780
rect 16632 23740 16638 23752
rect 17465 23749 17477 23752
rect 17511 23749 17523 23783
rect 17465 23743 17523 23749
rect 17681 23783 17739 23789
rect 17681 23749 17693 23783
rect 17727 23749 17739 23783
rect 19794 23780 19800 23792
rect 17681 23743 17739 23749
rect 18800 23752 19800 23780
rect 17696 23712 17724 23743
rect 18325 23715 18383 23721
rect 18325 23712 18337 23715
rect 17696 23684 18337 23712
rect 18325 23681 18337 23684
rect 18371 23712 18383 23715
rect 18690 23712 18696 23724
rect 18371 23684 18696 23712
rect 18371 23681 18383 23684
rect 18325 23675 18383 23681
rect 18690 23672 18696 23684
rect 18748 23672 18754 23724
rect 18800 23721 18828 23752
rect 19794 23740 19800 23752
rect 19852 23780 19858 23792
rect 20254 23780 20260 23792
rect 19852 23752 20260 23780
rect 19852 23740 19858 23752
rect 20254 23740 20260 23752
rect 20312 23740 20318 23792
rect 20809 23783 20867 23789
rect 20809 23749 20821 23783
rect 20855 23780 20867 23783
rect 20990 23780 20996 23792
rect 20855 23752 20996 23780
rect 20855 23749 20867 23752
rect 20809 23743 20867 23749
rect 20990 23740 20996 23752
rect 21048 23740 21054 23792
rect 26510 23740 26516 23792
rect 26568 23780 26574 23792
rect 26568 23752 27936 23780
rect 26568 23740 26574 23752
rect 18785 23715 18843 23721
rect 18785 23681 18797 23715
rect 18831 23681 18843 23715
rect 18785 23675 18843 23681
rect 18969 23715 19027 23721
rect 18969 23681 18981 23715
rect 19015 23681 19027 23715
rect 19886 23712 19892 23724
rect 19847 23684 19892 23712
rect 18969 23675 19027 23681
rect 18984 23644 19012 23675
rect 19886 23672 19892 23684
rect 19944 23672 19950 23724
rect 26878 23672 26884 23724
rect 26936 23712 26942 23724
rect 27433 23715 27491 23721
rect 27433 23712 27445 23715
rect 26936 23684 27445 23712
rect 26936 23672 26942 23684
rect 27433 23681 27445 23684
rect 27479 23712 27491 23715
rect 27614 23712 27620 23724
rect 27479 23684 27620 23712
rect 27479 23681 27491 23684
rect 27433 23675 27491 23681
rect 27614 23672 27620 23684
rect 27672 23672 27678 23724
rect 27908 23721 27936 23752
rect 27893 23715 27951 23721
rect 27893 23681 27905 23715
rect 27939 23681 27951 23715
rect 27893 23675 27951 23681
rect 17604 23616 19012 23644
rect 21085 23647 21143 23653
rect 17604 23588 17632 23616
rect 21085 23613 21097 23647
rect 21131 23644 21143 23647
rect 21174 23644 21180 23656
rect 21131 23616 21180 23644
rect 21131 23613 21143 23616
rect 21085 23607 21143 23613
rect 21174 23604 21180 23616
rect 21232 23644 21238 23656
rect 21634 23644 21640 23656
rect 21232 23616 21640 23644
rect 21232 23604 21238 23616
rect 21634 23604 21640 23616
rect 21692 23604 21698 23656
rect 17313 23579 17371 23585
rect 17313 23545 17325 23579
rect 17359 23576 17371 23579
rect 17586 23576 17592 23588
rect 17359 23548 17592 23576
rect 17359 23545 17371 23548
rect 17313 23539 17371 23545
rect 17586 23536 17592 23548
rect 17644 23536 17650 23588
rect 16390 23468 16396 23520
rect 16448 23508 16454 23520
rect 17497 23511 17555 23517
rect 17497 23508 17509 23511
rect 16448 23480 17509 23508
rect 16448 23468 16454 23480
rect 17497 23477 17509 23480
rect 17543 23477 17555 23511
rect 17497 23471 17555 23477
rect 17678 23468 17684 23520
rect 17736 23508 17742 23520
rect 18233 23511 18291 23517
rect 18233 23508 18245 23511
rect 17736 23480 18245 23508
rect 17736 23468 17742 23480
rect 18233 23477 18245 23480
rect 18279 23477 18291 23511
rect 18233 23471 18291 23477
rect 18874 23468 18880 23520
rect 18932 23508 18938 23520
rect 18969 23511 19027 23517
rect 18969 23508 18981 23511
rect 18932 23480 18981 23508
rect 18932 23468 18938 23480
rect 18969 23477 18981 23480
rect 19015 23477 19027 23511
rect 18969 23471 19027 23477
rect 26510 23468 26516 23520
rect 26568 23508 26574 23520
rect 26605 23511 26663 23517
rect 26605 23508 26617 23511
rect 26568 23480 26617 23508
rect 26568 23468 26574 23480
rect 26605 23477 26617 23480
rect 26651 23477 26663 23511
rect 26605 23471 26663 23477
rect 1104 23418 28888 23440
rect 1104 23366 4423 23418
rect 4475 23366 4487 23418
rect 4539 23366 4551 23418
rect 4603 23366 4615 23418
rect 4667 23366 4679 23418
rect 4731 23366 11369 23418
rect 11421 23366 11433 23418
rect 11485 23366 11497 23418
rect 11549 23366 11561 23418
rect 11613 23366 11625 23418
rect 11677 23366 18315 23418
rect 18367 23366 18379 23418
rect 18431 23366 18443 23418
rect 18495 23366 18507 23418
rect 18559 23366 18571 23418
rect 18623 23366 25261 23418
rect 25313 23366 25325 23418
rect 25377 23366 25389 23418
rect 25441 23366 25453 23418
rect 25505 23366 25517 23418
rect 25569 23366 28888 23418
rect 1104 23344 28888 23366
rect 17221 23307 17279 23313
rect 17221 23273 17233 23307
rect 17267 23304 17279 23307
rect 17310 23304 17316 23316
rect 17267 23276 17316 23304
rect 17267 23273 17279 23276
rect 17221 23267 17279 23273
rect 17310 23264 17316 23276
rect 17368 23264 17374 23316
rect 17497 23239 17555 23245
rect 17497 23205 17509 23239
rect 17543 23236 17555 23239
rect 18325 23239 18383 23245
rect 18325 23236 18337 23239
rect 17543 23208 18337 23236
rect 17543 23205 17555 23208
rect 17497 23199 17555 23205
rect 18325 23205 18337 23208
rect 18371 23205 18383 23239
rect 18325 23199 18383 23205
rect 23566 23196 23572 23248
rect 23624 23236 23630 23248
rect 23753 23239 23811 23245
rect 23753 23236 23765 23239
rect 23624 23208 23765 23236
rect 23624 23196 23630 23208
rect 23753 23205 23765 23208
rect 23799 23205 23811 23239
rect 23753 23199 23811 23205
rect 15856 23140 16528 23168
rect 15856 23109 15884 23140
rect 15657 23103 15715 23109
rect 15657 23069 15669 23103
rect 15703 23069 15715 23103
rect 15657 23063 15715 23069
rect 15841 23103 15899 23109
rect 15841 23069 15853 23103
rect 15887 23069 15899 23103
rect 16390 23100 16396 23112
rect 16351 23072 16396 23100
rect 15841 23063 15899 23069
rect 15672 23032 15700 23063
rect 16390 23060 16396 23072
rect 16448 23060 16454 23112
rect 16500 23109 16528 23140
rect 17218 23128 17224 23180
rect 17276 23128 17282 23180
rect 17678 23168 17684 23180
rect 17639 23140 17684 23168
rect 17678 23128 17684 23140
rect 17736 23128 17742 23180
rect 19794 23168 19800 23180
rect 17788 23140 19656 23168
rect 19755 23140 19800 23168
rect 16485 23103 16543 23109
rect 16485 23069 16497 23103
rect 16531 23100 16543 23103
rect 16574 23100 16580 23112
rect 16531 23072 16580 23100
rect 16531 23069 16543 23072
rect 16485 23063 16543 23069
rect 16574 23060 16580 23072
rect 16632 23060 16638 23112
rect 17034 23060 17040 23112
rect 17092 23100 17098 23112
rect 17236 23100 17264 23128
rect 17405 23103 17463 23109
rect 17405 23100 17417 23103
rect 17092 23072 17417 23100
rect 17092 23060 17098 23072
rect 17405 23069 17417 23072
rect 17451 23069 17463 23103
rect 17586 23100 17592 23112
rect 17547 23072 17592 23100
rect 17405 23063 17463 23069
rect 17586 23060 17592 23072
rect 17644 23100 17650 23112
rect 17788 23100 17816 23140
rect 17644 23072 17816 23100
rect 17644 23060 17650 23072
rect 17862 23060 17868 23112
rect 17920 23100 17926 23112
rect 18325 23103 18383 23109
rect 17920 23072 17965 23100
rect 17920 23060 17926 23072
rect 18325 23069 18337 23103
rect 18371 23069 18383 23103
rect 18325 23063 18383 23069
rect 18509 23103 18567 23109
rect 18509 23069 18521 23103
rect 18555 23100 18567 23103
rect 18690 23100 18696 23112
rect 18555 23072 18696 23100
rect 18555 23069 18567 23072
rect 18509 23063 18567 23069
rect 16206 23032 16212 23044
rect 15672 23004 16212 23032
rect 16206 22992 16212 23004
rect 16264 23032 16270 23044
rect 16408 23032 16436 23060
rect 16264 23004 16436 23032
rect 16669 23035 16727 23041
rect 16264 22992 16270 23004
rect 16669 23001 16681 23035
rect 16715 23032 16727 23035
rect 17218 23032 17224 23044
rect 16715 23004 17224 23032
rect 16715 23001 16727 23004
rect 16669 22995 16727 23001
rect 17218 22992 17224 23004
rect 17276 23032 17282 23044
rect 18340 23032 18368 23063
rect 18690 23060 18696 23072
rect 18748 23060 18754 23112
rect 19628 23109 19656 23140
rect 19794 23128 19800 23140
rect 19852 23128 19858 23180
rect 20162 23128 20168 23180
rect 20220 23168 20226 23180
rect 20530 23168 20536 23180
rect 20220 23140 20536 23168
rect 20220 23128 20226 23140
rect 20530 23128 20536 23140
rect 20588 23128 20594 23180
rect 25038 23168 25044 23180
rect 23676 23140 25044 23168
rect 23676 23112 23704 23140
rect 25038 23128 25044 23140
rect 25096 23168 25102 23180
rect 25225 23171 25283 23177
rect 25225 23168 25237 23171
rect 25096 23140 25237 23168
rect 25096 23128 25102 23140
rect 25225 23137 25237 23140
rect 25271 23168 25283 23171
rect 25774 23168 25780 23180
rect 25271 23140 25780 23168
rect 25271 23137 25283 23140
rect 25225 23131 25283 23137
rect 25774 23128 25780 23140
rect 25832 23128 25838 23180
rect 26510 23168 26516 23180
rect 26471 23140 26516 23168
rect 26510 23128 26516 23140
rect 26568 23128 26574 23180
rect 28353 23171 28411 23177
rect 28353 23137 28365 23171
rect 28399 23168 28411 23171
rect 29914 23168 29920 23180
rect 28399 23140 29920 23168
rect 28399 23137 28411 23140
rect 28353 23131 28411 23137
rect 29914 23128 29920 23140
rect 29972 23128 29978 23180
rect 19613 23103 19671 23109
rect 19613 23069 19625 23103
rect 19659 23069 19671 23103
rect 20714 23100 20720 23112
rect 20675 23072 20720 23100
rect 19613 23063 19671 23069
rect 20714 23060 20720 23072
rect 20772 23060 20778 23112
rect 23477 23103 23535 23109
rect 23477 23069 23489 23103
rect 23523 23100 23535 23103
rect 23658 23100 23664 23112
rect 23523 23072 23664 23100
rect 23523 23069 23535 23072
rect 23477 23063 23535 23069
rect 23658 23060 23664 23072
rect 23716 23060 23722 23112
rect 24670 23060 24676 23112
rect 24728 23100 24734 23112
rect 25133 23103 25191 23109
rect 25133 23100 25145 23103
rect 24728 23072 25145 23100
rect 24728 23060 24734 23072
rect 25133 23069 25145 23072
rect 25179 23069 25191 23103
rect 25133 23063 25191 23069
rect 23750 23032 23756 23044
rect 17276 23004 18368 23032
rect 23663 23004 23756 23032
rect 17276 22992 17282 23004
rect 23750 22992 23756 23004
rect 23808 23032 23814 23044
rect 26142 23032 26148 23044
rect 23808 23004 26148 23032
rect 23808 22992 23814 23004
rect 26142 22992 26148 23004
rect 26200 22992 26206 23044
rect 26697 23035 26755 23041
rect 26697 23001 26709 23035
rect 26743 23032 26755 23035
rect 27246 23032 27252 23044
rect 26743 23004 27252 23032
rect 26743 23001 26755 23004
rect 26697 22995 26755 23001
rect 27246 22992 27252 23004
rect 27304 22992 27310 23044
rect 15746 22964 15752 22976
rect 15707 22936 15752 22964
rect 15746 22924 15752 22936
rect 15804 22924 15810 22976
rect 19429 22967 19487 22973
rect 19429 22933 19441 22967
rect 19475 22964 19487 22967
rect 19978 22964 19984 22976
rect 19475 22936 19984 22964
rect 19475 22933 19487 22936
rect 19429 22927 19487 22933
rect 19978 22924 19984 22936
rect 20036 22924 20042 22976
rect 20898 22964 20904 22976
rect 20859 22936 20904 22964
rect 20898 22924 20904 22936
rect 20956 22924 20962 22976
rect 23474 22924 23480 22976
rect 23532 22964 23538 22976
rect 23569 22967 23627 22973
rect 23569 22964 23581 22967
rect 23532 22936 23581 22964
rect 23532 22924 23538 22936
rect 23569 22933 23581 22936
rect 23615 22964 23627 22967
rect 24670 22964 24676 22976
rect 23615 22936 24676 22964
rect 23615 22933 23627 22936
rect 23569 22927 23627 22933
rect 24670 22924 24676 22936
rect 24728 22924 24734 22976
rect 25501 22967 25559 22973
rect 25501 22933 25513 22967
rect 25547 22964 25559 22967
rect 25590 22964 25596 22976
rect 25547 22936 25596 22964
rect 25547 22933 25559 22936
rect 25501 22927 25559 22933
rect 25590 22924 25596 22936
rect 25648 22924 25654 22976
rect 1104 22874 29048 22896
rect 1104 22822 7896 22874
rect 7948 22822 7960 22874
rect 8012 22822 8024 22874
rect 8076 22822 8088 22874
rect 8140 22822 8152 22874
rect 8204 22822 14842 22874
rect 14894 22822 14906 22874
rect 14958 22822 14970 22874
rect 15022 22822 15034 22874
rect 15086 22822 15098 22874
rect 15150 22822 21788 22874
rect 21840 22822 21852 22874
rect 21904 22822 21916 22874
rect 21968 22822 21980 22874
rect 22032 22822 22044 22874
rect 22096 22822 28734 22874
rect 28786 22822 28798 22874
rect 28850 22822 28862 22874
rect 28914 22822 28926 22874
rect 28978 22822 28990 22874
rect 29042 22822 29048 22874
rect 1104 22800 29048 22822
rect 17034 22720 17040 22772
rect 17092 22760 17098 22772
rect 17092 22732 17908 22760
rect 17092 22720 17098 22732
rect 15746 22652 15752 22704
rect 15804 22692 15810 22704
rect 15804 22664 17172 22692
rect 15804 22652 15810 22664
rect 17034 22624 17040 22636
rect 16995 22596 17040 22624
rect 17034 22584 17040 22596
rect 17092 22584 17098 22636
rect 17144 22633 17172 22664
rect 17129 22627 17187 22633
rect 17129 22593 17141 22627
rect 17175 22593 17187 22627
rect 17129 22587 17187 22593
rect 17218 22584 17224 22636
rect 17276 22624 17282 22636
rect 17497 22627 17555 22633
rect 17276 22596 17321 22624
rect 17276 22584 17282 22596
rect 17497 22593 17509 22627
rect 17543 22624 17555 22627
rect 17770 22624 17776 22636
rect 17543 22596 17776 22624
rect 17543 22593 17555 22596
rect 17497 22587 17555 22593
rect 17770 22584 17776 22596
rect 17828 22584 17834 22636
rect 17880 22624 17908 22732
rect 18230 22720 18236 22772
rect 18288 22760 18294 22772
rect 18509 22763 18567 22769
rect 18509 22760 18521 22763
rect 18288 22732 18521 22760
rect 18288 22720 18294 22732
rect 18509 22729 18521 22732
rect 18555 22729 18567 22763
rect 20714 22760 20720 22772
rect 20675 22732 20720 22760
rect 18509 22723 18567 22729
rect 20714 22720 20720 22732
rect 20772 22720 20778 22772
rect 21174 22760 21180 22772
rect 21135 22732 21180 22760
rect 21174 22720 21180 22732
rect 21232 22720 21238 22772
rect 26142 22720 26148 22772
rect 26200 22760 26206 22772
rect 26513 22763 26571 22769
rect 26513 22760 26525 22763
rect 26200 22732 26525 22760
rect 26200 22720 26206 22732
rect 26513 22729 26525 22732
rect 26559 22729 26571 22763
rect 27246 22760 27252 22772
rect 27207 22732 27252 22760
rect 26513 22723 26571 22729
rect 27246 22720 27252 22732
rect 27304 22720 27310 22772
rect 21085 22695 21143 22701
rect 21085 22661 21097 22695
rect 21131 22692 21143 22695
rect 21266 22692 21272 22704
rect 21131 22664 21272 22692
rect 21131 22661 21143 22664
rect 21085 22655 21143 22661
rect 21266 22652 21272 22664
rect 21324 22652 21330 22704
rect 23382 22652 23388 22704
rect 23440 22692 23446 22704
rect 23440 22664 25176 22692
rect 23440 22652 23446 22664
rect 18690 22624 18696 22636
rect 17880 22596 18696 22624
rect 18690 22584 18696 22596
rect 18748 22584 18754 22636
rect 18874 22624 18880 22636
rect 18835 22596 18880 22624
rect 18874 22584 18880 22596
rect 18932 22584 18938 22636
rect 18966 22584 18972 22636
rect 19024 22624 19030 22636
rect 19153 22627 19211 22633
rect 19024 22596 19068 22624
rect 19024 22584 19030 22596
rect 19153 22593 19165 22627
rect 19199 22593 19211 22627
rect 19794 22624 19800 22636
rect 19755 22596 19800 22624
rect 19153 22587 19211 22593
rect 17310 22516 17316 22568
rect 17368 22556 17374 22568
rect 17788 22556 17816 22584
rect 19168 22556 19196 22587
rect 19794 22584 19800 22596
rect 19852 22584 19858 22636
rect 22646 22584 22652 22636
rect 22704 22624 22710 22636
rect 22741 22627 22799 22633
rect 22741 22624 22753 22627
rect 22704 22596 22753 22624
rect 22704 22584 22710 22596
rect 22741 22593 22753 22596
rect 22787 22593 22799 22627
rect 22741 22587 22799 22593
rect 22925 22627 22983 22633
rect 22925 22593 22937 22627
rect 22971 22624 22983 22627
rect 23750 22624 23756 22636
rect 22971 22596 23756 22624
rect 22971 22593 22983 22596
rect 22925 22587 22983 22593
rect 23750 22584 23756 22596
rect 23808 22584 23814 22636
rect 23845 22627 23903 22633
rect 23845 22593 23857 22627
rect 23891 22624 23903 22627
rect 23934 22624 23940 22636
rect 23891 22596 23940 22624
rect 23891 22593 23903 22596
rect 23845 22587 23903 22593
rect 23934 22584 23940 22596
rect 23992 22584 23998 22636
rect 24026 22584 24032 22636
rect 24084 22624 24090 22636
rect 24302 22624 24308 22636
rect 24084 22596 24129 22624
rect 24263 22596 24308 22624
rect 24084 22584 24090 22596
rect 24302 22584 24308 22596
rect 24360 22584 24366 22636
rect 25148 22633 25176 22664
rect 25133 22627 25191 22633
rect 25133 22593 25145 22627
rect 25179 22593 25191 22627
rect 25133 22587 25191 22593
rect 25222 22584 25228 22636
rect 25280 22624 25286 22636
rect 25389 22627 25447 22633
rect 25389 22624 25401 22627
rect 25280 22596 25401 22624
rect 25280 22584 25286 22596
rect 25389 22593 25401 22596
rect 25435 22593 25447 22627
rect 25389 22587 25447 22593
rect 27341 22627 27399 22633
rect 27341 22593 27353 22627
rect 27387 22624 27399 22627
rect 28626 22624 28632 22636
rect 27387 22596 28632 22624
rect 27387 22593 27399 22596
rect 27341 22587 27399 22593
rect 28626 22584 28632 22596
rect 28684 22584 28690 22636
rect 17368 22528 17413 22556
rect 17788 22528 19196 22556
rect 21361 22559 21419 22565
rect 17368 22516 17374 22528
rect 21361 22525 21373 22559
rect 21407 22556 21419 22559
rect 21634 22556 21640 22568
rect 21407 22528 21640 22556
rect 21407 22525 21419 22528
rect 21361 22519 21419 22525
rect 21634 22516 21640 22528
rect 21692 22516 21698 22568
rect 24118 22556 24124 22568
rect 24079 22528 24124 22556
rect 24118 22516 24124 22528
rect 24176 22516 24182 22568
rect 18785 22491 18843 22497
rect 18785 22457 18797 22491
rect 18831 22488 18843 22491
rect 19978 22488 19984 22500
rect 18831 22460 19984 22488
rect 18831 22457 18843 22460
rect 18785 22451 18843 22457
rect 19978 22448 19984 22460
rect 20036 22448 20042 22500
rect 23566 22448 23572 22500
rect 23624 22488 23630 22500
rect 23937 22491 23995 22497
rect 23937 22488 23949 22491
rect 23624 22460 23949 22488
rect 23624 22448 23630 22460
rect 23937 22457 23949 22460
rect 23983 22457 23995 22491
rect 23937 22451 23995 22457
rect 16850 22420 16856 22432
rect 16811 22392 16856 22420
rect 16850 22380 16856 22392
rect 16908 22380 16914 22432
rect 19058 22380 19064 22432
rect 19116 22420 19122 22432
rect 19705 22423 19763 22429
rect 19705 22420 19717 22423
rect 19116 22392 19717 22420
rect 19116 22380 19122 22392
rect 19705 22389 19717 22392
rect 19751 22389 19763 22423
rect 19705 22383 19763 22389
rect 22462 22380 22468 22432
rect 22520 22420 22526 22432
rect 22833 22423 22891 22429
rect 22833 22420 22845 22423
rect 22520 22392 22845 22420
rect 22520 22380 22526 22392
rect 22833 22389 22845 22392
rect 22879 22389 22891 22423
rect 22833 22383 22891 22389
rect 23661 22423 23719 22429
rect 23661 22389 23673 22423
rect 23707 22420 23719 22423
rect 23842 22420 23848 22432
rect 23707 22392 23848 22420
rect 23707 22389 23719 22392
rect 23661 22383 23719 22389
rect 23842 22380 23848 22392
rect 23900 22380 23906 22432
rect 28074 22420 28080 22432
rect 28035 22392 28080 22420
rect 28074 22380 28080 22392
rect 28132 22380 28138 22432
rect 1104 22330 28888 22352
rect 1104 22278 4423 22330
rect 4475 22278 4487 22330
rect 4539 22278 4551 22330
rect 4603 22278 4615 22330
rect 4667 22278 4679 22330
rect 4731 22278 11369 22330
rect 11421 22278 11433 22330
rect 11485 22278 11497 22330
rect 11549 22278 11561 22330
rect 11613 22278 11625 22330
rect 11677 22278 18315 22330
rect 18367 22278 18379 22330
rect 18431 22278 18443 22330
rect 18495 22278 18507 22330
rect 18559 22278 18571 22330
rect 18623 22278 25261 22330
rect 25313 22278 25325 22330
rect 25377 22278 25389 22330
rect 25441 22278 25453 22330
rect 25505 22278 25517 22330
rect 25569 22278 28888 22330
rect 1104 22256 28888 22278
rect 18690 22176 18696 22228
rect 18748 22216 18754 22228
rect 19613 22219 19671 22225
rect 19613 22216 19625 22219
rect 18748 22188 19625 22216
rect 18748 22176 18754 22188
rect 19613 22185 19625 22188
rect 19659 22185 19671 22219
rect 19613 22179 19671 22185
rect 23934 22176 23940 22228
rect 23992 22216 23998 22228
rect 24394 22216 24400 22228
rect 23992 22188 24400 22216
rect 23992 22176 23998 22188
rect 24394 22176 24400 22188
rect 24452 22176 24458 22228
rect 25130 22176 25136 22228
rect 25188 22216 25194 22228
rect 25225 22219 25283 22225
rect 25225 22216 25237 22219
rect 25188 22188 25237 22216
rect 25188 22176 25194 22188
rect 25225 22185 25237 22188
rect 25271 22185 25283 22219
rect 25225 22179 25283 22185
rect 17126 22080 17132 22092
rect 16040 22052 17132 22080
rect 16040 22021 16068 22052
rect 17126 22040 17132 22052
rect 17184 22040 17190 22092
rect 23937 22083 23995 22089
rect 23937 22049 23949 22083
rect 23983 22080 23995 22083
rect 27522 22080 27528 22092
rect 23983 22052 24808 22080
rect 27483 22052 27528 22080
rect 23983 22049 23995 22052
rect 23937 22043 23995 22049
rect 16025 22015 16083 22021
rect 16025 21981 16037 22015
rect 16071 21981 16083 22015
rect 16025 21975 16083 21981
rect 16209 22015 16267 22021
rect 16209 21981 16221 22015
rect 16255 22012 16267 22015
rect 16850 22012 16856 22024
rect 16255 21984 16856 22012
rect 16255 21981 16267 21984
rect 16209 21975 16267 21981
rect 16850 21972 16856 21984
rect 16908 21972 16914 22024
rect 18230 21972 18236 22024
rect 18288 22012 18294 22024
rect 19426 22012 19432 22024
rect 18288 21984 19432 22012
rect 18288 21972 18294 21984
rect 19426 21972 19432 21984
rect 19484 22012 19490 22024
rect 20441 22015 20499 22021
rect 20441 22012 20453 22015
rect 19484 21984 20453 22012
rect 19484 21972 19490 21984
rect 20441 21981 20453 21984
rect 20487 21981 20499 22015
rect 20441 21975 20499 21981
rect 21450 21972 21456 22024
rect 21508 22012 21514 22024
rect 22281 22015 22339 22021
rect 22281 22012 22293 22015
rect 21508 21984 22293 22012
rect 21508 21972 21514 21984
rect 22281 21981 22293 21984
rect 22327 21981 22339 22015
rect 22462 22012 22468 22024
rect 22423 21984 22468 22012
rect 22281 21975 22339 21981
rect 22462 21972 22468 21984
rect 22520 21972 22526 22024
rect 22557 22015 22615 22021
rect 22557 21981 22569 22015
rect 22603 22012 22615 22015
rect 22922 22012 22928 22024
rect 22603 21984 22928 22012
rect 22603 21981 22615 21984
rect 22557 21975 22615 21981
rect 22922 21972 22928 21984
rect 22980 21972 22986 22024
rect 23842 22012 23848 22024
rect 23803 21984 23848 22012
rect 23842 21972 23848 21984
rect 23900 21972 23906 22024
rect 24029 22015 24087 22021
rect 24029 21981 24041 22015
rect 24075 21981 24087 22015
rect 24029 21975 24087 21981
rect 19521 21947 19579 21953
rect 19521 21913 19533 21947
rect 19567 21944 19579 21947
rect 19702 21944 19708 21956
rect 19567 21916 19708 21944
rect 19567 21913 19579 21916
rect 19521 21907 19579 21913
rect 19702 21904 19708 21916
rect 19760 21904 19766 21956
rect 20714 21953 20720 21956
rect 20708 21907 20720 21953
rect 20772 21944 20778 21956
rect 20772 21916 20808 21944
rect 20714 21904 20720 21907
rect 20772 21904 20778 21916
rect 16114 21876 16120 21888
rect 16075 21848 16120 21876
rect 16114 21836 16120 21848
rect 16172 21836 16178 21888
rect 21266 21836 21272 21888
rect 21324 21876 21330 21888
rect 21821 21879 21879 21885
rect 21821 21876 21833 21879
rect 21324 21848 21833 21876
rect 21324 21836 21330 21848
rect 21821 21845 21833 21848
rect 21867 21845 21879 21879
rect 21821 21839 21879 21845
rect 22379 21879 22437 21885
rect 22379 21845 22391 21879
rect 22425 21876 22437 21879
rect 23106 21876 23112 21888
rect 22425 21848 23112 21876
rect 22425 21845 22437 21848
rect 22379 21839 22437 21845
rect 23106 21836 23112 21848
rect 23164 21836 23170 21888
rect 24044 21876 24072 21975
rect 24210 21972 24216 22024
rect 24268 22012 24274 22024
rect 24581 22015 24639 22021
rect 24581 22012 24593 22015
rect 24268 21984 24593 22012
rect 24268 21972 24274 21984
rect 24581 21981 24593 21984
rect 24627 22012 24639 22015
rect 24670 22012 24676 22024
rect 24627 21984 24676 22012
rect 24627 21981 24639 21984
rect 24581 21975 24639 21981
rect 24670 21972 24676 21984
rect 24728 21972 24734 22024
rect 24780 22021 24808 22052
rect 27522 22040 27528 22052
rect 27580 22040 27586 22092
rect 28074 22040 28080 22092
rect 28132 22080 28138 22092
rect 28353 22083 28411 22089
rect 28353 22080 28365 22083
rect 28132 22052 28365 22080
rect 28132 22040 28138 22052
rect 28353 22049 28365 22052
rect 28399 22049 28411 22083
rect 28353 22043 28411 22049
rect 24765 22015 24823 22021
rect 24765 21981 24777 22015
rect 24811 21981 24823 22015
rect 24765 21975 24823 21981
rect 24857 22015 24915 22021
rect 24857 21981 24869 22015
rect 24903 21981 24915 22015
rect 24857 21975 24915 21981
rect 24949 22015 25007 22021
rect 24949 21981 24961 22015
rect 24995 22012 25007 22015
rect 26142 22012 26148 22024
rect 24995 21984 26148 22012
rect 24995 21981 25007 21984
rect 24949 21975 25007 21981
rect 24872 21888 24900 21975
rect 26142 21972 26148 21984
rect 26200 21972 26206 22024
rect 27890 21904 27896 21956
rect 27948 21944 27954 21956
rect 28169 21947 28227 21953
rect 28169 21944 28181 21947
rect 27948 21916 28181 21944
rect 27948 21904 27954 21916
rect 28169 21913 28181 21916
rect 28215 21913 28227 21947
rect 28169 21907 28227 21913
rect 24854 21876 24860 21888
rect 24044 21848 24860 21876
rect 24854 21836 24860 21848
rect 24912 21836 24918 21888
rect 1104 21786 29048 21808
rect 1104 21734 7896 21786
rect 7948 21734 7960 21786
rect 8012 21734 8024 21786
rect 8076 21734 8088 21786
rect 8140 21734 8152 21786
rect 8204 21734 14842 21786
rect 14894 21734 14906 21786
rect 14958 21734 14970 21786
rect 15022 21734 15034 21786
rect 15086 21734 15098 21786
rect 15150 21734 21788 21786
rect 21840 21734 21852 21786
rect 21904 21734 21916 21786
rect 21968 21734 21980 21786
rect 22032 21734 22044 21786
rect 22096 21734 28734 21786
rect 28786 21734 28798 21786
rect 28850 21734 28862 21786
rect 28914 21734 28926 21786
rect 28978 21734 28990 21786
rect 29042 21734 29048 21786
rect 1104 21712 29048 21734
rect 16206 21632 16212 21684
rect 16264 21672 16270 21684
rect 18233 21675 18291 21681
rect 18233 21672 18245 21675
rect 16264 21644 18245 21672
rect 16264 21632 16270 21644
rect 18233 21641 18245 21644
rect 18279 21641 18291 21675
rect 20714 21672 20720 21684
rect 20675 21644 20720 21672
rect 18233 21635 18291 21641
rect 20714 21632 20720 21644
rect 20772 21632 20778 21684
rect 22922 21672 22928 21684
rect 22883 21644 22928 21672
rect 22922 21632 22928 21644
rect 22980 21632 22986 21684
rect 27890 21672 27896 21684
rect 27851 21644 27896 21672
rect 27890 21632 27896 21644
rect 27948 21632 27954 21684
rect 16114 21564 16120 21616
rect 16172 21604 16178 21616
rect 17098 21607 17156 21613
rect 17098 21604 17110 21607
rect 16172 21576 17110 21604
rect 16172 21564 16178 21576
rect 17098 21573 17110 21576
rect 17144 21573 17156 21607
rect 17098 21567 17156 21573
rect 24394 21564 24400 21616
rect 24452 21604 24458 21616
rect 25590 21604 25596 21616
rect 24452 21576 25176 21604
rect 24452 21564 24458 21576
rect 19521 21539 19579 21545
rect 19521 21505 19533 21539
rect 19567 21536 19579 21539
rect 19702 21536 19708 21548
rect 19567 21508 19708 21536
rect 19567 21505 19579 21508
rect 19521 21499 19579 21505
rect 19702 21496 19708 21508
rect 19760 21496 19766 21548
rect 20898 21536 20904 21548
rect 20859 21508 20904 21536
rect 20898 21496 20904 21508
rect 20956 21496 20962 21548
rect 22370 21496 22376 21548
rect 22428 21536 22434 21548
rect 22649 21539 22707 21545
rect 22649 21536 22661 21539
rect 22428 21508 22661 21536
rect 22428 21496 22434 21508
rect 22649 21505 22661 21508
rect 22695 21505 22707 21539
rect 22649 21499 22707 21505
rect 23658 21496 23664 21548
rect 23716 21536 23722 21548
rect 23845 21539 23903 21545
rect 23845 21536 23857 21539
rect 23716 21508 23857 21536
rect 23716 21496 23722 21508
rect 23845 21505 23857 21508
rect 23891 21505 23903 21539
rect 23845 21499 23903 21505
rect 24118 21496 24124 21548
rect 24176 21536 24182 21548
rect 24176 21508 24440 21536
rect 24176 21496 24182 21508
rect 16853 21471 16911 21477
rect 16853 21437 16865 21471
rect 16899 21437 16911 21471
rect 16853 21431 16911 21437
rect 16868 21332 16896 21431
rect 22002 21428 22008 21480
rect 22060 21468 22066 21480
rect 22281 21471 22339 21477
rect 22281 21468 22293 21471
rect 22060 21440 22293 21468
rect 22060 21428 22066 21440
rect 22281 21437 22293 21440
rect 22327 21437 22339 21471
rect 22738 21468 22744 21480
rect 22651 21440 22744 21468
rect 22281 21431 22339 21437
rect 22738 21428 22744 21440
rect 22796 21468 22802 21480
rect 23937 21471 23995 21477
rect 22796 21440 23152 21468
rect 22796 21428 22802 21440
rect 19797 21403 19855 21409
rect 19797 21369 19809 21403
rect 19843 21400 19855 21403
rect 22756 21400 22784 21428
rect 19843 21372 22784 21400
rect 19843 21369 19855 21372
rect 19797 21363 19855 21369
rect 18230 21332 18236 21344
rect 16868 21304 18236 21332
rect 18230 21292 18236 21304
rect 18288 21292 18294 21344
rect 23124 21332 23152 21440
rect 23937 21437 23949 21471
rect 23983 21437 23995 21471
rect 23937 21431 23995 21437
rect 24213 21471 24271 21477
rect 24213 21437 24225 21471
rect 24259 21468 24271 21471
rect 24302 21468 24308 21480
rect 24259 21440 24308 21468
rect 24259 21437 24271 21440
rect 24213 21431 24271 21437
rect 23952 21400 23980 21431
rect 24302 21428 24308 21440
rect 24360 21428 24366 21480
rect 24412 21468 24440 21508
rect 24854 21496 24860 21548
rect 24912 21536 24918 21548
rect 24949 21539 25007 21545
rect 24949 21536 24961 21539
rect 24912 21508 24961 21536
rect 24912 21496 24918 21508
rect 24949 21505 24961 21508
rect 24995 21536 25007 21539
rect 25038 21536 25044 21548
rect 24995 21508 25044 21536
rect 24995 21505 25007 21508
rect 24949 21499 25007 21505
rect 25038 21496 25044 21508
rect 25096 21496 25102 21548
rect 25148 21545 25176 21576
rect 25240 21576 25596 21604
rect 25240 21545 25268 21576
rect 25590 21564 25596 21576
rect 25648 21564 25654 21616
rect 25133 21539 25191 21545
rect 25133 21505 25145 21539
rect 25179 21505 25191 21539
rect 25133 21499 25191 21505
rect 25225 21539 25283 21545
rect 25225 21505 25237 21539
rect 25271 21505 25283 21539
rect 25225 21499 25283 21505
rect 25314 21496 25320 21548
rect 25372 21536 25378 21548
rect 25501 21539 25559 21545
rect 25501 21536 25513 21539
rect 25372 21508 25513 21536
rect 25372 21496 25378 21508
rect 25501 21505 25513 21508
rect 25547 21536 25559 21539
rect 25682 21536 25688 21548
rect 25547 21508 25688 21536
rect 25547 21505 25559 21508
rect 25501 21499 25559 21505
rect 25682 21496 25688 21508
rect 25740 21496 25746 21548
rect 27341 21539 27399 21545
rect 27341 21505 27353 21539
rect 27387 21536 27399 21539
rect 27430 21536 27436 21548
rect 27387 21508 27436 21536
rect 27387 21505 27399 21508
rect 27341 21499 27399 21505
rect 27430 21496 27436 21508
rect 27488 21496 27494 21548
rect 27798 21536 27804 21548
rect 27759 21508 27804 21536
rect 27798 21496 27804 21508
rect 27856 21536 27862 21548
rect 28166 21536 28172 21548
rect 27856 21508 28172 21536
rect 27856 21496 27862 21508
rect 28166 21496 28172 21508
rect 28224 21496 28230 21548
rect 25409 21471 25467 21477
rect 25409 21468 25421 21471
rect 24412 21440 25421 21468
rect 25409 21437 25421 21440
rect 25455 21468 25467 21471
rect 26970 21468 26976 21480
rect 25455 21440 26976 21468
rect 25455 21437 25467 21440
rect 25409 21431 25467 21437
rect 26970 21428 26976 21440
rect 27028 21428 27034 21480
rect 25314 21400 25320 21412
rect 23952 21372 25320 21400
rect 25314 21360 25320 21372
rect 25372 21360 25378 21412
rect 24026 21332 24032 21344
rect 23124 21304 24032 21332
rect 24026 21292 24032 21304
rect 24084 21292 24090 21344
rect 24949 21335 25007 21341
rect 24949 21301 24961 21335
rect 24995 21332 25007 21335
rect 25130 21332 25136 21344
rect 24995 21304 25136 21332
rect 24995 21301 25007 21304
rect 24949 21295 25007 21301
rect 25130 21292 25136 21304
rect 25188 21292 25194 21344
rect 26694 21292 26700 21344
rect 26752 21332 26758 21344
rect 27249 21335 27307 21341
rect 27249 21332 27261 21335
rect 26752 21304 27261 21332
rect 26752 21292 26758 21304
rect 27249 21301 27261 21304
rect 27295 21301 27307 21335
rect 27249 21295 27307 21301
rect 1104 21242 28888 21264
rect 1104 21190 4423 21242
rect 4475 21190 4487 21242
rect 4539 21190 4551 21242
rect 4603 21190 4615 21242
rect 4667 21190 4679 21242
rect 4731 21190 11369 21242
rect 11421 21190 11433 21242
rect 11485 21190 11497 21242
rect 11549 21190 11561 21242
rect 11613 21190 11625 21242
rect 11677 21190 18315 21242
rect 18367 21190 18379 21242
rect 18431 21190 18443 21242
rect 18495 21190 18507 21242
rect 18559 21190 18571 21242
rect 18623 21190 25261 21242
rect 25313 21190 25325 21242
rect 25377 21190 25389 21242
rect 25441 21190 25453 21242
rect 25505 21190 25517 21242
rect 25569 21190 28888 21242
rect 1104 21168 28888 21190
rect 20257 21063 20315 21069
rect 20257 21029 20269 21063
rect 20303 21029 20315 21063
rect 20257 21023 20315 21029
rect 20272 20992 20300 21023
rect 19628 20964 20300 20992
rect 20901 20995 20959 21001
rect 16022 20924 16028 20936
rect 15983 20896 16028 20924
rect 16022 20884 16028 20896
rect 16080 20884 16086 20936
rect 19628 20933 19656 20964
rect 20901 20961 20913 20995
rect 20947 20992 20959 20995
rect 21634 20992 21640 21004
rect 20947 20964 21640 20992
rect 20947 20961 20959 20964
rect 20901 20955 20959 20961
rect 21634 20952 21640 20964
rect 21692 20952 21698 21004
rect 23382 20992 23388 21004
rect 23343 20964 23388 20992
rect 23382 20952 23388 20964
rect 23440 20952 23446 21004
rect 26513 20995 26571 21001
rect 26513 20961 26525 20995
rect 26559 20992 26571 20995
rect 27706 20992 27712 21004
rect 26559 20964 27712 20992
rect 26559 20961 26571 20964
rect 26513 20955 26571 20961
rect 27706 20952 27712 20964
rect 27764 20952 27770 21004
rect 28350 20992 28356 21004
rect 28311 20964 28356 20992
rect 28350 20952 28356 20964
rect 28408 20952 28414 21004
rect 18693 20927 18751 20933
rect 18693 20893 18705 20927
rect 18739 20924 18751 20927
rect 19429 20927 19487 20933
rect 19429 20924 19441 20927
rect 18739 20896 19441 20924
rect 18739 20893 18751 20896
rect 18693 20887 18751 20893
rect 19429 20893 19441 20896
rect 19475 20893 19487 20927
rect 19429 20887 19487 20893
rect 19613 20927 19671 20933
rect 19613 20893 19625 20927
rect 19659 20893 19671 20927
rect 19613 20887 19671 20893
rect 19797 20927 19855 20933
rect 19797 20893 19809 20927
rect 19843 20924 19855 20927
rect 20530 20924 20536 20936
rect 19843 20896 20536 20924
rect 19843 20893 19855 20896
rect 19797 20887 19855 20893
rect 19334 20816 19340 20868
rect 19392 20856 19398 20868
rect 19812 20856 19840 20887
rect 20530 20884 20536 20896
rect 20588 20884 20594 20936
rect 23106 20884 23112 20936
rect 23164 20933 23170 20936
rect 23164 20924 23176 20933
rect 23164 20896 23209 20924
rect 23164 20887 23176 20896
rect 23164 20884 23170 20887
rect 19392 20828 19840 20856
rect 26697 20859 26755 20865
rect 19392 20816 19398 20828
rect 26697 20825 26709 20859
rect 26743 20856 26755 20859
rect 27338 20856 27344 20868
rect 26743 20828 27344 20856
rect 26743 20825 26755 20828
rect 26697 20819 26755 20825
rect 27338 20816 27344 20828
rect 27396 20816 27402 20868
rect 16209 20791 16267 20797
rect 16209 20757 16221 20791
rect 16255 20788 16267 20791
rect 16942 20788 16948 20800
rect 16255 20760 16948 20788
rect 16255 20757 16267 20760
rect 16209 20751 16267 20757
rect 16942 20748 16948 20760
rect 17000 20748 17006 20800
rect 18877 20791 18935 20797
rect 18877 20757 18889 20791
rect 18923 20788 18935 20791
rect 19518 20788 19524 20800
rect 18923 20760 19524 20788
rect 18923 20757 18935 20760
rect 18877 20751 18935 20757
rect 19518 20748 19524 20760
rect 19576 20748 19582 20800
rect 20346 20748 20352 20800
rect 20404 20788 20410 20800
rect 20625 20791 20683 20797
rect 20625 20788 20637 20791
rect 20404 20760 20637 20788
rect 20404 20748 20410 20760
rect 20625 20757 20637 20760
rect 20671 20757 20683 20791
rect 20625 20751 20683 20757
rect 20717 20791 20775 20797
rect 20717 20757 20729 20791
rect 20763 20788 20775 20791
rect 22002 20788 22008 20800
rect 20763 20760 22008 20788
rect 20763 20757 20775 20760
rect 20717 20751 20775 20757
rect 22002 20748 22008 20760
rect 22060 20748 22066 20800
rect 1104 20698 29048 20720
rect 1104 20646 7896 20698
rect 7948 20646 7960 20698
rect 8012 20646 8024 20698
rect 8076 20646 8088 20698
rect 8140 20646 8152 20698
rect 8204 20646 14842 20698
rect 14894 20646 14906 20698
rect 14958 20646 14970 20698
rect 15022 20646 15034 20698
rect 15086 20646 15098 20698
rect 15150 20646 21788 20698
rect 21840 20646 21852 20698
rect 21904 20646 21916 20698
rect 21968 20646 21980 20698
rect 22032 20646 22044 20698
rect 22096 20646 28734 20698
rect 28786 20646 28798 20698
rect 28850 20646 28862 20698
rect 28914 20646 28926 20698
rect 28978 20646 28990 20698
rect 29042 20646 29048 20698
rect 1104 20624 29048 20646
rect 15841 20587 15899 20593
rect 15841 20553 15853 20587
rect 15887 20584 15899 20587
rect 16022 20584 16028 20596
rect 15887 20556 16028 20584
rect 15887 20553 15899 20556
rect 15841 20547 15899 20553
rect 16022 20544 16028 20556
rect 16080 20544 16086 20596
rect 25682 20544 25688 20596
rect 25740 20584 25746 20596
rect 27341 20587 27399 20593
rect 27341 20584 27353 20587
rect 25740 20556 27353 20584
rect 25740 20544 25746 20556
rect 27341 20553 27353 20556
rect 27387 20553 27399 20587
rect 27341 20547 27399 20553
rect 18230 20516 18236 20528
rect 16868 20488 18236 20516
rect 1949 20451 2007 20457
rect 1949 20417 1961 20451
rect 1995 20448 2007 20451
rect 2038 20448 2044 20460
rect 1995 20420 2044 20448
rect 1995 20417 2007 20420
rect 1949 20411 2007 20417
rect 2038 20408 2044 20420
rect 2096 20408 2102 20460
rect 15194 20408 15200 20460
rect 15252 20448 15258 20460
rect 15473 20451 15531 20457
rect 15473 20448 15485 20451
rect 15252 20420 15485 20448
rect 15252 20408 15258 20420
rect 15473 20417 15485 20420
rect 15519 20417 15531 20451
rect 15473 20411 15531 20417
rect 15654 20408 15660 20460
rect 15712 20448 15718 20460
rect 15838 20448 15844 20460
rect 15712 20420 15844 20448
rect 15712 20408 15718 20420
rect 15838 20408 15844 20420
rect 15896 20408 15902 20460
rect 16868 20457 16896 20488
rect 18230 20476 18236 20488
rect 18288 20476 18294 20528
rect 19518 20525 19524 20528
rect 19512 20516 19524 20525
rect 19479 20488 19524 20516
rect 19512 20479 19524 20488
rect 19518 20476 19524 20479
rect 19576 20476 19582 20528
rect 25492 20519 25550 20525
rect 25492 20485 25504 20519
rect 25538 20516 25550 20519
rect 25590 20516 25596 20528
rect 25538 20488 25596 20516
rect 25538 20485 25550 20488
rect 25492 20479 25550 20485
rect 25590 20476 25596 20488
rect 25648 20476 25654 20528
rect 16853 20451 16911 20457
rect 16853 20417 16865 20451
rect 16899 20417 16911 20451
rect 16853 20411 16911 20417
rect 16942 20408 16948 20460
rect 17000 20448 17006 20460
rect 17109 20451 17167 20457
rect 17109 20448 17121 20451
rect 17000 20420 17121 20448
rect 17000 20408 17006 20420
rect 17109 20417 17121 20420
rect 17155 20417 17167 20451
rect 18248 20448 18276 20476
rect 19245 20451 19303 20457
rect 19245 20448 19257 20451
rect 18248 20420 19257 20448
rect 17109 20411 17167 20417
rect 19245 20417 19257 20420
rect 19291 20417 19303 20451
rect 27157 20451 27215 20457
rect 27157 20448 27169 20451
rect 19245 20411 19303 20417
rect 26620 20420 27169 20448
rect 23474 20340 23480 20392
rect 23532 20380 23538 20392
rect 25225 20383 25283 20389
rect 25225 20380 25237 20383
rect 23532 20352 25237 20380
rect 23532 20340 23538 20352
rect 25225 20349 25237 20352
rect 25271 20349 25283 20383
rect 25225 20343 25283 20349
rect 26620 20321 26648 20420
rect 27157 20417 27169 20420
rect 27203 20417 27215 20451
rect 27157 20411 27215 20417
rect 26605 20315 26663 20321
rect 26605 20281 26617 20315
rect 26651 20281 26663 20315
rect 26605 20275 26663 20281
rect 1762 20204 1768 20256
rect 1820 20244 1826 20256
rect 1857 20247 1915 20253
rect 1857 20244 1869 20247
rect 1820 20216 1869 20244
rect 1820 20204 1826 20216
rect 1857 20213 1869 20216
rect 1903 20213 1915 20247
rect 1857 20207 1915 20213
rect 15286 20204 15292 20256
rect 15344 20244 15350 20256
rect 18233 20247 18291 20253
rect 18233 20244 18245 20247
rect 15344 20216 18245 20244
rect 15344 20204 15350 20216
rect 18233 20213 18245 20216
rect 18279 20213 18291 20247
rect 18233 20207 18291 20213
rect 20346 20204 20352 20256
rect 20404 20244 20410 20256
rect 20625 20247 20683 20253
rect 20625 20244 20637 20247
rect 20404 20216 20637 20244
rect 20404 20204 20410 20216
rect 20625 20213 20637 20216
rect 20671 20213 20683 20247
rect 27890 20244 27896 20256
rect 27851 20216 27896 20244
rect 20625 20207 20683 20213
rect 27890 20204 27896 20216
rect 27948 20204 27954 20256
rect 1104 20154 28888 20176
rect 1104 20102 4423 20154
rect 4475 20102 4487 20154
rect 4539 20102 4551 20154
rect 4603 20102 4615 20154
rect 4667 20102 4679 20154
rect 4731 20102 11369 20154
rect 11421 20102 11433 20154
rect 11485 20102 11497 20154
rect 11549 20102 11561 20154
rect 11613 20102 11625 20154
rect 11677 20102 18315 20154
rect 18367 20102 18379 20154
rect 18431 20102 18443 20154
rect 18495 20102 18507 20154
rect 18559 20102 18571 20154
rect 18623 20102 25261 20154
rect 25313 20102 25325 20154
rect 25377 20102 25389 20154
rect 25441 20102 25453 20154
rect 25505 20102 25517 20154
rect 25569 20102 28888 20154
rect 1104 20080 28888 20102
rect 15194 20040 15200 20052
rect 15155 20012 15200 20040
rect 15194 20000 15200 20012
rect 15252 20000 15258 20052
rect 24670 19972 24676 19984
rect 21652 19944 24676 19972
rect 1762 19904 1768 19916
rect 1723 19876 1768 19904
rect 1762 19864 1768 19876
rect 1820 19864 1826 19916
rect 2774 19904 2780 19916
rect 2735 19876 2780 19904
rect 2774 19864 2780 19876
rect 2832 19864 2838 19916
rect 15470 19864 15476 19916
rect 15528 19904 15534 19916
rect 15749 19907 15807 19913
rect 15749 19904 15761 19907
rect 15528 19876 15761 19904
rect 15528 19864 15534 19876
rect 15749 19873 15761 19876
rect 15795 19873 15807 19907
rect 15749 19867 15807 19873
rect 1578 19836 1584 19848
rect 1539 19808 1584 19836
rect 1578 19796 1584 19808
rect 1636 19796 1642 19848
rect 15286 19796 15292 19848
rect 15344 19836 15350 19848
rect 15565 19839 15623 19845
rect 15565 19836 15577 19839
rect 15344 19808 15577 19836
rect 15344 19796 15350 19808
rect 15565 19805 15577 19808
rect 15611 19805 15623 19839
rect 21450 19836 21456 19848
rect 21411 19808 21456 19836
rect 15565 19799 15623 19805
rect 21450 19796 21456 19808
rect 21508 19796 21514 19848
rect 21652 19845 21680 19944
rect 24670 19932 24676 19944
rect 24728 19932 24734 19984
rect 24486 19864 24492 19916
rect 24544 19904 24550 19916
rect 26513 19907 26571 19913
rect 24544 19876 25268 19904
rect 24544 19864 24550 19876
rect 25240 19848 25268 19876
rect 26513 19873 26525 19907
rect 26559 19904 26571 19907
rect 27890 19904 27896 19916
rect 26559 19876 27896 19904
rect 26559 19873 26571 19876
rect 26513 19867 26571 19873
rect 27890 19864 27896 19876
rect 27948 19864 27954 19916
rect 28350 19904 28356 19916
rect 28311 19876 28356 19904
rect 28350 19864 28356 19876
rect 28408 19864 28414 19916
rect 21637 19839 21695 19845
rect 21637 19805 21649 19839
rect 21683 19805 21695 19839
rect 21637 19799 21695 19805
rect 21729 19839 21787 19845
rect 21729 19805 21741 19839
rect 21775 19805 21787 19839
rect 21729 19799 21787 19805
rect 14366 19728 14372 19780
rect 14424 19768 14430 19780
rect 21174 19768 21180 19780
rect 14424 19740 21180 19768
rect 14424 19728 14430 19740
rect 21174 19728 21180 19740
rect 21232 19728 21238 19780
rect 21744 19768 21772 19799
rect 21818 19796 21824 19848
rect 21876 19836 21882 19848
rect 22462 19836 22468 19848
rect 21876 19808 22468 19836
rect 21876 19796 21882 19808
rect 22462 19796 22468 19808
rect 22520 19796 22526 19848
rect 24762 19836 24768 19848
rect 24723 19808 24768 19836
rect 24762 19796 24768 19808
rect 24820 19796 24826 19848
rect 25038 19836 25044 19848
rect 24999 19808 25044 19836
rect 25038 19796 25044 19808
rect 25096 19796 25102 19848
rect 25222 19836 25228 19848
rect 25183 19808 25228 19836
rect 25222 19796 25228 19808
rect 25280 19796 25286 19848
rect 22370 19768 22376 19780
rect 21744 19740 22376 19768
rect 22370 19728 22376 19740
rect 22428 19728 22434 19780
rect 26694 19768 26700 19780
rect 26655 19740 26700 19768
rect 26694 19728 26700 19740
rect 26752 19728 26758 19780
rect 15654 19660 15660 19712
rect 15712 19700 15718 19712
rect 22097 19703 22155 19709
rect 15712 19672 15757 19700
rect 15712 19660 15718 19672
rect 22097 19669 22109 19703
rect 22143 19700 22155 19703
rect 23198 19700 23204 19712
rect 22143 19672 23204 19700
rect 22143 19669 22155 19672
rect 22097 19663 22155 19669
rect 23198 19660 23204 19672
rect 23256 19660 23262 19712
rect 24581 19703 24639 19709
rect 24581 19669 24593 19703
rect 24627 19700 24639 19703
rect 24854 19700 24860 19712
rect 24627 19672 24860 19700
rect 24627 19669 24639 19672
rect 24581 19663 24639 19669
rect 24854 19660 24860 19672
rect 24912 19660 24918 19712
rect 1104 19610 29048 19632
rect 1104 19558 7896 19610
rect 7948 19558 7960 19610
rect 8012 19558 8024 19610
rect 8076 19558 8088 19610
rect 8140 19558 8152 19610
rect 8204 19558 14842 19610
rect 14894 19558 14906 19610
rect 14958 19558 14970 19610
rect 15022 19558 15034 19610
rect 15086 19558 15098 19610
rect 15150 19558 21788 19610
rect 21840 19558 21852 19610
rect 21904 19558 21916 19610
rect 21968 19558 21980 19610
rect 22032 19558 22044 19610
rect 22096 19558 28734 19610
rect 28786 19558 28798 19610
rect 28850 19558 28862 19610
rect 28914 19558 28926 19610
rect 28978 19558 28990 19610
rect 29042 19558 29048 19610
rect 1104 19536 29048 19558
rect 16666 19456 16672 19508
rect 16724 19496 16730 19508
rect 16945 19499 17003 19505
rect 16945 19496 16957 19499
rect 16724 19468 16957 19496
rect 16724 19456 16730 19468
rect 16945 19465 16957 19468
rect 16991 19465 17003 19499
rect 16945 19459 17003 19465
rect 18075 19499 18133 19505
rect 18075 19465 18087 19499
rect 18121 19496 18133 19499
rect 18693 19499 18751 19505
rect 18693 19496 18705 19499
rect 18121 19468 18705 19496
rect 18121 19465 18133 19468
rect 18075 19459 18133 19465
rect 18693 19465 18705 19468
rect 18739 19465 18751 19499
rect 18693 19459 18751 19465
rect 22097 19499 22155 19505
rect 22097 19465 22109 19499
rect 22143 19496 22155 19499
rect 22462 19496 22468 19508
rect 22143 19468 22468 19496
rect 22143 19465 22155 19468
rect 22097 19459 22155 19465
rect 22462 19456 22468 19468
rect 22520 19456 22526 19508
rect 25590 19496 25596 19508
rect 25551 19468 25596 19496
rect 25590 19456 25596 19468
rect 25648 19456 25654 19508
rect 27338 19496 27344 19508
rect 27299 19468 27344 19496
rect 27338 19456 27344 19468
rect 27396 19456 27402 19508
rect 16209 19431 16267 19437
rect 16209 19397 16221 19431
rect 16255 19428 16267 19431
rect 17218 19428 17224 19440
rect 16255 19400 17224 19428
rect 16255 19397 16267 19400
rect 16209 19391 16267 19397
rect 17218 19388 17224 19400
rect 17276 19388 17282 19440
rect 17865 19431 17923 19437
rect 17865 19397 17877 19431
rect 17911 19428 17923 19431
rect 18874 19428 18880 19440
rect 17911 19400 18880 19428
rect 17911 19397 17923 19400
rect 17865 19391 17923 19397
rect 18874 19388 18880 19400
rect 18932 19388 18938 19440
rect 22278 19428 22284 19440
rect 20824 19400 22284 19428
rect 1578 19320 1584 19372
rect 1636 19360 1642 19372
rect 1673 19363 1731 19369
rect 1673 19360 1685 19363
rect 1636 19332 1685 19360
rect 1636 19320 1642 19332
rect 1673 19329 1685 19332
rect 1719 19329 1731 19363
rect 16114 19360 16120 19372
rect 16075 19332 16120 19360
rect 1673 19323 1731 19329
rect 16114 19320 16120 19332
rect 16172 19320 16178 19372
rect 16850 19360 16856 19372
rect 16811 19332 16856 19360
rect 16850 19320 16856 19332
rect 16908 19320 16914 19372
rect 17129 19363 17187 19369
rect 17129 19329 17141 19363
rect 17175 19360 17187 19363
rect 17402 19360 17408 19372
rect 17175 19332 17408 19360
rect 17175 19329 17187 19332
rect 17129 19323 17187 19329
rect 17402 19320 17408 19332
rect 17460 19320 17466 19372
rect 18966 19360 18972 19372
rect 17512 19332 18972 19360
rect 17129 19227 17187 19233
rect 17129 19193 17141 19227
rect 17175 19224 17187 19227
rect 17512 19224 17540 19332
rect 18966 19320 18972 19332
rect 19024 19320 19030 19372
rect 19061 19363 19119 19369
rect 19061 19329 19073 19363
rect 19107 19360 19119 19363
rect 19702 19360 19708 19372
rect 19107 19332 19380 19360
rect 19663 19332 19708 19360
rect 19107 19329 19119 19332
rect 19061 19323 19119 19329
rect 18878 19295 18936 19301
rect 18878 19261 18890 19295
rect 18924 19261 18936 19295
rect 18878 19255 18936 19261
rect 18690 19224 18696 19236
rect 17175 19196 17540 19224
rect 18064 19196 18696 19224
rect 17175 19193 17187 19196
rect 17129 19187 17187 19193
rect 18064 19165 18092 19196
rect 18690 19184 18696 19196
rect 18748 19184 18754 19236
rect 18782 19184 18788 19236
rect 18840 19224 18846 19236
rect 18892 19224 18920 19255
rect 19150 19252 19156 19304
rect 19208 19292 19214 19304
rect 19352 19292 19380 19332
rect 19702 19320 19708 19332
rect 19760 19320 19766 19372
rect 20625 19363 20683 19369
rect 20625 19329 20637 19363
rect 20671 19360 20683 19363
rect 20714 19360 20720 19372
rect 20671 19332 20720 19360
rect 20671 19329 20683 19332
rect 20625 19323 20683 19329
rect 20714 19320 20720 19332
rect 20772 19320 20778 19372
rect 20824 19369 20852 19400
rect 22278 19388 22284 19400
rect 22336 19388 22342 19440
rect 23198 19388 23204 19440
rect 23256 19437 23262 19440
rect 23256 19428 23268 19437
rect 23256 19400 23301 19428
rect 23256 19391 23268 19400
rect 23256 19388 23262 19391
rect 25038 19388 25044 19440
rect 25096 19428 25102 19440
rect 25096 19400 25268 19428
rect 25096 19388 25102 19400
rect 20809 19363 20867 19369
rect 20809 19329 20821 19363
rect 20855 19329 20867 19363
rect 20809 19323 20867 19329
rect 21174 19320 21180 19372
rect 21232 19360 21238 19372
rect 21269 19363 21327 19369
rect 21269 19360 21281 19363
rect 21232 19332 21281 19360
rect 21232 19320 21238 19332
rect 21269 19329 21281 19332
rect 21315 19329 21327 19363
rect 21269 19323 21327 19329
rect 21361 19363 21419 19369
rect 21361 19329 21373 19363
rect 21407 19360 21419 19363
rect 22094 19360 22100 19372
rect 21407 19332 22100 19360
rect 21407 19329 21419 19332
rect 21361 19323 21419 19329
rect 22094 19320 22100 19332
rect 22152 19320 22158 19372
rect 23474 19360 23480 19372
rect 23435 19332 23480 19360
rect 23474 19320 23480 19332
rect 23532 19320 23538 19372
rect 24670 19320 24676 19372
rect 24728 19360 24734 19372
rect 24949 19363 25007 19369
rect 24949 19360 24961 19363
rect 24728 19332 24961 19360
rect 24728 19320 24734 19332
rect 24949 19329 24961 19332
rect 24995 19329 25007 19363
rect 25130 19360 25136 19372
rect 25091 19332 25136 19360
rect 24949 19323 25007 19329
rect 25130 19320 25136 19332
rect 25188 19320 25194 19372
rect 25240 19369 25268 19400
rect 25225 19363 25283 19369
rect 25225 19329 25237 19363
rect 25271 19329 25283 19363
rect 25225 19323 25283 19329
rect 25317 19363 25375 19369
rect 25317 19329 25329 19363
rect 25363 19360 25375 19363
rect 25682 19360 25688 19372
rect 25363 19332 25688 19360
rect 25363 19329 25375 19332
rect 25317 19323 25375 19329
rect 25682 19320 25688 19332
rect 25740 19320 25746 19372
rect 27246 19320 27252 19372
rect 27304 19360 27310 19372
rect 27433 19363 27491 19369
rect 27433 19360 27445 19363
rect 27304 19332 27445 19360
rect 27304 19320 27310 19332
rect 27433 19329 27445 19332
rect 27479 19360 27491 19363
rect 27798 19360 27804 19372
rect 27479 19332 27804 19360
rect 27479 19329 27491 19332
rect 27433 19323 27491 19329
rect 27798 19320 27804 19332
rect 27856 19320 27862 19372
rect 19610 19292 19616 19304
rect 19208 19264 19253 19292
rect 19352 19264 19616 19292
rect 19208 19252 19214 19264
rect 19610 19252 19616 19264
rect 19668 19252 19674 19304
rect 19794 19252 19800 19304
rect 19852 19292 19858 19304
rect 19981 19295 20039 19301
rect 19981 19292 19993 19295
rect 19852 19264 19993 19292
rect 19852 19252 19858 19264
rect 19981 19261 19993 19264
rect 20027 19261 20039 19295
rect 19981 19255 20039 19261
rect 20070 19252 20076 19304
rect 20128 19292 20134 19304
rect 20128 19264 20668 19292
rect 20128 19252 20134 19264
rect 20640 19233 20668 19264
rect 27706 19252 27712 19304
rect 27764 19292 27770 19304
rect 27893 19295 27951 19301
rect 27893 19292 27905 19295
rect 27764 19264 27905 19292
rect 27764 19252 27770 19264
rect 27893 19261 27905 19264
rect 27939 19261 27951 19295
rect 27893 19255 27951 19261
rect 19889 19227 19947 19233
rect 19889 19224 19901 19227
rect 18840 19196 18920 19224
rect 19168 19196 19901 19224
rect 18840 19184 18846 19196
rect 19168 19168 19196 19196
rect 19889 19193 19901 19196
rect 19935 19193 19947 19227
rect 19889 19187 19947 19193
rect 20625 19227 20683 19233
rect 20625 19193 20637 19227
rect 20671 19193 20683 19227
rect 20625 19187 20683 19193
rect 18049 19159 18107 19165
rect 18049 19125 18061 19159
rect 18095 19125 18107 19159
rect 18049 19119 18107 19125
rect 18138 19116 18144 19168
rect 18196 19156 18202 19168
rect 18233 19159 18291 19165
rect 18233 19156 18245 19159
rect 18196 19128 18245 19156
rect 18196 19116 18202 19128
rect 18233 19125 18245 19128
rect 18279 19125 18291 19159
rect 18233 19119 18291 19125
rect 19150 19116 19156 19168
rect 19208 19116 19214 19168
rect 19242 19116 19248 19168
rect 19300 19156 19306 19168
rect 19797 19159 19855 19165
rect 19797 19156 19809 19159
rect 19300 19128 19809 19156
rect 19300 19116 19306 19128
rect 19797 19125 19809 19128
rect 19843 19156 19855 19159
rect 19978 19156 19984 19168
rect 19843 19128 19984 19156
rect 19843 19125 19855 19128
rect 19797 19119 19855 19125
rect 19978 19116 19984 19128
rect 20036 19116 20042 19168
rect 1104 19066 28888 19088
rect 1104 19014 4423 19066
rect 4475 19014 4487 19066
rect 4539 19014 4551 19066
rect 4603 19014 4615 19066
rect 4667 19014 4679 19066
rect 4731 19014 11369 19066
rect 11421 19014 11433 19066
rect 11485 19014 11497 19066
rect 11549 19014 11561 19066
rect 11613 19014 11625 19066
rect 11677 19014 18315 19066
rect 18367 19014 18379 19066
rect 18431 19014 18443 19066
rect 18495 19014 18507 19066
rect 18559 19014 18571 19066
rect 18623 19014 25261 19066
rect 25313 19014 25325 19066
rect 25377 19014 25389 19066
rect 25441 19014 25453 19066
rect 25505 19014 25517 19066
rect 25569 19014 28888 19066
rect 1104 18992 28888 19014
rect 18046 18952 18052 18964
rect 17052 18924 18052 18952
rect 1578 18748 1584 18760
rect 1539 18720 1584 18748
rect 1578 18708 1584 18720
rect 1636 18708 1642 18760
rect 17052 18757 17080 18924
rect 18046 18912 18052 18924
rect 18104 18912 18110 18964
rect 18432 18924 18736 18952
rect 17313 18887 17371 18893
rect 17313 18853 17325 18887
rect 17359 18884 17371 18887
rect 18432 18884 18460 18924
rect 17359 18856 18460 18884
rect 18708 18884 18736 18924
rect 18782 18912 18788 18964
rect 18840 18952 18846 18964
rect 19242 18952 19248 18964
rect 18840 18924 19248 18952
rect 18840 18912 18846 18924
rect 19242 18912 19248 18924
rect 19300 18912 19306 18964
rect 19521 18955 19579 18961
rect 19521 18921 19533 18955
rect 19567 18952 19579 18955
rect 19702 18952 19708 18964
rect 19567 18924 19708 18952
rect 19567 18921 19579 18924
rect 19521 18915 19579 18921
rect 19702 18912 19708 18924
rect 19760 18912 19766 18964
rect 27522 18952 27528 18964
rect 22066 18924 27528 18952
rect 22066 18884 22094 18924
rect 27522 18912 27528 18924
rect 27580 18952 27586 18964
rect 27709 18955 27767 18961
rect 27709 18952 27721 18955
rect 27580 18924 27721 18952
rect 27580 18912 27586 18924
rect 27709 18921 27721 18924
rect 27755 18921 27767 18955
rect 27709 18915 27767 18921
rect 18708 18856 22094 18884
rect 17359 18853 17371 18856
rect 17313 18847 17371 18853
rect 17954 18776 17960 18828
rect 18012 18816 18018 18828
rect 18012 18788 18552 18816
rect 18012 18776 18018 18788
rect 17037 18751 17095 18757
rect 17037 18717 17049 18751
rect 17083 18717 17095 18751
rect 17037 18711 17095 18717
rect 17129 18751 17187 18757
rect 17129 18717 17141 18751
rect 17175 18748 17187 18751
rect 17218 18748 17224 18760
rect 17175 18720 17224 18748
rect 17175 18717 17187 18720
rect 17129 18711 17187 18717
rect 17218 18708 17224 18720
rect 17276 18708 17282 18760
rect 17405 18751 17463 18757
rect 17405 18717 17417 18751
rect 17451 18748 17463 18751
rect 17678 18748 17684 18760
rect 17451 18720 17684 18748
rect 17451 18717 17463 18720
rect 17405 18711 17463 18717
rect 17678 18708 17684 18720
rect 17736 18708 17742 18760
rect 18046 18748 18052 18760
rect 18007 18720 18052 18748
rect 18046 18708 18052 18720
rect 18104 18708 18110 18760
rect 18524 18757 18552 18788
rect 18708 18757 18736 18856
rect 23290 18844 23296 18896
rect 23348 18884 23354 18896
rect 23385 18887 23443 18893
rect 23385 18884 23397 18887
rect 23348 18856 23397 18884
rect 23348 18844 23354 18856
rect 23385 18853 23397 18856
rect 23431 18853 23443 18887
rect 23385 18847 23443 18853
rect 19334 18776 19340 18828
rect 19392 18816 19398 18828
rect 19794 18816 19800 18828
rect 19392 18788 19800 18816
rect 19392 18776 19398 18788
rect 19794 18776 19800 18788
rect 19852 18776 19858 18828
rect 22094 18776 22100 18828
rect 22152 18816 22158 18828
rect 22152 18788 22197 18816
rect 22152 18776 22158 18788
rect 22278 18776 22284 18828
rect 22336 18816 22342 18828
rect 23198 18816 23204 18828
rect 22336 18788 23204 18816
rect 22336 18776 22342 18788
rect 23198 18776 23204 18788
rect 23256 18816 23262 18828
rect 23753 18819 23811 18825
rect 23753 18816 23765 18819
rect 23256 18788 23765 18816
rect 23256 18776 23262 18788
rect 23753 18785 23765 18788
rect 23799 18785 23811 18819
rect 23753 18779 23811 18785
rect 24578 18776 24584 18828
rect 24636 18816 24642 18828
rect 26329 18819 26387 18825
rect 26329 18816 26341 18819
rect 24636 18788 26341 18816
rect 24636 18776 24642 18788
rect 26329 18785 26341 18788
rect 26375 18785 26387 18819
rect 26329 18779 26387 18785
rect 18509 18751 18567 18757
rect 18509 18717 18521 18751
rect 18555 18717 18567 18751
rect 18509 18711 18567 18717
rect 18693 18751 18751 18757
rect 18693 18717 18705 18751
rect 18739 18717 18751 18751
rect 18693 18711 18751 18717
rect 18966 18708 18972 18760
rect 19024 18748 19030 18760
rect 19429 18751 19487 18757
rect 19429 18748 19441 18751
rect 19024 18720 19441 18748
rect 19024 18708 19030 18720
rect 19429 18717 19441 18720
rect 19475 18717 19487 18751
rect 19610 18748 19616 18760
rect 19571 18720 19616 18748
rect 19429 18711 19487 18717
rect 19610 18708 19616 18720
rect 19668 18708 19674 18760
rect 24765 18751 24823 18757
rect 24765 18748 24777 18751
rect 22296 18720 24777 18748
rect 3326 18640 3332 18692
rect 3384 18680 3390 18692
rect 20441 18683 20499 18689
rect 20441 18680 20453 18683
rect 3384 18652 20453 18680
rect 3384 18640 3390 18652
rect 20441 18649 20453 18652
rect 20487 18649 20499 18683
rect 20441 18643 20499 18649
rect 20714 18640 20720 18692
rect 20772 18680 20778 18692
rect 22296 18680 22324 18720
rect 24765 18717 24777 18720
rect 24811 18748 24823 18751
rect 24946 18748 24952 18760
rect 24811 18720 24952 18748
rect 24811 18717 24823 18720
rect 24765 18711 24823 18717
rect 24946 18708 24952 18720
rect 25004 18708 25010 18760
rect 28350 18748 28356 18760
rect 28311 18720 28356 18748
rect 28350 18708 28356 18720
rect 28408 18708 28414 18760
rect 20772 18652 22324 18680
rect 20772 18640 20778 18652
rect 22370 18640 22376 18692
rect 22428 18680 22434 18692
rect 23382 18680 23388 18692
rect 22428 18652 23388 18680
rect 22428 18640 22434 18652
rect 23382 18640 23388 18652
rect 23440 18680 23446 18692
rect 24581 18683 24639 18689
rect 24581 18680 24593 18683
rect 23440 18652 24593 18680
rect 23440 18640 23446 18652
rect 24581 18649 24593 18652
rect 24627 18649 24639 18683
rect 24581 18643 24639 18649
rect 26596 18683 26654 18689
rect 26596 18649 26608 18683
rect 26642 18680 26654 18683
rect 27982 18680 27988 18692
rect 26642 18652 27988 18680
rect 26642 18649 26654 18652
rect 26596 18643 26654 18649
rect 27982 18640 27988 18652
rect 28040 18640 28046 18692
rect 1765 18615 1823 18621
rect 1765 18581 1777 18615
rect 1811 18612 1823 18615
rect 15654 18612 15660 18624
rect 1811 18584 15660 18612
rect 1811 18581 1823 18584
rect 1765 18575 1823 18581
rect 15654 18572 15660 18584
rect 15712 18572 15718 18624
rect 16853 18615 16911 18621
rect 16853 18581 16865 18615
rect 16899 18612 16911 18615
rect 17218 18612 17224 18624
rect 16899 18584 17224 18612
rect 16899 18581 16911 18584
rect 16853 18575 16911 18581
rect 17218 18572 17224 18584
rect 17276 18572 17282 18624
rect 17494 18572 17500 18624
rect 17552 18612 17558 18624
rect 17957 18615 18015 18621
rect 17957 18612 17969 18615
rect 17552 18584 17969 18612
rect 17552 18572 17558 18584
rect 17957 18581 17969 18584
rect 18003 18581 18015 18615
rect 18506 18612 18512 18624
rect 18467 18584 18512 18612
rect 17957 18575 18015 18581
rect 18506 18572 18512 18584
rect 18564 18572 18570 18624
rect 23293 18615 23351 18621
rect 23293 18581 23305 18615
rect 23339 18612 23351 18615
rect 23658 18612 23664 18624
rect 23339 18584 23664 18612
rect 23339 18581 23351 18584
rect 23293 18575 23351 18581
rect 23658 18572 23664 18584
rect 23716 18572 23722 18624
rect 1104 18522 29048 18544
rect 1104 18470 7896 18522
rect 7948 18470 7960 18522
rect 8012 18470 8024 18522
rect 8076 18470 8088 18522
rect 8140 18470 8152 18522
rect 8204 18470 14842 18522
rect 14894 18470 14906 18522
rect 14958 18470 14970 18522
rect 15022 18470 15034 18522
rect 15086 18470 15098 18522
rect 15150 18470 21788 18522
rect 21840 18470 21852 18522
rect 21904 18470 21916 18522
rect 21968 18470 21980 18522
rect 22032 18470 22044 18522
rect 22096 18470 28734 18522
rect 28786 18470 28798 18522
rect 28850 18470 28862 18522
rect 28914 18470 28926 18522
rect 28978 18470 28990 18522
rect 29042 18470 29048 18522
rect 1104 18448 29048 18470
rect 16850 18408 16856 18420
rect 16811 18380 16856 18408
rect 16850 18368 16856 18380
rect 16908 18368 16914 18420
rect 17218 18408 17224 18420
rect 17179 18380 17224 18408
rect 17218 18368 17224 18380
rect 17276 18368 17282 18420
rect 21177 18411 21235 18417
rect 21177 18377 21189 18411
rect 21223 18408 21235 18411
rect 21450 18408 21456 18420
rect 21223 18380 21456 18408
rect 21223 18377 21235 18380
rect 21177 18371 21235 18377
rect 21450 18368 21456 18380
rect 21508 18368 21514 18420
rect 23474 18368 23480 18420
rect 23532 18408 23538 18420
rect 24578 18408 24584 18420
rect 23532 18380 24584 18408
rect 23532 18368 23538 18380
rect 24578 18368 24584 18380
rect 24636 18408 24642 18420
rect 24673 18411 24731 18417
rect 24673 18408 24685 18411
rect 24636 18380 24685 18408
rect 24636 18368 24642 18380
rect 24673 18377 24685 18380
rect 24719 18377 24731 18411
rect 27982 18408 27988 18420
rect 27943 18380 27988 18408
rect 24673 18371 24731 18377
rect 27982 18368 27988 18380
rect 28040 18368 28046 18420
rect 18506 18340 18512 18352
rect 17144 18312 18512 18340
rect 17144 18284 17172 18312
rect 18506 18300 18512 18312
rect 18564 18300 18570 18352
rect 19981 18343 20039 18349
rect 19981 18309 19993 18343
rect 20027 18340 20039 18343
rect 22554 18340 22560 18352
rect 20027 18312 22560 18340
rect 20027 18309 20039 18312
rect 19981 18303 20039 18309
rect 22554 18300 22560 18312
rect 22612 18340 22618 18352
rect 23385 18343 23443 18349
rect 23385 18340 23397 18343
rect 22612 18312 23397 18340
rect 22612 18300 22618 18312
rect 23385 18309 23397 18312
rect 23431 18309 23443 18343
rect 23385 18303 23443 18309
rect 15654 18272 15660 18284
rect 15615 18244 15660 18272
rect 15654 18232 15660 18244
rect 15712 18232 15718 18284
rect 15838 18232 15844 18284
rect 15896 18272 15902 18284
rect 17126 18272 17132 18284
rect 15896 18244 15989 18272
rect 17039 18244 17132 18272
rect 15896 18232 15902 18244
rect 17126 18232 17132 18244
rect 17184 18232 17190 18284
rect 17310 18272 17316 18284
rect 17271 18244 17316 18272
rect 17310 18232 17316 18244
rect 17368 18232 17374 18284
rect 17494 18272 17500 18284
rect 17455 18244 17500 18272
rect 17494 18232 17500 18244
rect 17552 18232 17558 18284
rect 20714 18232 20720 18284
rect 20772 18272 20778 18284
rect 20809 18275 20867 18281
rect 20809 18272 20821 18275
rect 20772 18244 20821 18272
rect 20772 18232 20778 18244
rect 20809 18241 20821 18244
rect 20855 18241 20867 18275
rect 20809 18235 20867 18241
rect 20993 18275 21051 18281
rect 20993 18241 21005 18275
rect 21039 18272 21051 18275
rect 21039 18244 22094 18272
rect 21039 18241 21051 18244
rect 20993 18235 21051 18241
rect 15856 18136 15884 18232
rect 16206 18164 16212 18216
rect 16264 18204 16270 18216
rect 17589 18207 17647 18213
rect 17589 18204 17601 18207
rect 16264 18176 17601 18204
rect 16264 18164 16270 18176
rect 17589 18173 17601 18176
rect 17635 18173 17647 18207
rect 18230 18204 18236 18216
rect 18191 18176 18236 18204
rect 17589 18167 17647 18173
rect 18230 18164 18236 18176
rect 18288 18164 18294 18216
rect 22066 18204 22094 18244
rect 22186 18232 22192 18284
rect 22244 18272 22250 18284
rect 22741 18275 22799 18281
rect 22741 18272 22753 18275
rect 22244 18244 22753 18272
rect 22244 18232 22250 18244
rect 22741 18241 22753 18244
rect 22787 18241 22799 18275
rect 22741 18235 22799 18241
rect 22925 18275 22983 18281
rect 22925 18241 22937 18275
rect 22971 18272 22983 18275
rect 23842 18272 23848 18284
rect 22971 18244 23848 18272
rect 22971 18241 22983 18244
rect 22925 18235 22983 18241
rect 23842 18232 23848 18244
rect 23900 18232 23906 18284
rect 27338 18272 27344 18284
rect 27299 18244 27344 18272
rect 27338 18232 27344 18244
rect 27396 18232 27402 18284
rect 27525 18275 27583 18281
rect 27525 18241 27537 18275
rect 27571 18272 27583 18275
rect 28169 18275 28227 18281
rect 28169 18272 28181 18275
rect 27571 18244 28181 18272
rect 27571 18241 27583 18244
rect 27525 18235 27583 18241
rect 28169 18241 28181 18244
rect 28215 18241 28227 18275
rect 28169 18235 28227 18241
rect 22278 18204 22284 18216
rect 22066 18176 22284 18204
rect 22278 18164 22284 18176
rect 22336 18164 22342 18216
rect 26510 18164 26516 18216
rect 26568 18204 26574 18216
rect 27157 18207 27215 18213
rect 27157 18204 27169 18207
rect 26568 18176 27169 18204
rect 26568 18164 26574 18176
rect 27157 18173 27169 18176
rect 27203 18173 27215 18207
rect 27157 18167 27215 18173
rect 23934 18136 23940 18148
rect 15856 18108 23940 18136
rect 23934 18096 23940 18108
rect 23992 18096 23998 18148
rect 1578 18028 1584 18080
rect 1636 18068 1642 18080
rect 1673 18071 1731 18077
rect 1673 18068 1685 18071
rect 1636 18040 1685 18068
rect 1636 18028 1642 18040
rect 1673 18037 1685 18040
rect 1719 18037 1731 18071
rect 1673 18031 1731 18037
rect 16025 18071 16083 18077
rect 16025 18037 16037 18071
rect 16071 18068 16083 18071
rect 16850 18068 16856 18080
rect 16071 18040 16856 18068
rect 16071 18037 16083 18040
rect 16025 18031 16083 18037
rect 16850 18028 16856 18040
rect 16908 18028 16914 18080
rect 22925 18071 22983 18077
rect 22925 18037 22937 18071
rect 22971 18068 22983 18071
rect 23658 18068 23664 18080
rect 22971 18040 23664 18068
rect 22971 18037 22983 18040
rect 22925 18031 22983 18037
rect 23658 18028 23664 18040
rect 23716 18028 23722 18080
rect 1104 17978 28888 18000
rect 1104 17926 4423 17978
rect 4475 17926 4487 17978
rect 4539 17926 4551 17978
rect 4603 17926 4615 17978
rect 4667 17926 4679 17978
rect 4731 17926 11369 17978
rect 11421 17926 11433 17978
rect 11485 17926 11497 17978
rect 11549 17926 11561 17978
rect 11613 17926 11625 17978
rect 11677 17926 18315 17978
rect 18367 17926 18379 17978
rect 18431 17926 18443 17978
rect 18495 17926 18507 17978
rect 18559 17926 18571 17978
rect 18623 17926 25261 17978
rect 25313 17926 25325 17978
rect 25377 17926 25389 17978
rect 25441 17926 25453 17978
rect 25505 17926 25517 17978
rect 25569 17926 28888 17978
rect 1104 17904 28888 17926
rect 2222 17824 2228 17876
rect 2280 17864 2286 17876
rect 5166 17864 5172 17876
rect 2280 17836 5172 17864
rect 2280 17824 2286 17836
rect 5166 17824 5172 17836
rect 5224 17824 5230 17876
rect 15381 17867 15439 17873
rect 15381 17833 15393 17867
rect 15427 17864 15439 17867
rect 15654 17864 15660 17876
rect 15427 17836 15660 17864
rect 15427 17833 15439 17836
rect 15381 17827 15439 17833
rect 15654 17824 15660 17836
rect 15712 17824 15718 17876
rect 17126 17824 17132 17876
rect 17184 17864 17190 17876
rect 17221 17867 17279 17873
rect 17221 17864 17233 17867
rect 17184 17836 17233 17864
rect 17184 17824 17190 17836
rect 17221 17833 17233 17836
rect 17267 17833 17279 17867
rect 17402 17864 17408 17876
rect 17363 17836 17408 17864
rect 17221 17827 17279 17833
rect 17402 17824 17408 17836
rect 17460 17824 17466 17876
rect 18417 17867 18475 17873
rect 18417 17833 18429 17867
rect 18463 17833 18475 17867
rect 18417 17827 18475 17833
rect 1854 17756 1860 17808
rect 1912 17796 1918 17808
rect 1912 17768 15884 17796
rect 1912 17756 1918 17768
rect 1578 17728 1584 17740
rect 1539 17700 1584 17728
rect 1578 17688 1584 17700
rect 1636 17688 1642 17740
rect 2774 17728 2780 17740
rect 2735 17700 2780 17728
rect 2774 17688 2780 17700
rect 2832 17688 2838 17740
rect 15856 17737 15884 17768
rect 15841 17731 15899 17737
rect 15841 17697 15853 17731
rect 15887 17697 15899 17731
rect 15841 17691 15899 17697
rect 15930 17688 15936 17740
rect 15988 17728 15994 17740
rect 16853 17731 16911 17737
rect 15988 17700 16033 17728
rect 15988 17688 15994 17700
rect 16853 17697 16865 17731
rect 16899 17728 16911 17731
rect 17218 17728 17224 17740
rect 16899 17700 17224 17728
rect 16899 17697 16911 17700
rect 16853 17691 16911 17697
rect 17218 17688 17224 17700
rect 17276 17688 17282 17740
rect 18432 17728 18460 17827
rect 19610 17824 19616 17876
rect 19668 17864 19674 17876
rect 19705 17867 19763 17873
rect 19705 17864 19717 17867
rect 19668 17836 19717 17864
rect 19668 17824 19674 17836
rect 19705 17833 19717 17836
rect 19751 17833 19763 17867
rect 19705 17827 19763 17833
rect 24578 17728 24584 17740
rect 18432 17700 19472 17728
rect 24539 17700 24584 17728
rect 18690 17620 18696 17672
rect 18748 17660 18754 17672
rect 19444 17669 19472 17700
rect 24578 17688 24584 17700
rect 24636 17688 24642 17740
rect 26142 17688 26148 17740
rect 26200 17728 26206 17740
rect 26513 17731 26571 17737
rect 26513 17728 26525 17731
rect 26200 17700 26525 17728
rect 26200 17688 26206 17700
rect 26513 17697 26525 17700
rect 26559 17697 26571 17731
rect 28350 17728 28356 17740
rect 28311 17700 28356 17728
rect 26513 17691 26571 17697
rect 28350 17688 28356 17700
rect 28408 17688 28414 17740
rect 18785 17663 18843 17669
rect 18785 17660 18797 17663
rect 18748 17632 18797 17660
rect 18748 17620 18754 17632
rect 18785 17629 18797 17632
rect 18831 17629 18843 17663
rect 18785 17623 18843 17629
rect 19429 17663 19487 17669
rect 19429 17629 19441 17663
rect 19475 17660 19487 17663
rect 19886 17660 19892 17672
rect 19475 17632 19892 17660
rect 19475 17629 19487 17632
rect 19429 17623 19487 17629
rect 1765 17595 1823 17601
rect 1765 17561 1777 17595
rect 1811 17592 1823 17595
rect 1946 17592 1952 17604
rect 1811 17564 1952 17592
rect 1811 17561 1823 17564
rect 1765 17555 1823 17561
rect 1946 17552 1952 17564
rect 2004 17552 2010 17604
rect 17221 17595 17279 17601
rect 17221 17561 17233 17595
rect 17267 17592 17279 17595
rect 17310 17592 17316 17604
rect 17267 17564 17316 17592
rect 17267 17561 17279 17564
rect 17221 17555 17279 17561
rect 17310 17552 17316 17564
rect 17368 17592 17374 17604
rect 18800 17592 18828 17623
rect 19886 17620 19892 17632
rect 19944 17620 19950 17672
rect 22649 17663 22707 17669
rect 22649 17629 22661 17663
rect 22695 17660 22707 17663
rect 23109 17663 23167 17669
rect 23109 17660 23121 17663
rect 22695 17632 23121 17660
rect 22695 17629 22707 17632
rect 22649 17623 22707 17629
rect 23109 17629 23121 17632
rect 23155 17629 23167 17663
rect 23109 17623 23167 17629
rect 23198 17620 23204 17672
rect 23256 17660 23262 17672
rect 23293 17663 23351 17669
rect 23293 17660 23305 17663
rect 23256 17632 23305 17660
rect 23256 17620 23262 17632
rect 23293 17629 23305 17632
rect 23339 17629 23351 17663
rect 23293 17623 23351 17629
rect 23382 17620 23388 17672
rect 23440 17660 23446 17672
rect 24854 17669 24860 17672
rect 23477 17663 23535 17669
rect 23477 17660 23489 17663
rect 23440 17632 23489 17660
rect 23440 17620 23446 17632
rect 23477 17629 23489 17632
rect 23523 17629 23535 17663
rect 24848 17660 24860 17669
rect 24815 17632 24860 17660
rect 23477 17623 23535 17629
rect 24848 17623 24860 17632
rect 24854 17620 24860 17623
rect 24912 17620 24918 17672
rect 19521 17595 19579 17601
rect 19521 17592 19533 17595
rect 17368 17564 18276 17592
rect 18800 17564 19533 17592
rect 17368 17552 17374 17564
rect 15749 17527 15807 17533
rect 15749 17493 15761 17527
rect 15795 17524 15807 17527
rect 17954 17524 17960 17536
rect 15795 17496 17960 17524
rect 15795 17493 15807 17496
rect 15749 17487 15807 17493
rect 17954 17484 17960 17496
rect 18012 17484 18018 17536
rect 18248 17533 18276 17564
rect 19521 17561 19533 17564
rect 19567 17561 19579 17595
rect 19521 17555 19579 17561
rect 19705 17595 19763 17601
rect 19705 17561 19717 17595
rect 19751 17592 19763 17595
rect 21450 17592 21456 17604
rect 19751 17564 21456 17592
rect 19751 17561 19763 17564
rect 19705 17555 19763 17561
rect 21450 17552 21456 17564
rect 21508 17552 21514 17604
rect 28166 17592 28172 17604
rect 28127 17564 28172 17592
rect 28166 17552 28172 17564
rect 28224 17552 28230 17604
rect 18233 17527 18291 17533
rect 18233 17493 18245 17527
rect 18279 17493 18291 17527
rect 18414 17524 18420 17536
rect 18375 17496 18420 17524
rect 18233 17487 18291 17493
rect 18414 17484 18420 17496
rect 18472 17484 18478 17536
rect 22278 17484 22284 17536
rect 22336 17524 22342 17536
rect 22465 17527 22523 17533
rect 22465 17524 22477 17527
rect 22336 17496 22477 17524
rect 22336 17484 22342 17496
rect 22465 17493 22477 17496
rect 22511 17524 22523 17527
rect 24118 17524 24124 17536
rect 22511 17496 24124 17524
rect 22511 17493 22523 17496
rect 22465 17487 22523 17493
rect 24118 17484 24124 17496
rect 24176 17484 24182 17536
rect 25038 17484 25044 17536
rect 25096 17524 25102 17536
rect 25961 17527 26019 17533
rect 25961 17524 25973 17527
rect 25096 17496 25973 17524
rect 25096 17484 25102 17496
rect 25961 17493 25973 17496
rect 26007 17493 26019 17527
rect 25961 17487 26019 17493
rect 1104 17434 29048 17456
rect 1104 17382 7896 17434
rect 7948 17382 7960 17434
rect 8012 17382 8024 17434
rect 8076 17382 8088 17434
rect 8140 17382 8152 17434
rect 8204 17382 14842 17434
rect 14894 17382 14906 17434
rect 14958 17382 14970 17434
rect 15022 17382 15034 17434
rect 15086 17382 15098 17434
rect 15150 17382 21788 17434
rect 21840 17382 21852 17434
rect 21904 17382 21916 17434
rect 21968 17382 21980 17434
rect 22032 17382 22044 17434
rect 22096 17382 28734 17434
rect 28786 17382 28798 17434
rect 28850 17382 28862 17434
rect 28914 17382 28926 17434
rect 28978 17382 28990 17434
rect 29042 17382 29048 17434
rect 1104 17360 29048 17382
rect 1946 17320 1952 17332
rect 1907 17292 1952 17320
rect 1946 17280 1952 17292
rect 2004 17280 2010 17332
rect 17957 17323 18015 17329
rect 17957 17289 17969 17323
rect 18003 17320 18015 17323
rect 18414 17320 18420 17332
rect 18003 17292 18420 17320
rect 18003 17289 18015 17292
rect 17957 17283 18015 17289
rect 18414 17280 18420 17292
rect 18472 17280 18478 17332
rect 19886 17320 19892 17332
rect 19847 17292 19892 17320
rect 19886 17280 19892 17292
rect 19944 17280 19950 17332
rect 24670 17320 24676 17332
rect 22066 17292 24676 17320
rect 15470 17212 15476 17264
rect 15528 17252 15534 17264
rect 16025 17255 16083 17261
rect 16025 17252 16037 17255
rect 15528 17224 16037 17252
rect 15528 17212 15534 17224
rect 16025 17221 16037 17224
rect 16071 17252 16083 17255
rect 17310 17252 17316 17264
rect 16071 17224 17316 17252
rect 16071 17221 16083 17224
rect 16025 17215 16083 17221
rect 17310 17212 17316 17224
rect 17368 17212 17374 17264
rect 19058 17252 19064 17264
rect 18708 17224 19064 17252
rect 2038 17184 2044 17196
rect 1999 17156 2044 17184
rect 2038 17144 2044 17156
rect 2096 17144 2102 17196
rect 15749 17187 15807 17193
rect 15749 17153 15761 17187
rect 15795 17184 15807 17187
rect 15838 17184 15844 17196
rect 15795 17156 15844 17184
rect 15795 17153 15807 17156
rect 15749 17147 15807 17153
rect 15838 17144 15844 17156
rect 15896 17144 15902 17196
rect 16850 17184 16856 17196
rect 16811 17156 16856 17184
rect 16850 17144 16856 17156
rect 16908 17144 16914 17196
rect 17773 17187 17831 17193
rect 17773 17153 17785 17187
rect 17819 17184 17831 17187
rect 17862 17184 17868 17196
rect 17819 17156 17868 17184
rect 17819 17153 17831 17156
rect 17773 17147 17831 17153
rect 17862 17144 17868 17156
rect 17920 17144 17926 17196
rect 18708 17193 18736 17224
rect 19058 17212 19064 17224
rect 19116 17212 19122 17264
rect 22066 17252 22094 17292
rect 24670 17280 24676 17292
rect 24728 17280 24734 17332
rect 27157 17323 27215 17329
rect 27157 17289 27169 17323
rect 27203 17320 27215 17323
rect 27338 17320 27344 17332
rect 27203 17292 27344 17320
rect 27203 17289 27215 17292
rect 27157 17283 27215 17289
rect 27338 17280 27344 17292
rect 27396 17280 27402 17332
rect 27522 17320 27528 17332
rect 27483 17292 27528 17320
rect 27522 17280 27528 17292
rect 27580 17280 27586 17332
rect 22020 17224 22094 17252
rect 17957 17187 18015 17193
rect 17957 17153 17969 17187
rect 18003 17184 18015 17187
rect 18693 17187 18751 17193
rect 18693 17184 18705 17187
rect 18003 17156 18705 17184
rect 18003 17153 18015 17156
rect 17957 17147 18015 17153
rect 18693 17153 18705 17156
rect 18739 17153 18751 17187
rect 18693 17147 18751 17153
rect 18782 17144 18788 17196
rect 18840 17184 18846 17196
rect 18969 17187 19027 17193
rect 18969 17184 18981 17187
rect 18840 17156 18981 17184
rect 18840 17144 18846 17156
rect 18969 17153 18981 17156
rect 19015 17184 19027 17187
rect 19521 17187 19579 17193
rect 19521 17184 19533 17187
rect 19015 17156 19533 17184
rect 19015 17153 19027 17156
rect 18969 17147 19027 17153
rect 19521 17153 19533 17156
rect 19567 17153 19579 17187
rect 19521 17147 19579 17153
rect 19610 17144 19616 17196
rect 19668 17184 19674 17196
rect 22020 17193 22048 17224
rect 23934 17212 23940 17264
rect 23992 17252 23998 17264
rect 25501 17255 25559 17261
rect 25501 17252 25513 17255
rect 23992 17224 25513 17252
rect 23992 17212 23998 17224
rect 25501 17221 25513 17224
rect 25547 17221 25559 17255
rect 25501 17215 25559 17221
rect 19705 17187 19763 17193
rect 19705 17184 19717 17187
rect 19668 17156 19717 17184
rect 19668 17144 19674 17156
rect 19705 17153 19717 17156
rect 19751 17153 19763 17187
rect 19705 17147 19763 17153
rect 22005 17187 22063 17193
rect 22005 17153 22017 17187
rect 22051 17153 22063 17187
rect 22186 17184 22192 17196
rect 22147 17156 22192 17184
rect 22005 17147 22063 17153
rect 22186 17144 22192 17156
rect 22244 17144 22250 17196
rect 22373 17187 22431 17193
rect 22373 17153 22385 17187
rect 22419 17184 22431 17187
rect 22833 17187 22891 17193
rect 22833 17184 22845 17187
rect 22419 17156 22845 17184
rect 22419 17153 22431 17156
rect 22373 17147 22431 17153
rect 22833 17153 22845 17156
rect 22879 17153 22891 17187
rect 22833 17147 22891 17153
rect 23474 17144 23480 17196
rect 23532 17184 23538 17196
rect 23569 17187 23627 17193
rect 23569 17184 23581 17187
rect 23532 17156 23581 17184
rect 23532 17144 23538 17156
rect 23569 17153 23581 17156
rect 23615 17153 23627 17187
rect 23569 17147 23627 17153
rect 23658 17144 23664 17196
rect 23716 17184 23722 17196
rect 23825 17187 23883 17193
rect 23825 17184 23837 17187
rect 23716 17156 23837 17184
rect 23716 17144 23722 17156
rect 23825 17153 23837 17156
rect 23871 17153 23883 17187
rect 23825 17147 23883 17153
rect 25869 17187 25927 17193
rect 25869 17153 25881 17187
rect 25915 17184 25927 17187
rect 26418 17184 26424 17196
rect 25915 17156 26424 17184
rect 25915 17153 25927 17156
rect 25869 17147 25927 17153
rect 26418 17144 26424 17156
rect 26476 17144 26482 17196
rect 17880 17116 17908 17144
rect 18601 17119 18659 17125
rect 18601 17116 18613 17119
rect 17880 17088 18613 17116
rect 18601 17085 18613 17088
rect 18647 17085 18659 17119
rect 18601 17079 18659 17085
rect 19061 17119 19119 17125
rect 19061 17085 19073 17119
rect 19107 17085 19119 17119
rect 19334 17116 19340 17128
rect 19247 17088 19340 17116
rect 19061 17079 19119 17085
rect 18417 17051 18475 17057
rect 18417 17017 18429 17051
rect 18463 17048 18475 17051
rect 18690 17048 18696 17060
rect 18463 17020 18696 17048
rect 18463 17017 18475 17020
rect 18417 17011 18475 17017
rect 18690 17008 18696 17020
rect 18748 17008 18754 17060
rect 19076 17048 19104 17079
rect 19306 17076 19340 17088
rect 19392 17116 19398 17128
rect 19628 17116 19656 17144
rect 27614 17116 27620 17128
rect 19392 17088 19656 17116
rect 27575 17088 27620 17116
rect 19392 17076 19398 17088
rect 27614 17076 27620 17088
rect 27672 17076 27678 17128
rect 27709 17119 27767 17125
rect 27709 17085 27721 17119
rect 27755 17085 27767 17119
rect 27709 17079 27767 17085
rect 19306 17048 19334 17076
rect 19076 17020 19334 17048
rect 25866 17008 25872 17060
rect 25924 17048 25930 17060
rect 27724 17048 27752 17079
rect 25924 17020 27752 17048
rect 25924 17008 25930 17020
rect 17037 16983 17095 16989
rect 17037 16949 17049 16983
rect 17083 16980 17095 16983
rect 17126 16980 17132 16992
rect 17083 16952 17132 16980
rect 17083 16949 17095 16952
rect 17037 16943 17095 16949
rect 17126 16940 17132 16952
rect 17184 16940 17190 16992
rect 17310 16940 17316 16992
rect 17368 16980 17374 16992
rect 17862 16980 17868 16992
rect 17368 16952 17868 16980
rect 17368 16940 17374 16952
rect 17862 16940 17868 16952
rect 17920 16940 17926 16992
rect 23014 16980 23020 16992
rect 22975 16952 23020 16980
rect 23014 16940 23020 16952
rect 23072 16940 23078 16992
rect 24946 16980 24952 16992
rect 24907 16952 24952 16980
rect 24946 16940 24952 16952
rect 25004 16940 25010 16992
rect 26510 16980 26516 16992
rect 26471 16952 26516 16980
rect 26510 16940 26516 16952
rect 26568 16940 26574 16992
rect 1104 16890 28888 16912
rect 1104 16838 4423 16890
rect 4475 16838 4487 16890
rect 4539 16838 4551 16890
rect 4603 16838 4615 16890
rect 4667 16838 4679 16890
rect 4731 16838 11369 16890
rect 11421 16838 11433 16890
rect 11485 16838 11497 16890
rect 11549 16838 11561 16890
rect 11613 16838 11625 16890
rect 11677 16838 18315 16890
rect 18367 16838 18379 16890
rect 18431 16838 18443 16890
rect 18495 16838 18507 16890
rect 18559 16838 18571 16890
rect 18623 16838 25261 16890
rect 25313 16838 25325 16890
rect 25377 16838 25389 16890
rect 25441 16838 25453 16890
rect 25505 16838 25517 16890
rect 25569 16838 28888 16890
rect 1104 16816 28888 16838
rect 13262 16776 13268 16788
rect 13223 16748 13268 16776
rect 13262 16736 13268 16748
rect 13320 16736 13326 16788
rect 18230 16776 18236 16788
rect 16868 16748 18236 16776
rect 2222 16640 2228 16652
rect 2148 16612 2228 16640
rect 2148 16581 2176 16612
rect 2222 16600 2228 16612
rect 2280 16600 2286 16652
rect 16868 16649 16896 16748
rect 18230 16736 18236 16748
rect 18288 16736 18294 16788
rect 18782 16776 18788 16788
rect 18743 16748 18788 16776
rect 18782 16736 18788 16748
rect 18840 16736 18846 16788
rect 25866 16776 25872 16788
rect 22066 16748 25872 16776
rect 17862 16668 17868 16720
rect 17920 16708 17926 16720
rect 22066 16708 22094 16748
rect 25866 16736 25872 16748
rect 25924 16736 25930 16788
rect 26418 16736 26424 16788
rect 26476 16776 26482 16788
rect 27157 16779 27215 16785
rect 27157 16776 27169 16779
rect 26476 16748 27169 16776
rect 26476 16736 26482 16748
rect 27157 16745 27169 16748
rect 27203 16745 27215 16779
rect 27157 16739 27215 16745
rect 27893 16779 27951 16785
rect 27893 16745 27905 16779
rect 27939 16776 27951 16779
rect 28166 16776 28172 16788
rect 27939 16748 28172 16776
rect 27939 16745 27951 16748
rect 27893 16739 27951 16745
rect 28166 16736 28172 16748
rect 28224 16736 28230 16788
rect 17920 16680 22094 16708
rect 17920 16668 17926 16680
rect 16853 16643 16911 16649
rect 16853 16609 16865 16643
rect 16899 16609 16911 16643
rect 20438 16640 20444 16652
rect 16853 16603 16911 16609
rect 18892 16612 20444 16640
rect 2133 16575 2191 16581
rect 2133 16541 2145 16575
rect 2179 16541 2191 16575
rect 13446 16572 13452 16584
rect 13407 16544 13452 16572
rect 2133 16535 2191 16541
rect 13446 16532 13452 16544
rect 13504 16532 13510 16584
rect 13722 16572 13728 16584
rect 13683 16544 13728 16572
rect 13722 16532 13728 16544
rect 13780 16532 13786 16584
rect 17126 16581 17132 16584
rect 17120 16572 17132 16581
rect 17087 16544 17132 16572
rect 17120 16535 17132 16544
rect 17126 16532 17132 16535
rect 17184 16532 17190 16584
rect 18892 16581 18920 16612
rect 20438 16600 20444 16612
rect 20496 16600 20502 16652
rect 21266 16640 21272 16652
rect 21227 16612 21272 16640
rect 21266 16600 21272 16612
rect 21324 16600 21330 16652
rect 23293 16643 23351 16649
rect 23293 16609 23305 16643
rect 23339 16640 23351 16643
rect 23474 16640 23480 16652
rect 23339 16612 23480 16640
rect 23339 16609 23351 16612
rect 23293 16603 23351 16609
rect 23474 16600 23480 16612
rect 23532 16600 23538 16652
rect 24026 16640 24032 16652
rect 23952 16612 24032 16640
rect 18877 16575 18935 16581
rect 18877 16541 18889 16575
rect 18923 16541 18935 16575
rect 18877 16535 18935 16541
rect 18966 16532 18972 16584
rect 19024 16572 19030 16584
rect 19705 16575 19763 16581
rect 19705 16572 19717 16575
rect 19024 16544 19717 16572
rect 19024 16532 19030 16544
rect 19705 16541 19717 16544
rect 19751 16541 19763 16575
rect 19705 16535 19763 16541
rect 16022 16464 16028 16516
rect 16080 16504 16086 16516
rect 19720 16504 19748 16535
rect 20806 16532 20812 16584
rect 20864 16572 20870 16584
rect 21361 16575 21419 16581
rect 21361 16572 21373 16575
rect 20864 16544 21373 16572
rect 20864 16532 20870 16544
rect 21361 16541 21373 16544
rect 21407 16541 21419 16575
rect 21361 16535 21419 16541
rect 23014 16532 23020 16584
rect 23072 16581 23078 16584
rect 23072 16572 23084 16581
rect 23750 16572 23756 16584
rect 23072 16544 23117 16572
rect 23711 16544 23756 16572
rect 23072 16535 23084 16544
rect 23072 16532 23078 16535
rect 23750 16532 23756 16544
rect 23808 16532 23814 16584
rect 23952 16581 23980 16612
rect 24026 16600 24032 16612
rect 24084 16600 24090 16652
rect 25777 16643 25835 16649
rect 25777 16640 25789 16643
rect 24872 16612 25789 16640
rect 24872 16581 24900 16612
rect 25777 16609 25789 16612
rect 25823 16640 25835 16643
rect 26510 16640 26516 16652
rect 25823 16612 26516 16640
rect 25823 16609 25835 16612
rect 25777 16603 25835 16609
rect 26510 16600 26516 16612
rect 26568 16600 26574 16652
rect 27890 16640 27896 16652
rect 27816 16612 27896 16640
rect 23937 16575 23995 16581
rect 23937 16541 23949 16575
rect 23983 16541 23995 16575
rect 24857 16575 24915 16581
rect 24857 16572 24869 16575
rect 23937 16535 23995 16541
rect 24596 16544 24869 16572
rect 23842 16504 23848 16516
rect 16080 16476 19656 16504
rect 19720 16476 23704 16504
rect 23803 16476 23848 16504
rect 16080 16464 16086 16476
rect 1854 16396 1860 16448
rect 1912 16436 1918 16448
rect 2041 16439 2099 16445
rect 2041 16436 2053 16439
rect 1912 16408 2053 16436
rect 1912 16396 1918 16408
rect 2041 16405 2053 16408
rect 2087 16405 2099 16439
rect 2041 16399 2099 16405
rect 13633 16439 13691 16445
rect 13633 16405 13645 16439
rect 13679 16436 13691 16439
rect 13814 16436 13820 16448
rect 13679 16408 13820 16436
rect 13679 16405 13691 16408
rect 13633 16399 13691 16405
rect 13814 16396 13820 16408
rect 13872 16396 13878 16448
rect 17954 16396 17960 16448
rect 18012 16436 18018 16448
rect 18233 16439 18291 16445
rect 18233 16436 18245 16439
rect 18012 16408 18245 16436
rect 18012 16396 18018 16408
rect 18233 16405 18245 16408
rect 18279 16405 18291 16439
rect 18233 16399 18291 16405
rect 19426 16396 19432 16448
rect 19484 16436 19490 16448
rect 19521 16439 19579 16445
rect 19521 16436 19533 16439
rect 19484 16408 19533 16436
rect 19484 16396 19490 16408
rect 19521 16405 19533 16408
rect 19567 16405 19579 16439
rect 19628 16436 19656 16476
rect 20791 16439 20849 16445
rect 20791 16436 20803 16439
rect 19628 16408 20803 16436
rect 19521 16399 19579 16405
rect 20791 16405 20803 16408
rect 20837 16405 20849 16439
rect 20791 16399 20849 16405
rect 21269 16439 21327 16445
rect 21269 16405 21281 16439
rect 21315 16436 21327 16439
rect 21913 16439 21971 16445
rect 21913 16436 21925 16439
rect 21315 16408 21925 16436
rect 21315 16405 21327 16408
rect 21269 16399 21327 16405
rect 21913 16405 21925 16408
rect 21959 16436 21971 16439
rect 22370 16436 22376 16448
rect 21959 16408 22376 16436
rect 21959 16405 21971 16408
rect 21913 16399 21971 16405
rect 22370 16396 22376 16408
rect 22428 16396 22434 16448
rect 23676 16436 23704 16476
rect 23842 16464 23848 16476
rect 23900 16464 23906 16516
rect 24596 16436 24624 16544
rect 24857 16541 24869 16544
rect 24903 16541 24915 16575
rect 25590 16572 25596 16584
rect 25551 16544 25596 16572
rect 24857 16535 24915 16541
rect 25590 16532 25596 16544
rect 25648 16532 25654 16584
rect 27338 16572 27344 16584
rect 27299 16544 27344 16572
rect 27338 16532 27344 16544
rect 27396 16532 27402 16584
rect 27816 16581 27844 16612
rect 27890 16600 27896 16612
rect 27948 16600 27954 16652
rect 27801 16575 27859 16581
rect 27801 16541 27813 16575
rect 27847 16541 27859 16575
rect 27801 16535 27859 16541
rect 23676 16408 24624 16436
rect 24670 16396 24676 16448
rect 24728 16436 24734 16448
rect 24728 16408 24773 16436
rect 24728 16396 24734 16408
rect 24854 16396 24860 16448
rect 24912 16436 24918 16448
rect 25409 16439 25467 16445
rect 25409 16436 25421 16439
rect 24912 16408 25421 16436
rect 24912 16396 24918 16408
rect 25409 16405 25421 16408
rect 25455 16405 25467 16439
rect 25409 16399 25467 16405
rect 1104 16346 29048 16368
rect 1104 16294 7896 16346
rect 7948 16294 7960 16346
rect 8012 16294 8024 16346
rect 8076 16294 8088 16346
rect 8140 16294 8152 16346
rect 8204 16294 14842 16346
rect 14894 16294 14906 16346
rect 14958 16294 14970 16346
rect 15022 16294 15034 16346
rect 15086 16294 15098 16346
rect 15150 16294 21788 16346
rect 21840 16294 21852 16346
rect 21904 16294 21916 16346
rect 21968 16294 21980 16346
rect 22032 16294 22044 16346
rect 22096 16294 28734 16346
rect 28786 16294 28798 16346
rect 28850 16294 28862 16346
rect 28914 16294 28926 16346
rect 28978 16294 28990 16346
rect 29042 16294 29048 16346
rect 1104 16272 29048 16294
rect 13722 16192 13728 16244
rect 13780 16232 13786 16244
rect 14093 16235 14151 16241
rect 14093 16232 14105 16235
rect 13780 16204 14105 16232
rect 13780 16192 13786 16204
rect 14093 16201 14105 16204
rect 14139 16201 14151 16235
rect 20346 16232 20352 16244
rect 20307 16204 20352 16232
rect 14093 16195 14151 16201
rect 20346 16192 20352 16204
rect 20404 16192 20410 16244
rect 22005 16235 22063 16241
rect 22005 16201 22017 16235
rect 22051 16232 22063 16235
rect 22186 16232 22192 16244
rect 22051 16204 22192 16232
rect 22051 16201 22063 16204
rect 22005 16195 22063 16201
rect 22186 16192 22192 16204
rect 22244 16192 22250 16244
rect 22370 16232 22376 16244
rect 22331 16204 22376 16232
rect 22370 16192 22376 16204
rect 22428 16192 22434 16244
rect 24765 16235 24823 16241
rect 24765 16201 24777 16235
rect 24811 16201 24823 16235
rect 24765 16195 24823 16201
rect 1854 16164 1860 16176
rect 1815 16136 1860 16164
rect 1854 16124 1860 16136
rect 1912 16124 1918 16176
rect 14369 16167 14427 16173
rect 14369 16133 14381 16167
rect 14415 16164 14427 16167
rect 16022 16164 16028 16176
rect 14415 16136 16028 16164
rect 14415 16133 14427 16136
rect 14369 16127 14427 16133
rect 16022 16124 16028 16136
rect 16080 16124 16086 16176
rect 16117 16167 16175 16173
rect 16117 16133 16129 16167
rect 16163 16164 16175 16167
rect 24486 16164 24492 16176
rect 16163 16136 24492 16164
rect 16163 16133 16175 16136
rect 16117 16127 16175 16133
rect 24486 16124 24492 16136
rect 24544 16124 24550 16176
rect 24780 16164 24808 16195
rect 25470 16167 25528 16173
rect 25470 16164 25482 16167
rect 24780 16136 25482 16164
rect 25470 16133 25482 16136
rect 25516 16133 25528 16167
rect 25470 16127 25528 16133
rect 14093 16099 14151 16105
rect 14093 16065 14105 16099
rect 14139 16065 14151 16099
rect 14093 16059 14151 16065
rect 14185 16099 14243 16105
rect 14185 16065 14197 16099
rect 14231 16096 14243 16099
rect 14274 16096 14280 16108
rect 14231 16068 14280 16096
rect 14231 16065 14243 16068
rect 14185 16059 14243 16065
rect 1670 16028 1676 16040
rect 1631 16000 1676 16028
rect 1670 15988 1676 16000
rect 1728 15988 1734 16040
rect 2774 16028 2780 16040
rect 2735 16000 2780 16028
rect 2774 15988 2780 16000
rect 2832 15988 2838 16040
rect 14108 16028 14136 16059
rect 14274 16056 14280 16068
rect 14332 16056 14338 16108
rect 15194 16056 15200 16108
rect 15252 16096 15258 16108
rect 15749 16099 15807 16105
rect 15749 16096 15761 16099
rect 15252 16068 15761 16096
rect 15252 16056 15258 16068
rect 15749 16065 15761 16068
rect 15795 16065 15807 16099
rect 15749 16059 15807 16065
rect 15838 16056 15844 16108
rect 15896 16096 15902 16108
rect 15933 16099 15991 16105
rect 15933 16096 15945 16099
rect 15896 16068 15945 16096
rect 15896 16056 15902 16068
rect 15933 16065 15945 16068
rect 15979 16065 15991 16099
rect 15933 16059 15991 16065
rect 20441 16099 20499 16105
rect 20441 16065 20453 16099
rect 20487 16096 20499 16099
rect 20806 16096 20812 16108
rect 20487 16068 20812 16096
rect 20487 16065 20499 16068
rect 20441 16059 20499 16065
rect 20806 16056 20812 16068
rect 20864 16056 20870 16108
rect 24581 16099 24639 16105
rect 24581 16065 24593 16099
rect 24627 16096 24639 16099
rect 24854 16096 24860 16108
rect 24627 16068 24860 16096
rect 24627 16065 24639 16068
rect 24581 16059 24639 16065
rect 24854 16056 24860 16068
rect 24912 16056 24918 16108
rect 27154 16056 27160 16108
rect 27212 16096 27218 16108
rect 27433 16099 27491 16105
rect 27433 16096 27445 16099
rect 27212 16068 27445 16096
rect 27212 16056 27218 16068
rect 27433 16065 27445 16068
rect 27479 16065 27491 16099
rect 27433 16059 27491 16065
rect 20625 16031 20683 16037
rect 14108 16000 14688 16028
rect 14660 15904 14688 16000
rect 20625 15997 20637 16031
rect 20671 16028 20683 16031
rect 20714 16028 20720 16040
rect 20671 16000 20720 16028
rect 20671 15997 20683 16000
rect 20625 15991 20683 15997
rect 20714 15988 20720 16000
rect 20772 15988 20778 16040
rect 22465 16031 22523 16037
rect 22465 15997 22477 16031
rect 22511 15997 22523 16031
rect 22465 15991 22523 15997
rect 22480 15960 22508 15991
rect 22554 15988 22560 16040
rect 22612 16028 22618 16040
rect 22612 16000 22657 16028
rect 22612 15988 22618 16000
rect 23474 15988 23480 16040
rect 23532 16028 23538 16040
rect 23842 16028 23848 16040
rect 23532 16000 23848 16028
rect 23532 15988 23538 16000
rect 23842 15988 23848 16000
rect 23900 16028 23906 16040
rect 25225 16031 25283 16037
rect 25225 16028 25237 16031
rect 23900 16000 25237 16028
rect 23900 15988 23906 16000
rect 25225 15997 25237 16000
rect 25271 15997 25283 16031
rect 25225 15991 25283 15997
rect 22830 15960 22836 15972
rect 22480 15932 22836 15960
rect 22830 15920 22836 15932
rect 22888 15920 22894 15972
rect 14642 15852 14648 15904
rect 14700 15892 14706 15904
rect 16298 15892 16304 15904
rect 14700 15864 16304 15892
rect 14700 15852 14706 15864
rect 16298 15852 16304 15864
rect 16356 15892 16362 15904
rect 19981 15895 20039 15901
rect 19981 15892 19993 15895
rect 16356 15864 19993 15892
rect 16356 15852 16362 15864
rect 19981 15861 19993 15864
rect 20027 15861 20039 15895
rect 26602 15892 26608 15904
rect 26563 15864 26608 15892
rect 19981 15855 20039 15861
rect 26602 15852 26608 15864
rect 26660 15852 26666 15904
rect 27525 15895 27583 15901
rect 27525 15861 27537 15895
rect 27571 15892 27583 15895
rect 28166 15892 28172 15904
rect 27571 15864 28172 15892
rect 27571 15861 27583 15864
rect 27525 15855 27583 15861
rect 28166 15852 28172 15864
rect 28224 15852 28230 15904
rect 28261 15895 28319 15901
rect 28261 15861 28273 15895
rect 28307 15892 28319 15895
rect 28350 15892 28356 15904
rect 28307 15864 28356 15892
rect 28307 15861 28319 15864
rect 28261 15855 28319 15861
rect 28350 15852 28356 15864
rect 28408 15852 28414 15904
rect 1104 15802 28888 15824
rect 1104 15750 4423 15802
rect 4475 15750 4487 15802
rect 4539 15750 4551 15802
rect 4603 15750 4615 15802
rect 4667 15750 4679 15802
rect 4731 15750 11369 15802
rect 11421 15750 11433 15802
rect 11485 15750 11497 15802
rect 11549 15750 11561 15802
rect 11613 15750 11625 15802
rect 11677 15750 18315 15802
rect 18367 15750 18379 15802
rect 18431 15750 18443 15802
rect 18495 15750 18507 15802
rect 18559 15750 18571 15802
rect 18623 15750 25261 15802
rect 25313 15750 25325 15802
rect 25377 15750 25389 15802
rect 25441 15750 25453 15802
rect 25505 15750 25517 15802
rect 25569 15750 28888 15802
rect 1104 15728 28888 15750
rect 1670 15688 1676 15700
rect 1631 15660 1676 15688
rect 1670 15648 1676 15660
rect 1728 15648 1734 15700
rect 13725 15691 13783 15697
rect 13725 15657 13737 15691
rect 13771 15688 13783 15691
rect 13814 15688 13820 15700
rect 13771 15660 13820 15688
rect 13771 15657 13783 15660
rect 13725 15651 13783 15657
rect 13814 15648 13820 15660
rect 13872 15648 13878 15700
rect 15746 15688 15752 15700
rect 15707 15660 15752 15688
rect 15746 15648 15752 15660
rect 15804 15648 15810 15700
rect 20438 15648 20444 15700
rect 20496 15688 20502 15700
rect 25317 15691 25375 15697
rect 20496 15660 22094 15688
rect 20496 15648 20502 15660
rect 19610 15580 19616 15632
rect 19668 15620 19674 15632
rect 21361 15623 21419 15629
rect 21361 15620 21373 15623
rect 19668 15592 21373 15620
rect 19668 15580 19674 15592
rect 21361 15589 21373 15592
rect 21407 15589 21419 15623
rect 21361 15583 21419 15589
rect 20625 15555 20683 15561
rect 14476 15524 16160 15552
rect 12894 15444 12900 15496
rect 12952 15484 12958 15496
rect 13541 15487 13599 15493
rect 13541 15484 13553 15487
rect 12952 15456 13553 15484
rect 12952 15444 12958 15456
rect 13541 15453 13553 15456
rect 13587 15453 13599 15487
rect 13722 15484 13728 15496
rect 13683 15456 13728 15484
rect 13541 15447 13599 15453
rect 13556 15416 13584 15447
rect 13722 15444 13728 15456
rect 13780 15444 13786 15496
rect 14366 15444 14372 15496
rect 14424 15484 14430 15496
rect 14476 15493 14504 15524
rect 14461 15487 14519 15493
rect 14461 15484 14473 15487
rect 14424 15456 14473 15484
rect 14424 15444 14430 15456
rect 14461 15453 14473 15456
rect 14507 15453 14519 15487
rect 14642 15484 14648 15496
rect 14603 15456 14648 15484
rect 14461 15447 14519 15453
rect 14642 15444 14648 15456
rect 14700 15444 14706 15496
rect 15286 15444 15292 15496
rect 15344 15484 15350 15496
rect 16025 15487 16083 15493
rect 16025 15484 16037 15487
rect 15344 15456 16037 15484
rect 15344 15444 15350 15456
rect 16025 15453 16037 15456
rect 16071 15453 16083 15487
rect 16025 15447 16083 15453
rect 14553 15419 14611 15425
rect 14553 15416 14565 15419
rect 13556 15388 14565 15416
rect 14553 15385 14565 15388
rect 14599 15385 14611 15419
rect 14553 15379 14611 15385
rect 16132 15360 16160 15524
rect 20625 15521 20637 15555
rect 20671 15552 20683 15555
rect 20990 15552 20996 15564
rect 20671 15524 20996 15552
rect 20671 15521 20683 15524
rect 20625 15515 20683 15521
rect 20990 15512 20996 15524
rect 21048 15512 21054 15564
rect 20714 15484 20720 15496
rect 20675 15456 20720 15484
rect 20714 15444 20720 15456
rect 20772 15444 20778 15496
rect 21542 15444 21548 15496
rect 21600 15484 21606 15496
rect 21637 15487 21695 15493
rect 21637 15484 21649 15487
rect 21600 15456 21649 15484
rect 21600 15444 21606 15456
rect 21637 15453 21649 15456
rect 21683 15453 21695 15487
rect 22066 15484 22094 15660
rect 25317 15657 25329 15691
rect 25363 15688 25375 15691
rect 25590 15688 25596 15700
rect 25363 15660 25596 15688
rect 25363 15657 25375 15660
rect 25317 15651 25375 15657
rect 25590 15648 25596 15660
rect 25648 15648 25654 15700
rect 25866 15552 25872 15564
rect 25827 15524 25872 15552
rect 25866 15512 25872 15524
rect 25924 15512 25930 15564
rect 27522 15552 27528 15564
rect 27483 15524 27528 15552
rect 27522 15512 27528 15524
rect 27580 15512 27586 15564
rect 28166 15552 28172 15564
rect 28127 15524 28172 15552
rect 28166 15512 28172 15524
rect 28224 15512 28230 15564
rect 28350 15552 28356 15564
rect 28311 15524 28356 15552
rect 28350 15512 28356 15524
rect 28408 15512 28414 15564
rect 25685 15487 25743 15493
rect 25685 15484 25697 15487
rect 22066 15456 25697 15484
rect 21637 15447 21695 15453
rect 25685 15453 25697 15456
rect 25731 15484 25743 15487
rect 26602 15484 26608 15496
rect 25731 15456 26608 15484
rect 25731 15453 25743 15456
rect 25685 15447 25743 15453
rect 26602 15444 26608 15456
rect 26660 15444 26666 15496
rect 20732 15416 20760 15444
rect 21913 15419 21971 15425
rect 21913 15416 21925 15419
rect 20732 15388 21925 15416
rect 21913 15385 21925 15388
rect 21959 15385 21971 15419
rect 21913 15379 21971 15385
rect 15470 15308 15476 15360
rect 15528 15348 15534 15360
rect 15565 15351 15623 15357
rect 15565 15348 15577 15351
rect 15528 15320 15577 15348
rect 15528 15308 15534 15320
rect 15565 15317 15577 15320
rect 15611 15317 15623 15351
rect 15565 15311 15623 15317
rect 16114 15308 16120 15360
rect 16172 15348 16178 15360
rect 20147 15351 20205 15357
rect 20147 15348 20159 15351
rect 16172 15320 20159 15348
rect 16172 15308 16178 15320
rect 20147 15317 20159 15320
rect 20193 15317 20205 15351
rect 20147 15311 20205 15317
rect 20530 15308 20536 15360
rect 20588 15348 20594 15360
rect 20625 15351 20683 15357
rect 20625 15348 20637 15351
rect 20588 15320 20637 15348
rect 20588 15308 20594 15320
rect 20625 15317 20637 15320
rect 20671 15317 20683 15351
rect 20625 15311 20683 15317
rect 21821 15351 21879 15357
rect 21821 15317 21833 15351
rect 21867 15348 21879 15351
rect 22646 15348 22652 15360
rect 21867 15320 22652 15348
rect 21867 15317 21879 15320
rect 21821 15311 21879 15317
rect 22646 15308 22652 15320
rect 22704 15308 22710 15360
rect 25777 15351 25835 15357
rect 25777 15317 25789 15351
rect 25823 15348 25835 15351
rect 25866 15348 25872 15360
rect 25823 15320 25872 15348
rect 25823 15317 25835 15320
rect 25777 15311 25835 15317
rect 25866 15308 25872 15320
rect 25924 15308 25930 15360
rect 1104 15258 29048 15280
rect 1104 15206 7896 15258
rect 7948 15206 7960 15258
rect 8012 15206 8024 15258
rect 8076 15206 8088 15258
rect 8140 15206 8152 15258
rect 8204 15206 14842 15258
rect 14894 15206 14906 15258
rect 14958 15206 14970 15258
rect 15022 15206 15034 15258
rect 15086 15206 15098 15258
rect 15150 15206 21788 15258
rect 21840 15206 21852 15258
rect 21904 15206 21916 15258
rect 21968 15206 21980 15258
rect 22032 15206 22044 15258
rect 22096 15206 28734 15258
rect 28786 15206 28798 15258
rect 28850 15206 28862 15258
rect 28914 15206 28926 15258
rect 28978 15206 28990 15258
rect 29042 15206 29048 15258
rect 1104 15184 29048 15206
rect 13446 15104 13452 15156
rect 13504 15144 13510 15156
rect 13633 15147 13691 15153
rect 13633 15144 13645 15147
rect 13504 15116 13645 15144
rect 13504 15104 13510 15116
rect 13633 15113 13645 15116
rect 13679 15113 13691 15147
rect 14366 15144 14372 15156
rect 14327 15116 14372 15144
rect 13633 15107 13691 15113
rect 14366 15104 14372 15116
rect 14424 15104 14430 15156
rect 15013 15147 15071 15153
rect 15013 15113 15025 15147
rect 15059 15144 15071 15147
rect 15657 15147 15715 15153
rect 15657 15144 15669 15147
rect 15059 15116 15669 15144
rect 15059 15113 15071 15116
rect 15013 15107 15071 15113
rect 15657 15113 15669 15116
rect 15703 15144 15715 15147
rect 15746 15144 15752 15156
rect 15703 15116 15752 15144
rect 15703 15113 15715 15116
rect 15657 15107 15715 15113
rect 15746 15104 15752 15116
rect 15804 15104 15810 15156
rect 16298 15144 16304 15156
rect 16259 15116 16304 15144
rect 16298 15104 16304 15116
rect 16356 15104 16362 15156
rect 13722 15036 13728 15088
rect 13780 15076 13786 15088
rect 19610 15076 19616 15088
rect 13780 15048 15240 15076
rect 13780 15036 13786 15048
rect 2038 15008 2044 15020
rect 1951 14980 2044 15008
rect 2038 14968 2044 14980
rect 2096 15008 2102 15020
rect 2498 15008 2504 15020
rect 2096 14980 2504 15008
rect 2096 14968 2102 14980
rect 2498 14968 2504 14980
rect 2556 14968 2562 15020
rect 13354 14968 13360 15020
rect 13412 15008 13418 15020
rect 13449 15011 13507 15017
rect 13449 15008 13461 15011
rect 13412 14980 13461 15008
rect 13412 14968 13418 14980
rect 13449 14977 13461 14980
rect 13495 15008 13507 15011
rect 13740 15008 13768 15036
rect 13495 14980 13768 15008
rect 14185 15011 14243 15017
rect 13495 14977 13507 14980
rect 13449 14971 13507 14977
rect 14185 14977 14197 15011
rect 14231 14977 14243 15011
rect 14185 14971 14243 14977
rect 12894 14900 12900 14952
rect 12952 14940 12958 14952
rect 13265 14943 13323 14949
rect 13265 14940 13277 14943
rect 12952 14912 13277 14940
rect 12952 14900 12958 14912
rect 13265 14909 13277 14912
rect 13311 14940 13323 14943
rect 14200 14940 14228 14971
rect 14274 14968 14280 15020
rect 14332 15008 14338 15020
rect 15212 15017 15240 15048
rect 17052 15048 19616 15076
rect 17052 15017 17080 15048
rect 19610 15036 19616 15048
rect 19668 15036 19674 15088
rect 19334 15017 19340 15020
rect 14461 15011 14519 15017
rect 14461 15008 14473 15011
rect 14332 14980 14473 15008
rect 14332 14968 14338 14980
rect 14461 14977 14473 14980
rect 14507 14977 14519 15011
rect 14461 14971 14519 14977
rect 14921 15011 14979 15017
rect 14921 14977 14933 15011
rect 14967 14977 14979 15011
rect 14921 14971 14979 14977
rect 15197 15011 15255 15017
rect 15197 14977 15209 15011
rect 15243 15008 15255 15011
rect 17037 15011 17095 15017
rect 17037 15008 17049 15011
rect 15243 14980 17049 15008
rect 15243 14977 15255 14980
rect 15197 14971 15255 14977
rect 17037 14977 17049 14980
rect 17083 14977 17095 15011
rect 17037 14971 17095 14977
rect 19328 14971 19340 15017
rect 19392 15008 19398 15020
rect 19392 14980 19428 15008
rect 13311 14912 14228 14940
rect 13311 14909 13323 14912
rect 13265 14903 13323 14909
rect 12618 14832 12624 14884
rect 12676 14872 12682 14884
rect 14642 14872 14648 14884
rect 12676 14844 14648 14872
rect 12676 14832 12682 14844
rect 14642 14832 14648 14844
rect 14700 14832 14706 14884
rect 14936 14872 14964 14971
rect 19334 14968 19340 14971
rect 19392 14968 19398 14980
rect 23106 14968 23112 15020
rect 23164 15008 23170 15020
rect 23578 15011 23636 15017
rect 23578 15008 23590 15011
rect 23164 14980 23590 15008
rect 23164 14968 23170 14980
rect 23578 14977 23590 14980
rect 23624 14977 23636 15011
rect 23842 15008 23848 15020
rect 23803 14980 23848 15008
rect 23578 14971 23636 14977
rect 23842 14968 23848 14980
rect 23900 14968 23906 15020
rect 26878 14968 26884 15020
rect 26936 15008 26942 15020
rect 27433 15011 27491 15017
rect 27433 15008 27445 15011
rect 26936 14980 27445 15008
rect 26936 14968 26942 14980
rect 27433 14977 27445 14980
rect 27479 15008 27491 15011
rect 27522 15008 27528 15020
rect 27479 14980 27528 15008
rect 27479 14977 27491 14980
rect 27433 14971 27491 14977
rect 27522 14968 27528 14980
rect 27580 14968 27586 15020
rect 15841 14943 15899 14949
rect 15841 14909 15853 14943
rect 15887 14909 15899 14943
rect 15841 14903 15899 14909
rect 15933 14943 15991 14949
rect 15933 14909 15945 14943
rect 15979 14940 15991 14943
rect 16114 14940 16120 14952
rect 15979 14912 16120 14940
rect 15979 14909 15991 14912
rect 15933 14903 15991 14909
rect 15194 14872 15200 14884
rect 14936 14844 15056 14872
rect 15155 14844 15200 14872
rect 1762 14764 1768 14816
rect 1820 14804 1826 14816
rect 1949 14807 2007 14813
rect 1949 14804 1961 14807
rect 1820 14776 1961 14804
rect 1820 14764 1826 14776
rect 1949 14773 1961 14776
rect 1995 14773 2007 14807
rect 1949 14767 2007 14773
rect 14185 14807 14243 14813
rect 14185 14773 14197 14807
rect 14231 14804 14243 14807
rect 14734 14804 14740 14816
rect 14231 14776 14740 14804
rect 14231 14773 14243 14776
rect 14185 14767 14243 14773
rect 14734 14764 14740 14776
rect 14792 14764 14798 14816
rect 15028 14804 15056 14844
rect 15194 14832 15200 14844
rect 15252 14832 15258 14884
rect 15856 14872 15884 14903
rect 16114 14900 16120 14912
rect 16172 14900 16178 14952
rect 19058 14940 19064 14952
rect 19019 14912 19064 14940
rect 19058 14900 19064 14912
rect 19116 14900 19122 14952
rect 16022 14872 16028 14884
rect 15856 14844 16028 14872
rect 16022 14832 16028 14844
rect 16080 14832 16086 14884
rect 15286 14804 15292 14816
rect 15028 14776 15292 14804
rect 15286 14764 15292 14776
rect 15344 14764 15350 14816
rect 15562 14764 15568 14816
rect 15620 14804 15626 14816
rect 16945 14807 17003 14813
rect 16945 14804 16957 14807
rect 15620 14776 16957 14804
rect 15620 14764 15626 14776
rect 16945 14773 16957 14776
rect 16991 14773 17003 14807
rect 20438 14804 20444 14816
rect 20399 14776 20444 14804
rect 16945 14767 17003 14773
rect 20438 14764 20444 14776
rect 20496 14764 20502 14816
rect 22370 14764 22376 14816
rect 22428 14804 22434 14816
rect 22465 14807 22523 14813
rect 22465 14804 22477 14807
rect 22428 14776 22477 14804
rect 22428 14764 22434 14776
rect 22465 14773 22477 14776
rect 22511 14773 22523 14807
rect 22465 14767 22523 14773
rect 26694 14764 26700 14816
rect 26752 14804 26758 14816
rect 27341 14807 27399 14813
rect 27341 14804 27353 14807
rect 26752 14776 27353 14804
rect 26752 14764 26758 14776
rect 27341 14773 27353 14776
rect 27387 14773 27399 14807
rect 27890 14804 27896 14816
rect 27851 14776 27896 14804
rect 27341 14767 27399 14773
rect 27890 14764 27896 14776
rect 27948 14764 27954 14816
rect 1104 14714 28888 14736
rect 1104 14662 4423 14714
rect 4475 14662 4487 14714
rect 4539 14662 4551 14714
rect 4603 14662 4615 14714
rect 4667 14662 4679 14714
rect 4731 14662 11369 14714
rect 11421 14662 11433 14714
rect 11485 14662 11497 14714
rect 11549 14662 11561 14714
rect 11613 14662 11625 14714
rect 11677 14662 18315 14714
rect 18367 14662 18379 14714
rect 18431 14662 18443 14714
rect 18495 14662 18507 14714
rect 18559 14662 18571 14714
rect 18623 14662 25261 14714
rect 25313 14662 25325 14714
rect 25377 14662 25389 14714
rect 25441 14662 25453 14714
rect 25505 14662 25517 14714
rect 25569 14662 28888 14714
rect 1104 14640 28888 14662
rect 14277 14603 14335 14609
rect 14277 14600 14289 14603
rect 11440 14572 14289 14600
rect 1762 14464 1768 14476
rect 1723 14436 1768 14464
rect 1762 14424 1768 14436
rect 1820 14424 1826 14476
rect 2774 14464 2780 14476
rect 2735 14436 2780 14464
rect 2774 14424 2780 14436
rect 2832 14424 2838 14476
rect 9674 14464 9680 14476
rect 9635 14436 9680 14464
rect 9674 14424 9680 14436
rect 9732 14424 9738 14476
rect 11440 14473 11468 14572
rect 14277 14569 14289 14572
rect 14323 14569 14335 14603
rect 14277 14563 14335 14569
rect 15933 14603 15991 14609
rect 15933 14569 15945 14603
rect 15979 14600 15991 14603
rect 20806 14600 20812 14612
rect 15979 14572 20392 14600
rect 20767 14572 20812 14600
rect 15979 14569 15991 14572
rect 15933 14563 15991 14569
rect 12437 14535 12495 14541
rect 12437 14501 12449 14535
rect 12483 14532 12495 14535
rect 12483 14504 13032 14532
rect 12483 14501 12495 14504
rect 12437 14495 12495 14501
rect 11425 14467 11483 14473
rect 11425 14433 11437 14467
rect 11471 14433 11483 14467
rect 12618 14464 12624 14476
rect 11425 14427 11483 14433
rect 12268 14436 12624 14464
rect 1578 14396 1584 14408
rect 1539 14368 1584 14396
rect 1578 14356 1584 14368
rect 1636 14356 1642 14408
rect 8386 14396 8392 14408
rect 8299 14368 8392 14396
rect 8386 14356 8392 14368
rect 8444 14356 8450 14408
rect 12268 14405 12296 14436
rect 12618 14424 12624 14436
rect 12676 14424 12682 14476
rect 12894 14464 12900 14476
rect 12855 14436 12900 14464
rect 12894 14424 12900 14436
rect 12952 14424 12958 14476
rect 13004 14464 13032 14504
rect 13078 14492 13084 14544
rect 13136 14532 13142 14544
rect 14826 14532 14832 14544
rect 13136 14504 14832 14532
rect 13136 14492 13142 14504
rect 14826 14492 14832 14504
rect 14884 14532 14890 14544
rect 16022 14532 16028 14544
rect 14884 14504 16028 14532
rect 14884 14492 14890 14504
rect 16022 14492 16028 14504
rect 16080 14492 16086 14544
rect 18046 14492 18052 14544
rect 18104 14532 18110 14544
rect 18233 14535 18291 14541
rect 18233 14532 18245 14535
rect 18104 14504 18245 14532
rect 18104 14492 18110 14504
rect 18233 14501 18245 14504
rect 18279 14501 18291 14535
rect 20364 14532 20392 14572
rect 20806 14560 20812 14572
rect 20864 14560 20870 14612
rect 26326 14600 26332 14612
rect 20916 14572 26332 14600
rect 20916 14532 20944 14572
rect 26326 14560 26332 14572
rect 26384 14560 26390 14612
rect 27890 14532 27896 14544
rect 20364 14504 20944 14532
rect 26528 14504 27896 14532
rect 18233 14495 18291 14501
rect 13004 14436 13124 14464
rect 12253 14399 12311 14405
rect 12253 14365 12265 14399
rect 12299 14365 12311 14399
rect 12253 14359 12311 14365
rect 12437 14399 12495 14405
rect 12437 14365 12449 14399
rect 12483 14365 12495 14399
rect 13096 14396 13124 14436
rect 14274 14424 14280 14476
rect 14332 14464 14338 14476
rect 14332 14436 15608 14464
rect 14332 14424 14338 14436
rect 13173 14399 13231 14405
rect 13173 14396 13185 14399
rect 13096 14368 13185 14396
rect 12437 14359 12495 14365
rect 13173 14365 13185 14368
rect 13219 14365 13231 14399
rect 13354 14396 13360 14408
rect 13315 14368 13360 14396
rect 13173 14359 13231 14365
rect 8404 14328 8432 14356
rect 10962 14328 10968 14340
rect 8404 14300 10968 14328
rect 10962 14288 10968 14300
rect 11020 14288 11026 14340
rect 11238 14328 11244 14340
rect 11199 14300 11244 14328
rect 11238 14288 11244 14300
rect 11296 14288 11302 14340
rect 12452 14328 12480 14359
rect 12894 14328 12900 14340
rect 12452 14300 12900 14328
rect 12894 14288 12900 14300
rect 12952 14288 12958 14340
rect 13188 14328 13216 14359
rect 13354 14356 13360 14368
rect 13412 14356 13418 14408
rect 14568 14405 14596 14436
rect 15580 14408 15608 14436
rect 18138 14424 18144 14476
rect 18196 14464 18202 14476
rect 18196 14436 18920 14464
rect 18196 14424 18202 14436
rect 14415 14399 14473 14405
rect 14415 14396 14427 14399
rect 13464 14368 14427 14396
rect 13464 14328 13492 14368
rect 14415 14365 14427 14368
rect 14461 14365 14473 14399
rect 14415 14359 14473 14365
rect 14553 14399 14611 14405
rect 14553 14365 14565 14399
rect 14599 14365 14611 14399
rect 14826 14396 14832 14408
rect 14787 14368 14832 14396
rect 14553 14359 14611 14365
rect 14826 14356 14832 14368
rect 14884 14356 14890 14408
rect 14921 14399 14979 14405
rect 14921 14365 14933 14399
rect 14967 14365 14979 14399
rect 15470 14396 15476 14408
rect 15431 14368 15476 14396
rect 14921 14359 14979 14365
rect 13188 14300 13492 14328
rect 13814 14288 13820 14340
rect 13872 14328 13878 14340
rect 14642 14328 14648 14340
rect 13872 14300 14648 14328
rect 13872 14288 13878 14300
rect 14642 14288 14648 14300
rect 14700 14288 14706 14340
rect 14936 14328 14964 14359
rect 15470 14356 15476 14368
rect 15528 14356 15534 14408
rect 15562 14356 15568 14408
rect 15620 14396 15626 14408
rect 15749 14399 15807 14405
rect 15620 14368 15665 14396
rect 15620 14356 15626 14368
rect 15749 14365 15761 14399
rect 15795 14396 15807 14399
rect 15838 14396 15844 14408
rect 15795 14368 15844 14396
rect 15795 14365 15807 14368
rect 15749 14359 15807 14365
rect 15764 14328 15792 14359
rect 15838 14356 15844 14368
rect 15896 14356 15902 14408
rect 16853 14399 16911 14405
rect 16853 14365 16865 14399
rect 16899 14396 16911 14399
rect 18230 14396 18236 14408
rect 16899 14368 18236 14396
rect 16899 14365 16911 14368
rect 16853 14359 16911 14365
rect 18230 14356 18236 14368
rect 18288 14356 18294 14408
rect 18892 14405 18920 14436
rect 23842 14424 23848 14476
rect 23900 14464 23906 14476
rect 24210 14464 24216 14476
rect 23900 14436 24216 14464
rect 23900 14424 23906 14436
rect 24210 14424 24216 14436
rect 24268 14464 24274 14476
rect 26528 14473 26556 14504
rect 27890 14492 27896 14504
rect 27948 14492 27954 14544
rect 24581 14467 24639 14473
rect 24581 14464 24593 14467
rect 24268 14436 24593 14464
rect 24268 14424 24274 14436
rect 24581 14433 24593 14436
rect 24627 14433 24639 14467
rect 24581 14427 24639 14433
rect 26513 14467 26571 14473
rect 26513 14433 26525 14467
rect 26559 14433 26571 14467
rect 26694 14464 26700 14476
rect 26655 14436 26700 14464
rect 26513 14427 26571 14433
rect 26694 14424 26700 14436
rect 26752 14424 26758 14476
rect 18877 14399 18935 14405
rect 18877 14365 18889 14399
rect 18923 14365 18935 14399
rect 18877 14359 18935 14365
rect 19058 14356 19064 14408
rect 19116 14396 19122 14408
rect 19429 14399 19487 14405
rect 19429 14396 19441 14399
rect 19116 14368 19441 14396
rect 19116 14356 19122 14368
rect 19429 14365 19441 14368
rect 19475 14396 19487 14399
rect 21266 14396 21272 14408
rect 19475 14368 21272 14396
rect 19475 14365 19487 14368
rect 19429 14359 19487 14365
rect 21266 14356 21272 14368
rect 21324 14356 21330 14408
rect 28350 14396 28356 14408
rect 28311 14368 28356 14396
rect 28350 14356 28356 14368
rect 28408 14356 28414 14408
rect 14936 14300 15792 14328
rect 8481 14263 8539 14269
rect 8481 14229 8493 14263
rect 8527 14260 8539 14263
rect 9950 14260 9956 14272
rect 8527 14232 9956 14260
rect 8527 14229 8539 14232
rect 8481 14223 8539 14229
rect 9950 14220 9956 14232
rect 10008 14220 10014 14272
rect 13078 14260 13084 14272
rect 13039 14232 13084 14260
rect 13078 14220 13084 14232
rect 13136 14220 13142 14272
rect 13446 14220 13452 14272
rect 13504 14260 13510 14272
rect 14936 14260 14964 14300
rect 16298 14288 16304 14340
rect 16356 14328 16362 14340
rect 19702 14337 19708 14340
rect 17098 14331 17156 14337
rect 17098 14328 17110 14331
rect 16356 14300 17110 14328
rect 16356 14288 16362 14300
rect 17098 14297 17110 14300
rect 17144 14297 17156 14331
rect 17098 14291 17156 14297
rect 19696 14291 19708 14337
rect 19760 14328 19766 14340
rect 21542 14337 21548 14340
rect 19760 14300 19796 14328
rect 19702 14288 19708 14291
rect 19760 14288 19766 14300
rect 21536 14291 21548 14337
rect 21600 14328 21606 14340
rect 21600 14300 21636 14328
rect 21542 14288 21548 14291
rect 21600 14288 21606 14300
rect 24578 14288 24584 14340
rect 24636 14328 24642 14340
rect 24826 14331 24884 14337
rect 24826 14328 24838 14331
rect 24636 14300 24838 14328
rect 24636 14288 24642 14300
rect 24826 14297 24838 14300
rect 24872 14297 24884 14331
rect 24826 14291 24884 14297
rect 13504 14232 14964 14260
rect 13504 14220 13510 14232
rect 18506 14220 18512 14272
rect 18564 14260 18570 14272
rect 18693 14263 18751 14269
rect 18693 14260 18705 14263
rect 18564 14232 18705 14260
rect 18564 14220 18570 14232
rect 18693 14229 18705 14232
rect 18739 14229 18751 14263
rect 22646 14260 22652 14272
rect 22607 14232 22652 14260
rect 18693 14223 18751 14229
rect 22646 14220 22652 14232
rect 22704 14220 22710 14272
rect 25958 14260 25964 14272
rect 25919 14232 25964 14260
rect 25958 14220 25964 14232
rect 26016 14220 26022 14272
rect 1104 14170 29048 14192
rect 1104 14118 7896 14170
rect 7948 14118 7960 14170
rect 8012 14118 8024 14170
rect 8076 14118 8088 14170
rect 8140 14118 8152 14170
rect 8204 14118 14842 14170
rect 14894 14118 14906 14170
rect 14958 14118 14970 14170
rect 15022 14118 15034 14170
rect 15086 14118 15098 14170
rect 15150 14118 21788 14170
rect 21840 14118 21852 14170
rect 21904 14118 21916 14170
rect 21968 14118 21980 14170
rect 22032 14118 22044 14170
rect 22096 14118 28734 14170
rect 28786 14118 28798 14170
rect 28850 14118 28862 14170
rect 28914 14118 28926 14170
rect 28978 14118 28990 14170
rect 29042 14118 29048 14170
rect 1104 14096 29048 14118
rect 13078 14056 13084 14068
rect 10152 14028 13084 14056
rect 9950 13988 9956 14000
rect 9911 13960 9956 13988
rect 9950 13948 9956 13960
rect 10008 13948 10014 14000
rect 1578 13880 1584 13932
rect 1636 13920 1642 13932
rect 1673 13923 1731 13929
rect 1673 13920 1685 13923
rect 1636 13892 1685 13920
rect 1636 13880 1642 13892
rect 1673 13889 1685 13892
rect 1719 13889 1731 13923
rect 1673 13883 1731 13889
rect 3694 13880 3700 13932
rect 3752 13920 3758 13932
rect 10152 13929 10180 14028
rect 13078 14016 13084 14028
rect 13136 14016 13142 14068
rect 15286 14056 15292 14068
rect 15247 14028 15292 14056
rect 15286 14016 15292 14028
rect 15344 14016 15350 14068
rect 16114 14056 16120 14068
rect 15488 14028 16120 14056
rect 11057 13991 11115 13997
rect 11057 13957 11069 13991
rect 11103 13988 11115 13991
rect 13357 13991 13415 13997
rect 13357 13988 13369 13991
rect 11103 13960 13369 13988
rect 11103 13957 11115 13960
rect 11057 13951 11115 13957
rect 13357 13957 13369 13960
rect 13403 13957 13415 13991
rect 15304 13988 15332 14016
rect 15488 13997 15516 14028
rect 16114 14016 16120 14028
rect 16172 14016 16178 14068
rect 16298 14056 16304 14068
rect 16259 14028 16304 14056
rect 16298 14016 16304 14028
rect 16356 14016 16362 14068
rect 17221 14059 17279 14065
rect 17221 14025 17233 14059
rect 17267 14056 17279 14059
rect 18046 14056 18052 14068
rect 17267 14028 18052 14056
rect 17267 14025 17279 14028
rect 17221 14019 17279 14025
rect 18046 14016 18052 14028
rect 18104 14016 18110 14068
rect 19518 14016 19524 14068
rect 19576 14056 19582 14068
rect 19613 14059 19671 14065
rect 19613 14056 19625 14059
rect 19576 14028 19625 14056
rect 19576 14016 19582 14028
rect 19613 14025 19625 14028
rect 19659 14025 19671 14059
rect 19613 14019 19671 14025
rect 27614 14016 27620 14068
rect 27672 14056 27678 14068
rect 28169 14059 28227 14065
rect 28169 14056 28181 14059
rect 27672 14028 28181 14056
rect 27672 14016 27678 14028
rect 28169 14025 28181 14028
rect 28215 14025 28227 14059
rect 28169 14019 28227 14025
rect 13357 13951 13415 13957
rect 14568 13960 15332 13988
rect 15473 13991 15531 13997
rect 10137 13923 10195 13929
rect 3752 13892 8800 13920
rect 3752 13880 3758 13892
rect 2501 13855 2559 13861
rect 2501 13821 2513 13855
rect 2547 13852 2559 13855
rect 3418 13852 3424 13864
rect 2547 13824 3424 13852
rect 2547 13821 2559 13824
rect 2501 13815 2559 13821
rect 3418 13812 3424 13824
rect 3476 13812 3482 13864
rect 8294 13852 8300 13864
rect 8255 13824 8300 13852
rect 8294 13812 8300 13824
rect 8352 13812 8358 13864
rect 8772 13852 8800 13892
rect 10137 13889 10149 13923
rect 10183 13889 10195 13923
rect 10962 13920 10968 13932
rect 10923 13892 10968 13920
rect 10137 13883 10195 13889
rect 10962 13880 10968 13892
rect 11020 13880 11026 13932
rect 11701 13855 11759 13861
rect 11701 13852 11713 13855
rect 8772 13824 11713 13852
rect 11701 13821 11713 13824
rect 11747 13821 11759 13855
rect 11701 13815 11759 13821
rect 13541 13855 13599 13861
rect 13541 13821 13553 13855
rect 13587 13852 13599 13855
rect 14277 13855 14335 13861
rect 14277 13852 14289 13855
rect 13587 13824 14289 13852
rect 13587 13821 13599 13824
rect 13541 13815 13599 13821
rect 14277 13821 14289 13824
rect 14323 13821 14335 13855
rect 14458 13852 14464 13864
rect 14419 13824 14464 13852
rect 14277 13815 14335 13821
rect 14458 13812 14464 13824
rect 14516 13812 14522 13864
rect 14568 13861 14596 13960
rect 15473 13957 15485 13991
rect 15519 13957 15531 13991
rect 15473 13951 15531 13957
rect 15657 13991 15715 13997
rect 15657 13957 15669 13991
rect 15703 13988 15715 13991
rect 16022 13988 16028 14000
rect 15703 13960 16028 13988
rect 15703 13957 15715 13960
rect 15657 13951 15715 13957
rect 14737 13923 14795 13929
rect 14737 13889 14749 13923
rect 14783 13920 14795 13923
rect 15010 13920 15016 13932
rect 14783 13892 15016 13920
rect 14783 13889 14795 13892
rect 14737 13883 14795 13889
rect 15010 13880 15016 13892
rect 15068 13880 15074 13932
rect 15102 13880 15108 13932
rect 15160 13920 15166 13932
rect 15672 13920 15700 13951
rect 16022 13948 16028 13960
rect 16080 13948 16086 14000
rect 19058 13988 19064 14000
rect 18340 13960 19064 13988
rect 15160 13892 15700 13920
rect 16117 13923 16175 13929
rect 15160 13880 15166 13892
rect 16117 13889 16129 13923
rect 16163 13920 16175 13923
rect 16574 13920 16580 13932
rect 16163 13892 16580 13920
rect 16163 13889 16175 13892
rect 16117 13883 16175 13889
rect 16574 13880 16580 13892
rect 16632 13880 16638 13932
rect 17313 13923 17371 13929
rect 17313 13889 17325 13923
rect 17359 13920 17371 13923
rect 17586 13920 17592 13932
rect 17359 13892 17592 13920
rect 17359 13889 17371 13892
rect 17313 13883 17371 13889
rect 17586 13880 17592 13892
rect 17644 13880 17650 13932
rect 18230 13920 18236 13932
rect 18143 13892 18236 13920
rect 18230 13880 18236 13892
rect 18288 13920 18294 13932
rect 18340 13920 18368 13960
rect 19058 13948 19064 13960
rect 19116 13948 19122 14000
rect 21634 13948 21640 14000
rect 21692 13988 21698 14000
rect 22250 13991 22308 13997
rect 22250 13988 22262 13991
rect 21692 13960 22262 13988
rect 21692 13948 21698 13960
rect 22250 13957 22262 13960
rect 22296 13957 22308 13991
rect 22250 13951 22308 13957
rect 18506 13929 18512 13932
rect 18500 13920 18512 13929
rect 18288 13892 18368 13920
rect 18467 13892 18512 13920
rect 18288 13880 18294 13892
rect 18500 13883 18512 13892
rect 18506 13880 18512 13883
rect 18564 13880 18570 13932
rect 21266 13880 21272 13932
rect 21324 13920 21330 13932
rect 22005 13923 22063 13929
rect 22005 13920 22017 13923
rect 21324 13892 22017 13920
rect 21324 13880 21330 13892
rect 22005 13889 22017 13892
rect 22051 13889 22063 13923
rect 24210 13920 24216 13932
rect 24171 13892 24216 13920
rect 22005 13883 22063 13889
rect 24210 13880 24216 13892
rect 24268 13880 24274 13932
rect 24480 13923 24538 13929
rect 24480 13889 24492 13923
rect 24526 13920 24538 13923
rect 24762 13920 24768 13932
rect 24526 13892 24768 13920
rect 24526 13889 24538 13892
rect 24480 13883 24538 13889
rect 24762 13880 24768 13892
rect 24820 13880 24826 13932
rect 27154 13880 27160 13932
rect 27212 13920 27218 13932
rect 27341 13923 27399 13929
rect 27341 13920 27353 13923
rect 27212 13892 27353 13920
rect 27212 13880 27218 13892
rect 27341 13889 27353 13892
rect 27387 13889 27399 13923
rect 27341 13883 27399 13889
rect 28353 13923 28411 13929
rect 28353 13889 28365 13923
rect 28399 13920 28411 13923
rect 28442 13920 28448 13932
rect 28399 13892 28448 13920
rect 28399 13889 28411 13892
rect 28353 13883 28411 13889
rect 28442 13880 28448 13892
rect 28500 13880 28506 13932
rect 14553 13855 14611 13861
rect 14553 13821 14565 13855
rect 14599 13821 14611 13855
rect 14553 13815 14611 13821
rect 14642 13812 14648 13864
rect 14700 13852 14706 13864
rect 17405 13855 17463 13861
rect 14700 13824 14745 13852
rect 14700 13812 14706 13824
rect 17405 13821 17417 13855
rect 17451 13821 17463 13855
rect 17405 13815 17463 13821
rect 17310 13744 17316 13796
rect 17368 13784 17374 13796
rect 17420 13784 17448 13815
rect 17368 13756 17448 13784
rect 17368 13744 17374 13756
rect 16758 13676 16764 13728
rect 16816 13716 16822 13728
rect 16853 13719 16911 13725
rect 16853 13716 16865 13719
rect 16816 13688 16865 13716
rect 16816 13676 16822 13688
rect 16853 13685 16865 13688
rect 16899 13685 16911 13719
rect 23382 13716 23388 13728
rect 23343 13688 23388 13716
rect 16853 13679 16911 13685
rect 23382 13676 23388 13688
rect 23440 13676 23446 13728
rect 25590 13716 25596 13728
rect 25551 13688 25596 13716
rect 25590 13676 25596 13688
rect 25648 13676 25654 13728
rect 26694 13676 26700 13728
rect 26752 13716 26758 13728
rect 27249 13719 27307 13725
rect 27249 13716 27261 13719
rect 26752 13688 27261 13716
rect 26752 13676 26758 13688
rect 27249 13685 27261 13688
rect 27295 13685 27307 13719
rect 27249 13679 27307 13685
rect 1104 13626 28888 13648
rect 1104 13574 4423 13626
rect 4475 13574 4487 13626
rect 4539 13574 4551 13626
rect 4603 13574 4615 13626
rect 4667 13574 4679 13626
rect 4731 13574 11369 13626
rect 11421 13574 11433 13626
rect 11485 13574 11497 13626
rect 11549 13574 11561 13626
rect 11613 13574 11625 13626
rect 11677 13574 18315 13626
rect 18367 13574 18379 13626
rect 18431 13574 18443 13626
rect 18495 13574 18507 13626
rect 18559 13574 18571 13626
rect 18623 13574 25261 13626
rect 25313 13574 25325 13626
rect 25377 13574 25389 13626
rect 25441 13574 25453 13626
rect 25505 13574 25517 13626
rect 25569 13574 28888 13626
rect 1104 13552 28888 13574
rect 9769 13515 9827 13521
rect 9769 13481 9781 13515
rect 9815 13512 9827 13515
rect 11238 13512 11244 13524
rect 9815 13484 11244 13512
rect 9815 13481 9827 13484
rect 9769 13475 9827 13481
rect 11238 13472 11244 13484
rect 11296 13472 11302 13524
rect 14369 13515 14427 13521
rect 14369 13481 14381 13515
rect 14415 13512 14427 13515
rect 14458 13512 14464 13524
rect 14415 13484 14464 13512
rect 14415 13481 14427 13484
rect 14369 13475 14427 13481
rect 14458 13472 14464 13484
rect 14516 13472 14522 13524
rect 16574 13512 16580 13524
rect 16535 13484 16580 13512
rect 16574 13472 16580 13484
rect 16632 13472 16638 13524
rect 19426 13472 19432 13524
rect 19484 13512 19490 13524
rect 19794 13512 19800 13524
rect 19484 13484 19800 13512
rect 19484 13472 19490 13484
rect 19794 13472 19800 13484
rect 19852 13472 19858 13524
rect 1578 13376 1584 13388
rect 1539 13348 1584 13376
rect 1578 13336 1584 13348
rect 1636 13336 1642 13388
rect 3418 13376 3424 13388
rect 3379 13348 3424 13376
rect 3418 13336 3424 13348
rect 3476 13336 3482 13388
rect 16945 13379 17003 13385
rect 16945 13345 16957 13379
rect 16991 13376 17003 13379
rect 19444 13376 19472 13472
rect 26694 13376 26700 13388
rect 16991 13348 19472 13376
rect 26655 13348 26700 13376
rect 16991 13345 17003 13348
rect 16945 13339 17003 13345
rect 26694 13336 26700 13348
rect 26752 13336 26758 13388
rect 28074 13376 28080 13388
rect 28035 13348 28080 13376
rect 28074 13336 28080 13348
rect 28132 13336 28138 13388
rect 9677 13311 9735 13317
rect 9677 13277 9689 13311
rect 9723 13308 9735 13311
rect 9766 13308 9772 13320
rect 9723 13280 9772 13308
rect 9723 13277 9735 13280
rect 9677 13271 9735 13277
rect 9766 13268 9772 13280
rect 9824 13308 9830 13320
rect 13538 13308 13544 13320
rect 9824 13280 13544 13308
rect 9824 13268 9830 13280
rect 13538 13268 13544 13280
rect 13596 13268 13602 13320
rect 14277 13311 14335 13317
rect 14277 13277 14289 13311
rect 14323 13308 14335 13311
rect 14366 13308 14372 13320
rect 14323 13280 14372 13308
rect 14323 13277 14335 13280
rect 14277 13271 14335 13277
rect 14366 13268 14372 13280
rect 14424 13268 14430 13320
rect 14461 13311 14519 13317
rect 14461 13277 14473 13311
rect 14507 13308 14519 13311
rect 14550 13308 14556 13320
rect 14507 13280 14556 13308
rect 14507 13277 14519 13280
rect 14461 13271 14519 13277
rect 14550 13268 14556 13280
rect 14608 13268 14614 13320
rect 14734 13268 14740 13320
rect 14792 13308 14798 13320
rect 14921 13311 14979 13317
rect 14921 13308 14933 13311
rect 14792 13280 14933 13308
rect 14792 13268 14798 13280
rect 14921 13277 14933 13280
rect 14967 13277 14979 13311
rect 15102 13308 15108 13320
rect 15063 13280 15108 13308
rect 14921 13271 14979 13277
rect 15102 13268 15108 13280
rect 15160 13268 15166 13320
rect 16758 13308 16764 13320
rect 16719 13280 16764 13308
rect 16758 13268 16764 13280
rect 16816 13268 16822 13320
rect 26513 13311 26571 13317
rect 26513 13308 26525 13311
rect 22066 13280 26525 13308
rect 2038 13200 2044 13252
rect 2096 13240 2102 13252
rect 3237 13243 3295 13249
rect 3237 13240 3249 13243
rect 2096 13212 3249 13240
rect 2096 13200 2102 13212
rect 3237 13209 3249 13212
rect 3283 13209 3295 13243
rect 15010 13240 15016 13252
rect 14923 13212 15016 13240
rect 3237 13203 3295 13209
rect 15010 13200 15016 13212
rect 15068 13240 15074 13252
rect 22066 13240 22094 13280
rect 26513 13277 26525 13280
rect 26559 13277 26571 13311
rect 26513 13271 26571 13277
rect 15068 13212 22094 13240
rect 15068 13200 15074 13212
rect 1104 13082 29048 13104
rect 1104 13030 7896 13082
rect 7948 13030 7960 13082
rect 8012 13030 8024 13082
rect 8076 13030 8088 13082
rect 8140 13030 8152 13082
rect 8204 13030 14842 13082
rect 14894 13030 14906 13082
rect 14958 13030 14970 13082
rect 15022 13030 15034 13082
rect 15086 13030 15098 13082
rect 15150 13030 21788 13082
rect 21840 13030 21852 13082
rect 21904 13030 21916 13082
rect 21968 13030 21980 13082
rect 22032 13030 22044 13082
rect 22096 13030 28734 13082
rect 28786 13030 28798 13082
rect 28850 13030 28862 13082
rect 28914 13030 28926 13082
rect 28978 13030 28990 13082
rect 29042 13030 29048 13082
rect 1104 13008 29048 13030
rect 2038 12968 2044 12980
rect 1999 12940 2044 12968
rect 2038 12928 2044 12940
rect 2096 12928 2102 12980
rect 19334 12928 19340 12980
rect 19392 12968 19398 12980
rect 19429 12971 19487 12977
rect 19429 12968 19441 12971
rect 19392 12940 19441 12968
rect 19392 12928 19398 12940
rect 19429 12937 19441 12940
rect 19475 12937 19487 12971
rect 24762 12968 24768 12980
rect 24723 12940 24768 12968
rect 19429 12931 19487 12937
rect 24762 12928 24768 12940
rect 24820 12928 24826 12980
rect 24670 12900 24676 12912
rect 24136 12872 24676 12900
rect 2130 12832 2136 12844
rect 2091 12804 2136 12832
rect 2130 12792 2136 12804
rect 2188 12792 2194 12844
rect 19610 12832 19616 12844
rect 19571 12804 19616 12832
rect 19610 12792 19616 12804
rect 19668 12792 19674 12844
rect 22278 12792 22284 12844
rect 22336 12832 22342 12844
rect 22557 12835 22615 12841
rect 22557 12832 22569 12835
rect 22336 12804 22569 12832
rect 22336 12792 22342 12804
rect 22557 12801 22569 12804
rect 22603 12801 22615 12835
rect 22738 12832 22744 12844
rect 22699 12804 22744 12832
rect 22557 12795 22615 12801
rect 22738 12792 22744 12804
rect 22796 12792 22802 12844
rect 24136 12841 24164 12872
rect 24670 12860 24676 12872
rect 24728 12860 24734 12912
rect 24121 12835 24179 12841
rect 24121 12801 24133 12835
rect 24167 12801 24179 12835
rect 24302 12832 24308 12844
rect 24263 12804 24308 12832
rect 24121 12795 24179 12801
rect 24136 12764 24164 12795
rect 24302 12792 24308 12804
rect 24360 12792 24366 12844
rect 24397 12835 24455 12841
rect 24397 12801 24409 12835
rect 24443 12801 24455 12835
rect 24397 12795 24455 12801
rect 24210 12764 24216 12776
rect 24136 12736 24216 12764
rect 24210 12724 24216 12736
rect 24268 12724 24274 12776
rect 24412 12764 24440 12795
rect 24486 12792 24492 12844
rect 24544 12832 24550 12844
rect 24544 12804 24589 12832
rect 24544 12792 24550 12804
rect 27246 12792 27252 12844
rect 27304 12832 27310 12844
rect 27433 12835 27491 12841
rect 27433 12832 27445 12835
rect 27304 12804 27445 12832
rect 27304 12792 27310 12804
rect 27433 12801 27445 12804
rect 27479 12801 27491 12835
rect 27433 12795 27491 12801
rect 25682 12764 25688 12776
rect 24412 12736 25688 12764
rect 25682 12724 25688 12736
rect 25740 12724 25746 12776
rect 26510 12656 26516 12708
rect 26568 12696 26574 12708
rect 27893 12699 27951 12705
rect 27893 12696 27905 12699
rect 26568 12668 27905 12696
rect 26568 12656 26574 12668
rect 27893 12665 27905 12668
rect 27939 12665 27951 12699
rect 27893 12659 27951 12665
rect 22741 12631 22799 12637
rect 22741 12597 22753 12631
rect 22787 12628 22799 12631
rect 23474 12628 23480 12640
rect 22787 12600 23480 12628
rect 22787 12597 22799 12600
rect 22741 12591 22799 12597
rect 23474 12588 23480 12600
rect 23532 12588 23538 12640
rect 23842 12588 23848 12640
rect 23900 12628 23906 12640
rect 24486 12628 24492 12640
rect 23900 12600 24492 12628
rect 23900 12588 23906 12600
rect 24486 12588 24492 12600
rect 24544 12588 24550 12640
rect 26694 12588 26700 12640
rect 26752 12628 26758 12640
rect 27341 12631 27399 12637
rect 27341 12628 27353 12631
rect 26752 12600 27353 12628
rect 26752 12588 26758 12600
rect 27341 12597 27353 12600
rect 27387 12597 27399 12631
rect 27341 12591 27399 12597
rect 1104 12538 28888 12560
rect 1104 12486 4423 12538
rect 4475 12486 4487 12538
rect 4539 12486 4551 12538
rect 4603 12486 4615 12538
rect 4667 12486 4679 12538
rect 4731 12486 11369 12538
rect 11421 12486 11433 12538
rect 11485 12486 11497 12538
rect 11549 12486 11561 12538
rect 11613 12486 11625 12538
rect 11677 12486 18315 12538
rect 18367 12486 18379 12538
rect 18431 12486 18443 12538
rect 18495 12486 18507 12538
rect 18559 12486 18571 12538
rect 18623 12486 25261 12538
rect 25313 12486 25325 12538
rect 25377 12486 25389 12538
rect 25441 12486 25453 12538
rect 25505 12486 25517 12538
rect 25569 12486 28888 12538
rect 1104 12464 28888 12486
rect 3602 12384 3608 12436
rect 3660 12424 3666 12436
rect 9674 12424 9680 12436
rect 3660 12396 9680 12424
rect 3660 12384 3666 12396
rect 9674 12384 9680 12396
rect 9732 12384 9738 12436
rect 19613 12427 19671 12433
rect 19613 12393 19625 12427
rect 19659 12424 19671 12427
rect 19702 12424 19708 12436
rect 19659 12396 19708 12424
rect 19659 12393 19671 12396
rect 19613 12387 19671 12393
rect 19702 12384 19708 12396
rect 19760 12384 19766 12436
rect 21542 12424 21548 12436
rect 21503 12396 21548 12424
rect 21542 12384 21548 12396
rect 21600 12384 21606 12436
rect 23566 12424 23572 12436
rect 23400 12396 23572 12424
rect 23400 12368 23428 12396
rect 23566 12384 23572 12396
rect 23624 12384 23630 12436
rect 24578 12424 24584 12436
rect 24539 12396 24584 12424
rect 24578 12384 24584 12396
rect 24636 12384 24642 12436
rect 25682 12424 25688 12436
rect 25643 12396 25688 12424
rect 25682 12384 25688 12396
rect 25740 12384 25746 12436
rect 23382 12356 23388 12368
rect 22664 12328 23388 12356
rect 20990 12288 20996 12300
rect 20903 12260 20996 12288
rect 20990 12248 20996 12260
rect 21048 12288 21054 12300
rect 22554 12288 22560 12300
rect 21048 12260 22560 12288
rect 21048 12248 21054 12260
rect 22554 12248 22560 12260
rect 22612 12248 22618 12300
rect 19426 12220 19432 12232
rect 19387 12192 19432 12220
rect 19426 12180 19432 12192
rect 19484 12180 19490 12232
rect 20717 12223 20775 12229
rect 20717 12189 20729 12223
rect 20763 12220 20775 12223
rect 20806 12220 20812 12232
rect 20763 12192 20812 12220
rect 20763 12189 20775 12192
rect 20717 12183 20775 12189
rect 20806 12180 20812 12192
rect 20864 12180 20870 12232
rect 21082 12180 21088 12232
rect 21140 12220 21146 12232
rect 21729 12223 21787 12229
rect 21729 12220 21741 12223
rect 21140 12192 21741 12220
rect 21140 12180 21146 12192
rect 21729 12189 21741 12192
rect 21775 12189 21787 12223
rect 21729 12183 21787 12189
rect 22278 12180 22284 12232
rect 22336 12220 22342 12232
rect 22373 12223 22431 12229
rect 22373 12220 22385 12223
rect 22336 12192 22385 12220
rect 22336 12180 22342 12192
rect 22373 12189 22385 12192
rect 22419 12189 22431 12223
rect 22373 12183 22431 12189
rect 22388 12152 22416 12183
rect 22462 12180 22468 12232
rect 22520 12220 22526 12232
rect 22664 12220 22692 12328
rect 23382 12316 23388 12328
rect 23440 12316 23446 12368
rect 23750 12356 23756 12368
rect 23584 12328 23756 12356
rect 22738 12248 22744 12300
rect 22796 12288 22802 12300
rect 23584 12297 23612 12328
rect 23750 12316 23756 12328
rect 23808 12356 23814 12368
rect 24394 12356 24400 12368
rect 23808 12328 24400 12356
rect 23808 12316 23814 12328
rect 24394 12316 24400 12328
rect 24452 12316 24458 12368
rect 23477 12291 23535 12297
rect 23477 12288 23489 12291
rect 22796 12260 23489 12288
rect 22796 12248 22802 12260
rect 23477 12257 23489 12260
rect 23523 12257 23535 12291
rect 23477 12251 23535 12257
rect 23569 12291 23627 12297
rect 23569 12257 23581 12291
rect 23615 12257 23627 12291
rect 24026 12288 24032 12300
rect 23569 12251 23627 12257
rect 23676 12260 24032 12288
rect 23676 12232 23704 12260
rect 24026 12248 24032 12260
rect 24084 12248 24090 12300
rect 24486 12248 24492 12300
rect 24544 12288 24550 12300
rect 26510 12288 26516 12300
rect 24544 12260 24992 12288
rect 26471 12260 26516 12288
rect 24544 12248 24550 12260
rect 22520 12192 22692 12220
rect 22833 12223 22891 12229
rect 22520 12180 22526 12192
rect 22833 12189 22845 12223
rect 22879 12220 22891 12223
rect 22922 12220 22928 12232
rect 22879 12192 22928 12220
rect 22879 12189 22891 12192
rect 22833 12183 22891 12189
rect 22922 12180 22928 12192
rect 22980 12220 22986 12232
rect 23382 12220 23388 12232
rect 22980 12192 23388 12220
rect 22980 12180 22986 12192
rect 23382 12180 23388 12192
rect 23440 12180 23446 12232
rect 23658 12220 23664 12232
rect 23619 12192 23664 12220
rect 23658 12180 23664 12192
rect 23716 12180 23722 12232
rect 23753 12223 23811 12229
rect 23753 12189 23765 12223
rect 23799 12189 23811 12223
rect 24854 12220 24860 12232
rect 24815 12192 24860 12220
rect 23753 12183 23811 12189
rect 20824 12124 22324 12152
rect 22388 12124 23428 12152
rect 20346 12084 20352 12096
rect 20307 12056 20352 12084
rect 20346 12044 20352 12056
rect 20404 12044 20410 12096
rect 20824 12093 20852 12124
rect 20809 12087 20867 12093
rect 20809 12053 20821 12087
rect 20855 12053 20867 12087
rect 22186 12084 22192 12096
rect 22147 12056 22192 12084
rect 20809 12047 20867 12053
rect 22186 12044 22192 12056
rect 22244 12044 22250 12096
rect 22296 12084 22324 12124
rect 22370 12084 22376 12096
rect 22296 12056 22376 12084
rect 22370 12044 22376 12056
rect 22428 12084 22434 12096
rect 22554 12084 22560 12096
rect 22428 12056 22560 12084
rect 22428 12044 22434 12056
rect 22554 12044 22560 12056
rect 22612 12044 22618 12096
rect 22741 12087 22799 12093
rect 22741 12053 22753 12087
rect 22787 12084 22799 12087
rect 23014 12084 23020 12096
rect 22787 12056 23020 12084
rect 22787 12053 22799 12056
rect 22741 12047 22799 12053
rect 23014 12044 23020 12056
rect 23072 12044 23078 12096
rect 23290 12084 23296 12096
rect 23251 12056 23296 12084
rect 23290 12044 23296 12056
rect 23348 12044 23354 12096
rect 23400 12084 23428 12124
rect 23566 12112 23572 12164
rect 23624 12152 23630 12164
rect 23768 12152 23796 12183
rect 24854 12180 24860 12192
rect 24912 12180 24918 12232
rect 24964 12229 24992 12260
rect 26510 12248 26516 12260
rect 26568 12248 26574 12300
rect 26694 12288 26700 12300
rect 26655 12260 26700 12288
rect 26694 12248 26700 12260
rect 26752 12248 26758 12300
rect 28350 12288 28356 12300
rect 28311 12260 28356 12288
rect 28350 12248 28356 12260
rect 28408 12248 28414 12300
rect 24949 12223 25007 12229
rect 24949 12189 24961 12223
rect 24995 12189 25007 12223
rect 24949 12183 25007 12189
rect 25041 12223 25099 12229
rect 25041 12189 25053 12223
rect 25087 12220 25099 12223
rect 25130 12220 25136 12232
rect 25087 12192 25136 12220
rect 25087 12189 25099 12192
rect 25041 12183 25099 12189
rect 25130 12180 25136 12192
rect 25188 12180 25194 12232
rect 25225 12223 25283 12229
rect 25225 12189 25237 12223
rect 25271 12189 25283 12223
rect 25225 12183 25283 12189
rect 23624 12124 23796 12152
rect 23624 12112 23630 12124
rect 24210 12112 24216 12164
rect 24268 12152 24274 12164
rect 25240 12152 25268 12183
rect 25590 12180 25596 12232
rect 25648 12220 25654 12232
rect 25958 12220 25964 12232
rect 25648 12192 25820 12220
rect 25919 12192 25964 12220
rect 25648 12180 25654 12192
rect 24268 12124 25268 12152
rect 25685 12155 25743 12161
rect 24268 12112 24274 12124
rect 25685 12121 25697 12155
rect 25731 12121 25743 12155
rect 25792 12152 25820 12192
rect 25958 12180 25964 12192
rect 26016 12180 26022 12232
rect 25869 12155 25927 12161
rect 25869 12152 25881 12155
rect 25792 12124 25881 12152
rect 25685 12115 25743 12121
rect 25869 12121 25881 12124
rect 25915 12121 25927 12155
rect 25869 12115 25927 12121
rect 25700 12084 25728 12115
rect 23400 12056 25728 12084
rect 1104 11994 29048 12016
rect 1104 11942 7896 11994
rect 7948 11942 7960 11994
rect 8012 11942 8024 11994
rect 8076 11942 8088 11994
rect 8140 11942 8152 11994
rect 8204 11942 14842 11994
rect 14894 11942 14906 11994
rect 14958 11942 14970 11994
rect 15022 11942 15034 11994
rect 15086 11942 15098 11994
rect 15150 11942 21788 11994
rect 21840 11942 21852 11994
rect 21904 11942 21916 11994
rect 21968 11942 21980 11994
rect 22032 11942 22044 11994
rect 22096 11942 28734 11994
rect 28786 11942 28798 11994
rect 28850 11942 28862 11994
rect 28914 11942 28926 11994
rect 28978 11942 28990 11994
rect 29042 11942 29048 11994
rect 1104 11920 29048 11942
rect 19426 11880 19432 11892
rect 19387 11852 19432 11880
rect 19426 11840 19432 11852
rect 19484 11840 19490 11892
rect 20438 11840 20444 11892
rect 20496 11880 20502 11892
rect 20809 11883 20867 11889
rect 20809 11880 20821 11883
rect 20496 11852 20821 11880
rect 20496 11840 20502 11852
rect 20809 11849 20821 11852
rect 20855 11849 20867 11883
rect 20809 11843 20867 11849
rect 21634 11840 21640 11892
rect 21692 11880 21698 11892
rect 22005 11883 22063 11889
rect 22005 11880 22017 11883
rect 21692 11852 22017 11880
rect 21692 11840 21698 11852
rect 22005 11849 22017 11852
rect 22051 11849 22063 11883
rect 22005 11843 22063 11849
rect 22370 11840 22376 11892
rect 22428 11840 22434 11892
rect 23106 11880 23112 11892
rect 23067 11852 23112 11880
rect 23106 11840 23112 11852
rect 23164 11840 23170 11892
rect 23198 11840 23204 11892
rect 23256 11880 23262 11892
rect 24213 11883 24271 11889
rect 23256 11852 23428 11880
rect 23256 11840 23262 11852
rect 19613 11747 19671 11753
rect 19613 11713 19625 11747
rect 19659 11744 19671 11747
rect 20346 11744 20352 11756
rect 19659 11716 20352 11744
rect 19659 11713 19671 11716
rect 19613 11707 19671 11713
rect 20346 11704 20352 11716
rect 20404 11704 20410 11756
rect 22388 11753 22416 11840
rect 23290 11812 23296 11824
rect 22572 11784 23296 11812
rect 22281 11747 22339 11753
rect 22281 11713 22293 11747
rect 22327 11713 22339 11747
rect 22281 11707 22339 11713
rect 22373 11747 22431 11753
rect 22373 11713 22385 11747
rect 22419 11713 22431 11747
rect 22373 11707 22431 11713
rect 22465 11747 22523 11753
rect 22465 11713 22477 11747
rect 22511 11744 22523 11747
rect 22572 11744 22600 11784
rect 23290 11772 23296 11784
rect 23348 11772 23354 11824
rect 23400 11812 23428 11852
rect 24213 11849 24225 11883
rect 24259 11880 24271 11883
rect 24302 11880 24308 11892
rect 24259 11852 24308 11880
rect 24259 11849 24271 11852
rect 24213 11843 24271 11849
rect 24302 11840 24308 11852
rect 24360 11840 24366 11892
rect 24854 11840 24860 11892
rect 24912 11880 24918 11892
rect 25317 11883 25375 11889
rect 25317 11880 25329 11883
rect 24912 11852 25329 11880
rect 24912 11840 24918 11852
rect 25317 11849 25329 11852
rect 25363 11849 25375 11883
rect 25317 11843 25375 11849
rect 23842 11812 23848 11824
rect 23400 11784 23848 11812
rect 23400 11753 23428 11784
rect 23842 11772 23848 11784
rect 23900 11772 23906 11824
rect 24026 11772 24032 11824
rect 24084 11812 24090 11824
rect 24084 11784 24532 11812
rect 24084 11772 24090 11784
rect 22511 11716 22600 11744
rect 22649 11747 22707 11753
rect 22511 11713 22523 11716
rect 22465 11707 22523 11713
rect 22649 11713 22661 11747
rect 22695 11744 22707 11747
rect 23385 11747 23443 11753
rect 22695 11716 23336 11744
rect 22695 11713 22707 11716
rect 22649 11707 22707 11713
rect 1670 11676 1676 11688
rect 1631 11648 1676 11676
rect 1670 11636 1676 11648
rect 1728 11636 1734 11688
rect 1857 11679 1915 11685
rect 1857 11645 1869 11679
rect 1903 11676 1915 11679
rect 2406 11676 2412 11688
rect 1903 11648 2412 11676
rect 1903 11645 1915 11648
rect 1857 11639 1915 11645
rect 2406 11636 2412 11648
rect 2464 11636 2470 11688
rect 2774 11676 2780 11688
rect 2735 11648 2780 11676
rect 2774 11636 2780 11648
rect 2832 11636 2838 11688
rect 19794 11676 19800 11688
rect 19755 11648 19800 11676
rect 19794 11636 19800 11648
rect 19852 11636 19858 11688
rect 20901 11679 20959 11685
rect 20901 11645 20913 11679
rect 20947 11645 20959 11679
rect 20901 11639 20959 11645
rect 20916 11608 20944 11639
rect 20990 11636 20996 11688
rect 21048 11676 21054 11688
rect 22296 11676 22324 11707
rect 21048 11648 21093 11676
rect 22296 11648 22416 11676
rect 21048 11636 21054 11648
rect 22388 11608 22416 11648
rect 23198 11608 23204 11620
rect 20916 11580 21036 11608
rect 22388 11580 23204 11608
rect 19702 11500 19708 11552
rect 19760 11540 19766 11552
rect 20441 11543 20499 11549
rect 20441 11540 20453 11543
rect 19760 11512 20453 11540
rect 19760 11500 19766 11512
rect 20441 11509 20453 11512
rect 20487 11509 20499 11543
rect 21008 11540 21036 11580
rect 23198 11568 23204 11580
rect 23256 11568 23262 11620
rect 23308 11608 23336 11716
rect 23385 11713 23397 11747
rect 23431 11713 23443 11747
rect 23477 11747 23535 11753
rect 23477 11722 23489 11747
rect 23523 11722 23535 11747
rect 23385 11707 23443 11713
rect 23474 11670 23480 11722
rect 23532 11670 23538 11722
rect 23566 11704 23572 11756
rect 23624 11744 23630 11756
rect 23753 11747 23811 11753
rect 23624 11716 23669 11744
rect 23624 11704 23630 11716
rect 23753 11713 23765 11747
rect 23799 11744 23811 11747
rect 24210 11744 24216 11756
rect 23799 11716 24216 11744
rect 23799 11713 23811 11716
rect 23753 11707 23811 11713
rect 23768 11608 23796 11707
rect 24210 11704 24216 11716
rect 24268 11704 24274 11756
rect 24504 11753 24532 11784
rect 24489 11747 24547 11753
rect 24489 11713 24501 11747
rect 24535 11713 24547 11747
rect 24489 11707 24547 11713
rect 24581 11747 24639 11753
rect 24581 11713 24593 11747
rect 24627 11744 24639 11747
rect 24854 11744 24860 11756
rect 24627 11716 24860 11744
rect 24627 11713 24639 11716
rect 24581 11707 24639 11713
rect 24854 11704 24860 11716
rect 24912 11744 24918 11756
rect 25409 11747 25467 11753
rect 25409 11744 25421 11747
rect 24912 11716 25421 11744
rect 24912 11704 24918 11716
rect 25409 11713 25421 11716
rect 25455 11744 25467 11747
rect 25958 11744 25964 11756
rect 25455 11716 25964 11744
rect 25455 11713 25467 11716
rect 25409 11707 25467 11713
rect 25958 11704 25964 11716
rect 26016 11704 26022 11756
rect 24394 11676 24400 11688
rect 24307 11648 24400 11676
rect 24394 11636 24400 11648
rect 24452 11636 24458 11688
rect 24673 11679 24731 11685
rect 24673 11645 24685 11679
rect 24719 11676 24731 11679
rect 25590 11676 25596 11688
rect 24719 11648 25596 11676
rect 24719 11645 24731 11648
rect 24673 11639 24731 11645
rect 23308 11580 23796 11608
rect 24412 11608 24440 11636
rect 24762 11608 24768 11620
rect 24412 11580 24768 11608
rect 24762 11568 24768 11580
rect 24820 11568 24826 11620
rect 23106 11540 23112 11552
rect 21008 11512 23112 11540
rect 20441 11503 20499 11509
rect 23106 11500 23112 11512
rect 23164 11540 23170 11552
rect 24872 11540 24900 11648
rect 25590 11636 25596 11648
rect 25648 11636 25654 11688
rect 23164 11512 24900 11540
rect 23164 11500 23170 11512
rect 1104 11450 28888 11472
rect 1104 11398 4423 11450
rect 4475 11398 4487 11450
rect 4539 11398 4551 11450
rect 4603 11398 4615 11450
rect 4667 11398 4679 11450
rect 4731 11398 11369 11450
rect 11421 11398 11433 11450
rect 11485 11398 11497 11450
rect 11549 11398 11561 11450
rect 11613 11398 11625 11450
rect 11677 11398 18315 11450
rect 18367 11398 18379 11450
rect 18431 11398 18443 11450
rect 18495 11398 18507 11450
rect 18559 11398 18571 11450
rect 18623 11398 25261 11450
rect 25313 11398 25325 11450
rect 25377 11398 25389 11450
rect 25441 11398 25453 11450
rect 25505 11398 25517 11450
rect 25569 11398 28888 11450
rect 1104 11376 28888 11398
rect 1670 11336 1676 11348
rect 1631 11308 1676 11336
rect 1670 11296 1676 11308
rect 1728 11296 1734 11348
rect 2406 11336 2412 11348
rect 2367 11308 2412 11336
rect 2406 11296 2412 11308
rect 2464 11296 2470 11348
rect 19521 11339 19579 11345
rect 19521 11305 19533 11339
rect 19567 11336 19579 11339
rect 19610 11336 19616 11348
rect 19567 11308 19616 11336
rect 19567 11305 19579 11308
rect 19521 11299 19579 11305
rect 19610 11296 19616 11308
rect 19668 11296 19674 11348
rect 22370 11336 22376 11348
rect 22331 11308 22376 11336
rect 22370 11296 22376 11308
rect 22428 11296 22434 11348
rect 23382 11296 23388 11348
rect 23440 11296 23446 11348
rect 23566 11336 23572 11348
rect 23527 11308 23572 11336
rect 23566 11296 23572 11308
rect 23624 11296 23630 11348
rect 25130 11336 25136 11348
rect 25091 11308 25136 11336
rect 25130 11296 25136 11308
rect 25188 11296 25194 11348
rect 23106 11228 23112 11280
rect 23164 11268 23170 11280
rect 23400 11268 23428 11296
rect 24854 11268 24860 11280
rect 23164 11240 23336 11268
rect 23400 11240 24860 11268
rect 23164 11228 23170 11240
rect 20990 11160 20996 11212
rect 21048 11200 21054 11212
rect 21637 11203 21695 11209
rect 21637 11200 21649 11203
rect 21048 11172 21649 11200
rect 21048 11160 21054 11172
rect 21637 11169 21649 11172
rect 21683 11169 21695 11203
rect 22462 11200 22468 11212
rect 21637 11163 21695 11169
rect 22066 11172 22468 11200
rect 2222 11092 2228 11144
rect 2280 11132 2286 11144
rect 2501 11135 2559 11141
rect 2501 11132 2513 11135
rect 2280 11104 2513 11132
rect 2280 11092 2286 11104
rect 2501 11101 2513 11104
rect 2547 11132 2559 11135
rect 9766 11132 9772 11144
rect 2547 11104 9772 11132
rect 2547 11101 2559 11104
rect 2501 11095 2559 11101
rect 9766 11092 9772 11104
rect 9824 11092 9830 11144
rect 19702 11132 19708 11144
rect 19663 11104 19708 11132
rect 19702 11092 19708 11104
rect 19760 11092 19766 11144
rect 19794 11092 19800 11144
rect 19852 11132 19858 11144
rect 19889 11135 19947 11141
rect 19889 11132 19901 11135
rect 19852 11104 19901 11132
rect 19852 11092 19858 11104
rect 19889 11101 19901 11104
rect 19935 11132 19947 11135
rect 20714 11132 20720 11144
rect 19935 11104 20720 11132
rect 19935 11101 19947 11104
rect 19889 11095 19947 11101
rect 20714 11092 20720 11104
rect 20772 11092 20778 11144
rect 21545 11135 21603 11141
rect 21545 11101 21557 11135
rect 21591 11132 21603 11135
rect 22066 11132 22094 11172
rect 22462 11160 22468 11172
rect 22520 11160 22526 11212
rect 23308 11209 23336 11240
rect 23293 11203 23351 11209
rect 23293 11169 23305 11203
rect 23339 11169 23351 11203
rect 23293 11163 23351 11169
rect 23382 11160 23388 11212
rect 23440 11200 23446 11212
rect 24688 11209 24716 11240
rect 24854 11228 24860 11240
rect 24912 11228 24918 11280
rect 24946 11228 24952 11280
rect 25004 11228 25010 11280
rect 24673 11203 24731 11209
rect 23440 11172 23485 11200
rect 23440 11160 23446 11172
rect 24673 11169 24685 11203
rect 24719 11169 24731 11203
rect 24673 11163 24731 11169
rect 24765 11203 24823 11209
rect 24765 11169 24777 11203
rect 24811 11200 24823 11203
rect 24964 11200 24992 11228
rect 25590 11200 25596 11212
rect 24811 11172 25596 11200
rect 24811 11169 24823 11172
rect 24765 11163 24823 11169
rect 25590 11160 25596 11172
rect 25648 11160 25654 11212
rect 27522 11200 27528 11212
rect 27483 11172 27528 11200
rect 27522 11160 27528 11172
rect 27580 11160 27586 11212
rect 21591 11104 22094 11132
rect 21591 11101 21603 11104
rect 21545 11095 21603 11101
rect 22186 11092 22192 11144
rect 22244 11132 22250 11144
rect 22281 11135 22339 11141
rect 22281 11132 22293 11135
rect 22244 11104 22293 11132
rect 22244 11092 22250 11104
rect 22281 11101 22293 11104
rect 22327 11101 22339 11135
rect 22281 11095 22339 11101
rect 22925 11135 22983 11141
rect 22925 11101 22937 11135
rect 22971 11132 22983 11135
rect 24394 11132 24400 11144
rect 22971 11104 24400 11132
rect 22971 11101 22983 11104
rect 22925 11095 22983 11101
rect 24394 11092 24400 11104
rect 24452 11092 24458 11144
rect 24857 11135 24915 11141
rect 24857 11101 24869 11135
rect 24903 11101 24915 11135
rect 24857 11095 24915 11101
rect 21453 11067 21511 11073
rect 21453 11033 21465 11067
rect 21499 11064 21511 11067
rect 22646 11064 22652 11076
rect 21499 11036 22652 11064
rect 21499 11033 21511 11036
rect 21453 11027 21511 11033
rect 22646 11024 22652 11036
rect 22704 11024 22710 11076
rect 23017 11067 23075 11073
rect 23017 11033 23029 11067
rect 23063 11064 23075 11067
rect 23658 11064 23664 11076
rect 23063 11036 23664 11064
rect 23063 11033 23075 11036
rect 23017 11027 23075 11033
rect 23658 11024 23664 11036
rect 23716 11064 23722 11076
rect 24872 11064 24900 11095
rect 24946 11092 24952 11144
rect 25004 11132 25010 11144
rect 25004 11104 25049 11132
rect 25004 11092 25010 11104
rect 28350 11092 28356 11144
rect 28408 11132 28414 11144
rect 28408 11104 28453 11132
rect 28408 11092 28414 11104
rect 23716 11036 24900 11064
rect 23716 11024 23722 11036
rect 27706 11024 27712 11076
rect 27764 11064 27770 11076
rect 28169 11067 28227 11073
rect 28169 11064 28181 11067
rect 27764 11036 28181 11064
rect 27764 11024 27770 11036
rect 28169 11033 28181 11036
rect 28215 11033 28227 11067
rect 28169 11027 28227 11033
rect 20898 10956 20904 11008
rect 20956 10996 20962 11008
rect 21085 10999 21143 11005
rect 21085 10996 21097 10999
rect 20956 10968 21097 10996
rect 20956 10956 20962 10968
rect 21085 10965 21097 10968
rect 21131 10965 21143 10999
rect 21085 10959 21143 10965
rect 23201 10999 23259 11005
rect 23201 10965 23213 10999
rect 23247 10996 23259 10999
rect 23290 10996 23296 11008
rect 23247 10968 23296 10996
rect 23247 10965 23259 10968
rect 23201 10959 23259 10965
rect 23290 10956 23296 10968
rect 23348 10956 23354 11008
rect 1104 10906 29048 10928
rect 1104 10854 7896 10906
rect 7948 10854 7960 10906
rect 8012 10854 8024 10906
rect 8076 10854 8088 10906
rect 8140 10854 8152 10906
rect 8204 10854 14842 10906
rect 14894 10854 14906 10906
rect 14958 10854 14970 10906
rect 15022 10854 15034 10906
rect 15086 10854 15098 10906
rect 15150 10854 21788 10906
rect 21840 10854 21852 10906
rect 21904 10854 21916 10906
rect 21968 10854 21980 10906
rect 22032 10854 22044 10906
rect 22096 10854 28734 10906
rect 28786 10854 28798 10906
rect 28850 10854 28862 10906
rect 28914 10854 28926 10906
rect 28978 10854 28990 10906
rect 29042 10854 29048 10906
rect 1104 10832 29048 10854
rect 21082 10792 21088 10804
rect 21043 10764 21088 10792
rect 21082 10752 21088 10764
rect 21140 10752 21146 10804
rect 22738 10792 22744 10804
rect 22699 10764 22744 10792
rect 22738 10752 22744 10764
rect 22796 10752 22802 10804
rect 13538 10684 13544 10736
rect 13596 10724 13602 10736
rect 22370 10724 22376 10736
rect 13596 10696 21036 10724
rect 22331 10696 22376 10724
rect 13596 10684 13602 10696
rect 20714 10656 20720 10668
rect 20675 10628 20720 10656
rect 20714 10616 20720 10628
rect 20772 10616 20778 10668
rect 20898 10656 20904 10668
rect 20859 10628 20904 10656
rect 20898 10616 20904 10628
rect 20956 10616 20962 10668
rect 21008 10656 21036 10696
rect 22370 10684 22376 10696
rect 22428 10684 22434 10736
rect 22589 10727 22647 10733
rect 22589 10693 22601 10727
rect 22635 10724 22647 10727
rect 23290 10724 23296 10736
rect 22635 10696 23296 10724
rect 22635 10693 22647 10696
rect 22589 10687 22647 10693
rect 23290 10684 23296 10696
rect 23348 10684 23354 10736
rect 26421 10659 26479 10665
rect 26421 10656 26433 10659
rect 21008 10628 26433 10656
rect 26421 10625 26433 10628
rect 26467 10625 26479 10659
rect 26421 10619 26479 10625
rect 28077 10659 28135 10665
rect 28077 10625 28089 10659
rect 28123 10656 28135 10659
rect 28350 10656 28356 10668
rect 28123 10628 28356 10656
rect 28123 10625 28135 10628
rect 28077 10619 28135 10625
rect 28350 10616 28356 10628
rect 28408 10616 28414 10668
rect 22370 10548 22376 10600
rect 22428 10588 22434 10600
rect 22554 10588 22560 10600
rect 22428 10560 22560 10588
rect 22428 10548 22434 10560
rect 22554 10548 22560 10560
rect 22612 10588 22618 10600
rect 23382 10588 23388 10600
rect 22612 10560 23388 10588
rect 22612 10548 22618 10560
rect 23382 10548 23388 10560
rect 23440 10548 23446 10600
rect 22557 10455 22615 10461
rect 22557 10421 22569 10455
rect 22603 10452 22615 10455
rect 23106 10452 23112 10464
rect 22603 10424 23112 10452
rect 22603 10421 22615 10424
rect 22557 10415 22615 10421
rect 23106 10412 23112 10424
rect 23164 10412 23170 10464
rect 26513 10455 26571 10461
rect 26513 10421 26525 10455
rect 26559 10452 26571 10455
rect 26694 10452 26700 10464
rect 26559 10424 26700 10452
rect 26559 10421 26571 10424
rect 26513 10415 26571 10421
rect 26694 10412 26700 10424
rect 26752 10412 26758 10464
rect 27154 10452 27160 10464
rect 27115 10424 27160 10452
rect 27154 10412 27160 10424
rect 27212 10412 27218 10464
rect 1104 10362 28888 10384
rect 1104 10310 4423 10362
rect 4475 10310 4487 10362
rect 4539 10310 4551 10362
rect 4603 10310 4615 10362
rect 4667 10310 4679 10362
rect 4731 10310 11369 10362
rect 11421 10310 11433 10362
rect 11485 10310 11497 10362
rect 11549 10310 11561 10362
rect 11613 10310 11625 10362
rect 11677 10310 18315 10362
rect 18367 10310 18379 10362
rect 18431 10310 18443 10362
rect 18495 10310 18507 10362
rect 18559 10310 18571 10362
rect 18623 10310 25261 10362
rect 25313 10310 25325 10362
rect 25377 10310 25389 10362
rect 25441 10310 25453 10362
rect 25505 10310 25517 10362
rect 25569 10310 28888 10362
rect 1104 10288 28888 10310
rect 27154 10180 27160 10192
rect 26528 10152 27160 10180
rect 26528 10121 26556 10152
rect 27154 10140 27160 10152
rect 27212 10140 27218 10192
rect 26513 10115 26571 10121
rect 26513 10081 26525 10115
rect 26559 10081 26571 10115
rect 26694 10112 26700 10124
rect 26655 10084 26700 10112
rect 26513 10075 26571 10081
rect 26694 10072 26700 10084
rect 26752 10072 26758 10124
rect 28353 10115 28411 10121
rect 28353 10081 28365 10115
rect 28399 10112 28411 10115
rect 29914 10112 29920 10124
rect 28399 10084 29920 10112
rect 28399 10081 28411 10084
rect 28353 10075 28411 10081
rect 29914 10072 29920 10084
rect 29972 10072 29978 10124
rect 1670 10004 1676 10056
rect 1728 10044 1734 10056
rect 1765 10047 1823 10053
rect 1765 10044 1777 10047
rect 1728 10016 1777 10044
rect 1728 10004 1734 10016
rect 1765 10013 1777 10016
rect 1811 10013 1823 10047
rect 3050 10044 3056 10056
rect 3011 10016 3056 10044
rect 1765 10007 1823 10013
rect 3050 10004 3056 10016
rect 3108 10004 3114 10056
rect 1104 9818 29048 9840
rect 1104 9766 7896 9818
rect 7948 9766 7960 9818
rect 8012 9766 8024 9818
rect 8076 9766 8088 9818
rect 8140 9766 8152 9818
rect 8204 9766 14842 9818
rect 14894 9766 14906 9818
rect 14958 9766 14970 9818
rect 15022 9766 15034 9818
rect 15086 9766 15098 9818
rect 15150 9766 21788 9818
rect 21840 9766 21852 9818
rect 21904 9766 21916 9818
rect 21968 9766 21980 9818
rect 22032 9766 22044 9818
rect 22096 9766 28734 9818
rect 28786 9766 28798 9818
rect 28850 9766 28862 9818
rect 28914 9766 28926 9818
rect 28978 9766 28990 9818
rect 29042 9766 29048 9818
rect 1104 9744 29048 9766
rect 25682 9636 25688 9648
rect 2884 9608 25688 9636
rect 2498 9568 2504 9580
rect 2411 9540 2504 9568
rect 2498 9528 2504 9540
rect 2556 9568 2562 9580
rect 2884 9568 2912 9608
rect 25682 9596 25688 9608
rect 25740 9596 25746 9648
rect 27706 9636 27712 9648
rect 27667 9608 27712 9636
rect 27706 9596 27712 9608
rect 27764 9596 27770 9648
rect 3050 9568 3056 9580
rect 2556 9540 2912 9568
rect 3011 9540 3056 9568
rect 2556 9528 2562 9540
rect 3050 9528 3056 9540
rect 3108 9528 3114 9580
rect 21358 9528 21364 9580
rect 21416 9568 21422 9580
rect 25961 9571 26019 9577
rect 25961 9568 25973 9571
rect 21416 9540 25973 9568
rect 21416 9528 21422 9540
rect 25961 9537 25973 9540
rect 26007 9537 26019 9571
rect 27614 9568 27620 9580
rect 27575 9540 27620 9568
rect 25961 9531 26019 9537
rect 27614 9528 27620 9540
rect 27672 9528 27678 9580
rect 3237 9503 3295 9509
rect 3237 9469 3249 9503
rect 3283 9500 3295 9503
rect 4062 9500 4068 9512
rect 3283 9472 4068 9500
rect 3283 9469 3295 9472
rect 3237 9463 3295 9469
rect 4062 9460 4068 9472
rect 4120 9460 4126 9512
rect 4154 9460 4160 9512
rect 4212 9500 4218 9512
rect 4212 9472 4257 9500
rect 4212 9460 4218 9472
rect 1578 9324 1584 9376
rect 1636 9364 1642 9376
rect 1673 9367 1731 9373
rect 1673 9364 1685 9367
rect 1636 9336 1685 9364
rect 1636 9324 1642 9336
rect 1673 9333 1685 9336
rect 1719 9333 1731 9367
rect 1673 9327 1731 9333
rect 1762 9324 1768 9376
rect 1820 9364 1826 9376
rect 2409 9367 2467 9373
rect 2409 9364 2421 9367
rect 1820 9336 2421 9364
rect 1820 9324 1826 9336
rect 2409 9333 2421 9336
rect 2455 9333 2467 9367
rect 2409 9327 2467 9333
rect 25774 9324 25780 9376
rect 25832 9364 25838 9376
rect 25869 9367 25927 9373
rect 25869 9364 25881 9367
rect 25832 9336 25881 9364
rect 25832 9324 25838 9336
rect 25869 9333 25881 9336
rect 25915 9333 25927 9367
rect 25869 9327 25927 9333
rect 1104 9274 28888 9296
rect 1104 9222 4423 9274
rect 4475 9222 4487 9274
rect 4539 9222 4551 9274
rect 4603 9222 4615 9274
rect 4667 9222 4679 9274
rect 4731 9222 11369 9274
rect 11421 9222 11433 9274
rect 11485 9222 11497 9274
rect 11549 9222 11561 9274
rect 11613 9222 11625 9274
rect 11677 9222 18315 9274
rect 18367 9222 18379 9274
rect 18431 9222 18443 9274
rect 18495 9222 18507 9274
rect 18559 9222 18571 9274
rect 18623 9222 25261 9274
rect 25313 9222 25325 9274
rect 25377 9222 25389 9274
rect 25441 9222 25453 9274
rect 25505 9222 25517 9274
rect 25569 9222 28888 9274
rect 1104 9200 28888 9222
rect 4062 9160 4068 9172
rect 4023 9132 4068 9160
rect 4062 9120 4068 9132
rect 4120 9120 4126 9172
rect 1578 9024 1584 9036
rect 1539 8996 1584 9024
rect 1578 8984 1584 8996
rect 1636 8984 1642 9036
rect 1762 9024 1768 9036
rect 1723 8996 1768 9024
rect 1762 8984 1768 8996
rect 1820 8984 1826 9036
rect 2774 9024 2780 9036
rect 2735 8996 2780 9024
rect 2774 8984 2780 8996
rect 2832 8984 2838 9036
rect 25590 9024 25596 9036
rect 25551 8996 25596 9024
rect 25590 8984 25596 8996
rect 25648 8984 25654 9036
rect 25774 9024 25780 9036
rect 25735 8996 25780 9024
rect 25774 8984 25780 8996
rect 25832 8984 25838 9036
rect 4157 8959 4215 8965
rect 4157 8925 4169 8959
rect 4203 8956 4215 8959
rect 4338 8956 4344 8968
rect 4203 8928 4344 8956
rect 4203 8925 4215 8928
rect 4157 8919 4215 8925
rect 4338 8916 4344 8928
rect 4396 8916 4402 8968
rect 28077 8959 28135 8965
rect 28077 8925 28089 8959
rect 28123 8956 28135 8959
rect 28350 8956 28356 8968
rect 28123 8928 28356 8956
rect 28123 8925 28135 8928
rect 28077 8919 28135 8925
rect 28350 8916 28356 8928
rect 28408 8916 28414 8968
rect 27433 8891 27491 8897
rect 27433 8857 27445 8891
rect 27479 8888 27491 8891
rect 29914 8888 29920 8900
rect 27479 8860 29920 8888
rect 27479 8857 27491 8860
rect 27433 8851 27491 8857
rect 29914 8848 29920 8860
rect 29972 8848 29978 8900
rect 1104 8730 29048 8752
rect 1104 8678 7896 8730
rect 7948 8678 7960 8730
rect 8012 8678 8024 8730
rect 8076 8678 8088 8730
rect 8140 8678 8152 8730
rect 8204 8678 14842 8730
rect 14894 8678 14906 8730
rect 14958 8678 14970 8730
rect 15022 8678 15034 8730
rect 15086 8678 15098 8730
rect 15150 8678 21788 8730
rect 21840 8678 21852 8730
rect 21904 8678 21916 8730
rect 21968 8678 21980 8730
rect 22032 8678 22044 8730
rect 22096 8678 28734 8730
rect 28786 8678 28798 8730
rect 28850 8678 28862 8730
rect 28914 8678 28926 8730
rect 28978 8678 28990 8730
rect 29042 8678 29048 8730
rect 1104 8656 29048 8678
rect 12710 8548 12716 8560
rect 4816 8520 12716 8548
rect 1670 8480 1676 8492
rect 1631 8452 1676 8480
rect 1670 8440 1676 8452
rect 1728 8440 1734 8492
rect 4816 8489 4844 8520
rect 12710 8508 12716 8520
rect 12768 8508 12774 8560
rect 4801 8483 4859 8489
rect 4801 8449 4813 8483
rect 4847 8449 4859 8483
rect 9309 8483 9367 8489
rect 9309 8480 9321 8483
rect 4801 8443 4859 8449
rect 6886 8452 9321 8480
rect 1854 8412 1860 8424
rect 1815 8384 1860 8412
rect 1854 8372 1860 8384
rect 1912 8372 1918 8424
rect 2774 8412 2780 8424
rect 2735 8384 2780 8412
rect 2774 8372 2780 8384
rect 2832 8372 2838 8424
rect 4338 8372 4344 8424
rect 4396 8412 4402 8424
rect 6886 8412 6914 8452
rect 9309 8449 9321 8452
rect 9355 8449 9367 8483
rect 27706 8480 27712 8492
rect 27619 8452 27712 8480
rect 9309 8443 9367 8449
rect 27706 8440 27712 8452
rect 27764 8480 27770 8492
rect 28534 8480 28540 8492
rect 27764 8452 28540 8480
rect 27764 8440 27770 8452
rect 28534 8440 28540 8452
rect 28592 8440 28598 8492
rect 4396 8384 6914 8412
rect 4396 8372 4402 8384
rect 9398 8344 9404 8356
rect 9359 8316 9404 8344
rect 9398 8304 9404 8316
rect 9456 8304 9462 8356
rect 3970 8276 3976 8288
rect 3931 8248 3976 8276
rect 3970 8236 3976 8248
rect 4028 8236 4034 8288
rect 4154 8236 4160 8288
rect 4212 8276 4218 8288
rect 4709 8279 4767 8285
rect 4709 8276 4721 8279
rect 4212 8248 4721 8276
rect 4212 8236 4218 8248
rect 4709 8245 4721 8248
rect 4755 8245 4767 8279
rect 26602 8276 26608 8288
rect 26563 8248 26608 8276
rect 4709 8239 4767 8245
rect 26602 8236 26608 8248
rect 26660 8236 26666 8288
rect 27801 8279 27859 8285
rect 27801 8245 27813 8279
rect 27847 8276 27859 8279
rect 28166 8276 28172 8288
rect 27847 8248 28172 8276
rect 27847 8245 27859 8248
rect 27801 8239 27859 8245
rect 28166 8236 28172 8248
rect 28224 8236 28230 8288
rect 1104 8186 28888 8208
rect 1104 8134 4423 8186
rect 4475 8134 4487 8186
rect 4539 8134 4551 8186
rect 4603 8134 4615 8186
rect 4667 8134 4679 8186
rect 4731 8134 11369 8186
rect 11421 8134 11433 8186
rect 11485 8134 11497 8186
rect 11549 8134 11561 8186
rect 11613 8134 11625 8186
rect 11677 8134 18315 8186
rect 18367 8134 18379 8186
rect 18431 8134 18443 8186
rect 18495 8134 18507 8186
rect 18559 8134 18571 8186
rect 18623 8134 25261 8186
rect 25313 8134 25325 8186
rect 25377 8134 25389 8186
rect 25441 8134 25453 8186
rect 25505 8134 25517 8186
rect 25569 8134 28888 8186
rect 1104 8112 28888 8134
rect 1854 8032 1860 8084
rect 1912 8072 1918 8084
rect 2133 8075 2191 8081
rect 2133 8072 2145 8075
rect 1912 8044 2145 8072
rect 1912 8032 1918 8044
rect 2133 8041 2145 8044
rect 2179 8041 2191 8075
rect 2133 8035 2191 8041
rect 3970 7936 3976 7948
rect 3931 7908 3976 7936
rect 3970 7896 3976 7908
rect 4028 7896 4034 7948
rect 4154 7936 4160 7948
rect 4115 7908 4160 7936
rect 4154 7896 4160 7908
rect 4212 7896 4218 7948
rect 5534 7936 5540 7948
rect 5495 7908 5540 7936
rect 5534 7896 5540 7908
rect 5592 7896 5598 7948
rect 27522 7936 27528 7948
rect 27483 7908 27528 7936
rect 27522 7896 27528 7908
rect 27580 7896 27586 7948
rect 28166 7936 28172 7948
rect 28127 7908 28172 7936
rect 28166 7896 28172 7908
rect 28224 7896 28230 7948
rect 28350 7936 28356 7948
rect 28311 7908 28356 7936
rect 28350 7896 28356 7908
rect 28408 7896 28414 7948
rect 2225 7871 2283 7877
rect 2225 7837 2237 7871
rect 2271 7868 2283 7871
rect 2406 7868 2412 7880
rect 2271 7840 2412 7868
rect 2271 7837 2283 7840
rect 2225 7831 2283 7837
rect 2406 7828 2412 7840
rect 2464 7828 2470 7880
rect 1104 7642 29048 7664
rect 1104 7590 7896 7642
rect 7948 7590 7960 7642
rect 8012 7590 8024 7642
rect 8076 7590 8088 7642
rect 8140 7590 8152 7642
rect 8204 7590 14842 7642
rect 14894 7590 14906 7642
rect 14958 7590 14970 7642
rect 15022 7590 15034 7642
rect 15086 7590 15098 7642
rect 15150 7590 21788 7642
rect 21840 7590 21852 7642
rect 21904 7590 21916 7642
rect 21968 7590 21980 7642
rect 22032 7590 22044 7642
rect 22096 7590 28734 7642
rect 28786 7590 28798 7642
rect 28850 7590 28862 7642
rect 28914 7590 28926 7642
rect 28978 7590 28990 7642
rect 29042 7590 29048 7642
rect 1104 7568 29048 7590
rect 2222 7392 2228 7404
rect 2183 7364 2228 7392
rect 2222 7352 2228 7364
rect 2280 7352 2286 7404
rect 26602 7352 26608 7404
rect 26660 7392 26666 7404
rect 27617 7395 27675 7401
rect 26660 7364 26705 7392
rect 26660 7352 26666 7364
rect 27617 7361 27629 7395
rect 27663 7392 27675 7395
rect 28258 7392 28264 7404
rect 27663 7364 28264 7392
rect 27663 7361 27675 7364
rect 27617 7355 27675 7361
rect 28258 7352 28264 7364
rect 28316 7352 28322 7404
rect 26142 7324 26148 7336
rect 26103 7296 26148 7324
rect 26142 7284 26148 7296
rect 26200 7284 26206 7336
rect 26421 7327 26479 7333
rect 26421 7293 26433 7327
rect 26467 7324 26479 7327
rect 27709 7327 27767 7333
rect 27709 7324 27721 7327
rect 26467 7296 27721 7324
rect 26467 7293 26479 7296
rect 26421 7287 26479 7293
rect 27709 7293 27721 7296
rect 27755 7293 27767 7327
rect 27709 7287 27767 7293
rect 1762 7148 1768 7200
rect 1820 7188 1826 7200
rect 2133 7191 2191 7197
rect 2133 7188 2145 7191
rect 1820 7160 2145 7188
rect 1820 7148 1826 7160
rect 2133 7157 2145 7160
rect 2179 7157 2191 7191
rect 2133 7151 2191 7157
rect 2958 7148 2964 7200
rect 3016 7188 3022 7200
rect 3053 7191 3111 7197
rect 3053 7188 3065 7191
rect 3016 7160 3065 7188
rect 3016 7148 3022 7160
rect 3053 7157 3065 7160
rect 3099 7157 3111 7191
rect 3053 7151 3111 7157
rect 1104 7098 28888 7120
rect 1104 7046 4423 7098
rect 4475 7046 4487 7098
rect 4539 7046 4551 7098
rect 4603 7046 4615 7098
rect 4667 7046 4679 7098
rect 4731 7046 11369 7098
rect 11421 7046 11433 7098
rect 11485 7046 11497 7098
rect 11549 7046 11561 7098
rect 11613 7046 11625 7098
rect 11677 7046 18315 7098
rect 18367 7046 18379 7098
rect 18431 7046 18443 7098
rect 18495 7046 18507 7098
rect 18559 7046 18571 7098
rect 18623 7046 25261 7098
rect 25313 7046 25325 7098
rect 25377 7046 25389 7098
rect 25441 7046 25453 7098
rect 25505 7046 25517 7098
rect 25569 7046 28888 7098
rect 1104 7024 28888 7046
rect 1762 6848 1768 6860
rect 1723 6820 1768 6848
rect 1762 6808 1768 6820
rect 1820 6808 1826 6860
rect 2774 6848 2780 6860
rect 2735 6820 2780 6848
rect 2774 6808 2780 6820
rect 2832 6808 2838 6860
rect 19610 6808 19616 6860
rect 19668 6848 19674 6860
rect 24581 6851 24639 6857
rect 24581 6848 24593 6851
rect 19668 6820 24593 6848
rect 19668 6808 19674 6820
rect 24581 6817 24593 6820
rect 24627 6817 24639 6851
rect 25130 6848 25136 6860
rect 25091 6820 25136 6848
rect 24581 6811 24639 6817
rect 25130 6808 25136 6820
rect 25188 6808 25194 6860
rect 1578 6780 1584 6792
rect 1539 6752 1584 6780
rect 1578 6740 1584 6752
rect 1636 6740 1642 6792
rect 23845 6783 23903 6789
rect 23845 6749 23857 6783
rect 23891 6749 23903 6783
rect 23845 6743 23903 6749
rect 23860 6656 23888 6743
rect 26602 6740 26608 6792
rect 26660 6780 26666 6792
rect 27617 6783 27675 6789
rect 27617 6780 27629 6783
rect 26660 6752 27629 6780
rect 26660 6740 26666 6752
rect 27617 6749 27629 6752
rect 27663 6749 27675 6783
rect 27617 6743 27675 6749
rect 23937 6715 23995 6721
rect 23937 6681 23949 6715
rect 23983 6712 23995 6715
rect 24765 6715 24823 6721
rect 24765 6712 24777 6715
rect 23983 6684 24777 6712
rect 23983 6681 23995 6684
rect 23937 6675 23995 6681
rect 24765 6681 24777 6684
rect 24811 6681 24823 6715
rect 24765 6675 24823 6681
rect 23842 6644 23848 6656
rect 23755 6616 23848 6644
rect 23842 6604 23848 6616
rect 23900 6644 23906 6656
rect 27338 6644 27344 6656
rect 23900 6616 27344 6644
rect 23900 6604 23906 6616
rect 27338 6604 27344 6616
rect 27396 6604 27402 6656
rect 1104 6554 29048 6576
rect 1104 6502 7896 6554
rect 7948 6502 7960 6554
rect 8012 6502 8024 6554
rect 8076 6502 8088 6554
rect 8140 6502 8152 6554
rect 8204 6502 14842 6554
rect 14894 6502 14906 6554
rect 14958 6502 14970 6554
rect 15022 6502 15034 6554
rect 15086 6502 15098 6554
rect 15150 6502 21788 6554
rect 21840 6502 21852 6554
rect 21904 6502 21916 6554
rect 21968 6502 21980 6554
rect 22032 6502 22044 6554
rect 22096 6502 28734 6554
rect 28786 6502 28798 6554
rect 28850 6502 28862 6554
rect 28914 6502 28926 6554
rect 28978 6502 28990 6554
rect 29042 6502 29048 6554
rect 1104 6480 29048 6502
rect 26421 6375 26479 6381
rect 26421 6341 26433 6375
rect 26467 6372 26479 6375
rect 27525 6375 27583 6381
rect 27525 6372 27537 6375
rect 26467 6344 27537 6372
rect 26467 6341 26479 6344
rect 26421 6335 26479 6341
rect 27525 6341 27537 6344
rect 27571 6341 27583 6375
rect 27525 6335 27583 6341
rect 1578 6264 1584 6316
rect 1636 6304 1642 6316
rect 1673 6307 1731 6313
rect 1673 6304 1685 6307
rect 1636 6276 1685 6304
rect 1636 6264 1642 6276
rect 1673 6273 1685 6276
rect 1719 6273 1731 6307
rect 2314 6304 2320 6316
rect 2227 6276 2320 6304
rect 1673 6267 1731 6273
rect 2314 6264 2320 6276
rect 2372 6264 2378 6316
rect 2958 6304 2964 6316
rect 2919 6276 2964 6304
rect 2958 6264 2964 6276
rect 3016 6264 3022 6316
rect 26602 6264 26608 6316
rect 26660 6304 26666 6316
rect 26660 6276 26705 6304
rect 26660 6264 26666 6276
rect 27338 6264 27344 6316
rect 27396 6304 27402 6316
rect 27433 6307 27491 6313
rect 27433 6304 27445 6307
rect 27396 6276 27445 6304
rect 27396 6264 27402 6276
rect 27433 6273 27445 6276
rect 27479 6273 27491 6307
rect 27433 6267 27491 6273
rect 2332 6168 2360 6264
rect 2409 6239 2467 6245
rect 2409 6205 2421 6239
rect 2455 6236 2467 6239
rect 3145 6239 3203 6245
rect 3145 6236 3157 6239
rect 2455 6208 3157 6236
rect 2455 6205 2467 6208
rect 2409 6199 2467 6205
rect 3145 6205 3157 6208
rect 3191 6205 3203 6239
rect 4154 6236 4160 6248
rect 4115 6208 4160 6236
rect 3145 6199 3203 6205
rect 4154 6196 4160 6208
rect 4212 6196 4218 6248
rect 26142 6236 26148 6248
rect 26103 6208 26148 6236
rect 26142 6196 26148 6208
rect 26200 6196 26206 6248
rect 5350 6168 5356 6180
rect 2332 6140 5356 6168
rect 5350 6128 5356 6140
rect 5408 6128 5414 6180
rect 1104 6010 28888 6032
rect 1104 5958 4423 6010
rect 4475 5958 4487 6010
rect 4539 5958 4551 6010
rect 4603 5958 4615 6010
rect 4667 5958 4679 6010
rect 4731 5958 11369 6010
rect 11421 5958 11433 6010
rect 11485 5958 11497 6010
rect 11549 5958 11561 6010
rect 11613 5958 11625 6010
rect 11677 5958 18315 6010
rect 18367 5958 18379 6010
rect 18431 5958 18443 6010
rect 18495 5958 18507 6010
rect 18559 5958 18571 6010
rect 18623 5958 25261 6010
rect 25313 5958 25325 6010
rect 25377 5958 25389 6010
rect 25441 5958 25453 6010
rect 25505 5958 25517 6010
rect 25569 5958 28888 6010
rect 1104 5936 28888 5958
rect 25682 5788 25688 5840
rect 25740 5828 25746 5840
rect 27706 5828 27712 5840
rect 25740 5800 27712 5828
rect 25740 5788 25746 5800
rect 3050 5760 3056 5772
rect 3011 5732 3056 5760
rect 3050 5720 3056 5732
rect 3108 5720 3114 5772
rect 25884 5769 25912 5800
rect 27706 5788 27712 5800
rect 27764 5788 27770 5840
rect 25869 5763 25927 5769
rect 25869 5729 25881 5763
rect 25915 5729 25927 5763
rect 25869 5723 25927 5729
rect 1578 5692 1584 5704
rect 1539 5664 1584 5692
rect 1578 5652 1584 5664
rect 1636 5652 1642 5704
rect 4154 5652 4160 5704
rect 4212 5692 4218 5704
rect 4709 5695 4767 5701
rect 4709 5692 4721 5695
rect 4212 5664 4721 5692
rect 4212 5652 4218 5664
rect 4709 5661 4721 5664
rect 4755 5661 4767 5695
rect 4709 5655 4767 5661
rect 24946 5652 24952 5704
rect 25004 5692 25010 5704
rect 25317 5695 25375 5701
rect 25317 5692 25329 5695
rect 25004 5664 25329 5692
rect 25004 5652 25010 5664
rect 25317 5661 25329 5664
rect 25363 5692 25375 5695
rect 26234 5692 26240 5704
rect 25363 5664 26240 5692
rect 25363 5661 25375 5664
rect 25317 5655 25375 5661
rect 26234 5652 26240 5664
rect 26292 5652 26298 5704
rect 26418 5692 26424 5704
rect 26379 5664 26424 5692
rect 26418 5652 26424 5664
rect 26476 5652 26482 5704
rect 1762 5624 1768 5636
rect 1723 5596 1768 5624
rect 1762 5584 1768 5596
rect 1820 5584 1826 5636
rect 26602 5624 26608 5636
rect 26563 5596 26608 5624
rect 26602 5584 26608 5596
rect 26660 5584 26666 5636
rect 28261 5627 28319 5633
rect 28261 5593 28273 5627
rect 28307 5624 28319 5627
rect 29914 5624 29920 5636
rect 28307 5596 29920 5624
rect 28307 5593 28319 5596
rect 28261 5587 28319 5593
rect 29914 5584 29920 5596
rect 29972 5584 29978 5636
rect 1104 5466 29048 5488
rect 1104 5414 7896 5466
rect 7948 5414 7960 5466
rect 8012 5414 8024 5466
rect 8076 5414 8088 5466
rect 8140 5414 8152 5466
rect 8204 5414 14842 5466
rect 14894 5414 14906 5466
rect 14958 5414 14970 5466
rect 15022 5414 15034 5466
rect 15086 5414 15098 5466
rect 15150 5414 21788 5466
rect 21840 5414 21852 5466
rect 21904 5414 21916 5466
rect 21968 5414 21980 5466
rect 22032 5414 22044 5466
rect 22096 5414 28734 5466
rect 28786 5414 28798 5466
rect 28850 5414 28862 5466
rect 28914 5414 28926 5466
rect 28978 5414 28990 5466
rect 29042 5414 29048 5466
rect 1104 5392 29048 5414
rect 1762 5312 1768 5364
rect 1820 5352 1826 5364
rect 2409 5355 2467 5361
rect 2409 5352 2421 5355
rect 1820 5324 2421 5352
rect 1820 5312 1826 5324
rect 2409 5321 2421 5324
rect 2455 5321 2467 5355
rect 2409 5315 2467 5321
rect 26421 5355 26479 5361
rect 26421 5321 26433 5355
rect 26467 5352 26479 5355
rect 26602 5352 26608 5364
rect 26467 5324 26608 5352
rect 26467 5321 26479 5324
rect 26421 5315 26479 5321
rect 26602 5312 26608 5324
rect 26660 5312 26666 5364
rect 2038 5244 2044 5296
rect 2096 5284 2102 5296
rect 10502 5284 10508 5296
rect 2096 5256 10508 5284
rect 2096 5244 2102 5256
rect 1578 5176 1584 5228
rect 1636 5216 1642 5228
rect 2516 5225 2544 5256
rect 10502 5244 10508 5256
rect 10560 5244 10566 5296
rect 26234 5244 26240 5296
rect 26292 5284 26298 5296
rect 27062 5284 27068 5296
rect 26292 5256 27068 5284
rect 26292 5244 26298 5256
rect 1673 5219 1731 5225
rect 1673 5216 1685 5219
rect 1636 5188 1685 5216
rect 1636 5176 1642 5188
rect 1673 5185 1685 5188
rect 1719 5185 1731 5219
rect 1673 5179 1731 5185
rect 2501 5219 2559 5225
rect 2501 5185 2513 5219
rect 2547 5185 2559 5219
rect 5350 5216 5356 5228
rect 5311 5188 5356 5216
rect 2501 5179 2559 5185
rect 5350 5176 5356 5188
rect 5408 5176 5414 5228
rect 26344 5225 26372 5256
rect 27062 5244 27068 5256
rect 27120 5244 27126 5296
rect 26329 5219 26387 5225
rect 26329 5185 26341 5219
rect 26375 5185 26387 5219
rect 26329 5179 26387 5185
rect 26418 5176 26424 5228
rect 26476 5216 26482 5228
rect 27157 5219 27215 5225
rect 27157 5216 27169 5219
rect 26476 5188 27169 5216
rect 26476 5176 26482 5188
rect 27157 5185 27169 5188
rect 27203 5185 27215 5219
rect 27157 5179 27215 5185
rect 2958 5148 2964 5160
rect 2919 5120 2964 5148
rect 2958 5108 2964 5120
rect 3016 5108 3022 5160
rect 3142 5148 3148 5160
rect 3103 5120 3148 5148
rect 3142 5108 3148 5120
rect 3200 5108 3206 5160
rect 4798 5148 4804 5160
rect 4759 5120 4804 5148
rect 4798 5108 4804 5120
rect 4856 5108 4862 5160
rect 5442 5012 5448 5024
rect 5403 4984 5448 5012
rect 5442 4972 5448 4984
rect 5500 4972 5506 5024
rect 26602 4972 26608 5024
rect 26660 5012 26666 5024
rect 27893 5015 27951 5021
rect 27893 5012 27905 5015
rect 26660 4984 27905 5012
rect 26660 4972 26666 4984
rect 27893 4981 27905 4984
rect 27939 4981 27951 5015
rect 27893 4975 27951 4981
rect 1104 4922 28888 4944
rect 1104 4870 4423 4922
rect 4475 4870 4487 4922
rect 4539 4870 4551 4922
rect 4603 4870 4615 4922
rect 4667 4870 4679 4922
rect 4731 4870 11369 4922
rect 11421 4870 11433 4922
rect 11485 4870 11497 4922
rect 11549 4870 11561 4922
rect 11613 4870 11625 4922
rect 11677 4870 18315 4922
rect 18367 4870 18379 4922
rect 18431 4870 18443 4922
rect 18495 4870 18507 4922
rect 18559 4870 18571 4922
rect 18623 4870 25261 4922
rect 25313 4870 25325 4922
rect 25377 4870 25389 4922
rect 25441 4870 25453 4922
rect 25505 4870 25517 4922
rect 25569 4870 28888 4922
rect 1104 4848 28888 4870
rect 2958 4808 2964 4820
rect 2919 4780 2964 4808
rect 2958 4768 2964 4780
rect 3016 4768 3022 4820
rect 5442 4672 5448 4684
rect 5403 4644 5448 4672
rect 5442 4632 5448 4644
rect 5500 4632 5506 4684
rect 5810 4672 5816 4684
rect 5771 4644 5816 4672
rect 5810 4632 5816 4644
rect 5868 4632 5874 4684
rect 23937 4675 23995 4681
rect 23937 4641 23949 4675
rect 23983 4672 23995 4675
rect 25038 4672 25044 4684
rect 23983 4644 25044 4672
rect 23983 4641 23995 4644
rect 23937 4635 23995 4641
rect 25038 4632 25044 4644
rect 25096 4632 25102 4684
rect 27430 4672 27436 4684
rect 27391 4644 27436 4672
rect 27430 4632 27436 4644
rect 27488 4632 27494 4684
rect 1578 4604 1584 4616
rect 1539 4576 1584 4604
rect 1578 4564 1584 4576
rect 1636 4564 1642 4616
rect 2409 4607 2467 4613
rect 2409 4573 2421 4607
rect 2455 4604 2467 4607
rect 2498 4604 2504 4616
rect 2455 4576 2504 4604
rect 2455 4573 2467 4576
rect 2409 4567 2467 4573
rect 2498 4564 2504 4576
rect 2556 4564 2562 4616
rect 3694 4564 3700 4616
rect 3752 4604 3758 4616
rect 3973 4607 4031 4613
rect 3973 4604 3985 4607
rect 3752 4576 3985 4604
rect 3752 4564 3758 4576
rect 3973 4573 3985 4576
rect 4019 4573 4031 4607
rect 3973 4567 4031 4573
rect 4801 4607 4859 4613
rect 4801 4573 4813 4607
rect 4847 4604 4859 4607
rect 5261 4607 5319 4613
rect 5261 4604 5273 4607
rect 4847 4576 5273 4604
rect 4847 4573 4859 4576
rect 4801 4567 4859 4573
rect 5261 4573 5273 4576
rect 5307 4573 5319 4607
rect 5261 4567 5319 4573
rect 28350 4564 28356 4616
rect 28408 4604 28414 4616
rect 28408 4576 28453 4604
rect 28408 4564 28414 4576
rect 22097 4539 22155 4545
rect 22097 4505 22109 4539
rect 22143 4536 22155 4539
rect 22186 4536 22192 4548
rect 22143 4508 22192 4536
rect 22143 4505 22155 4508
rect 22097 4499 22155 4505
rect 22186 4496 22192 4508
rect 22244 4496 22250 4548
rect 23750 4536 23756 4548
rect 23711 4508 23756 4536
rect 23750 4496 23756 4508
rect 23808 4496 23814 4548
rect 28166 4536 28172 4548
rect 28127 4508 28172 4536
rect 28166 4496 28172 4508
rect 28224 4496 28230 4548
rect 1946 4428 1952 4480
rect 2004 4468 2010 4480
rect 2317 4471 2375 4477
rect 2317 4468 2329 4471
rect 2004 4440 2329 4468
rect 2004 4428 2010 4440
rect 2317 4437 2329 4440
rect 2363 4437 2375 4471
rect 2317 4431 2375 4437
rect 1104 4378 29048 4400
rect 1104 4326 7896 4378
rect 7948 4326 7960 4378
rect 8012 4326 8024 4378
rect 8076 4326 8088 4378
rect 8140 4326 8152 4378
rect 8204 4326 14842 4378
rect 14894 4326 14906 4378
rect 14958 4326 14970 4378
rect 15022 4326 15034 4378
rect 15086 4326 15098 4378
rect 15150 4326 21788 4378
rect 21840 4326 21852 4378
rect 21904 4326 21916 4378
rect 21968 4326 21980 4378
rect 22032 4326 22044 4378
rect 22096 4326 28734 4378
rect 28786 4326 28798 4378
rect 28850 4326 28862 4378
rect 28914 4326 28926 4378
rect 28978 4326 28990 4378
rect 29042 4326 29048 4378
rect 1104 4304 29048 4326
rect 2498 4264 2504 4276
rect 1964 4236 2504 4264
rect 1964 4137 1992 4236
rect 2498 4224 2504 4236
rect 2556 4264 2562 4276
rect 4430 4264 4436 4276
rect 2556 4236 4436 4264
rect 2556 4224 2562 4236
rect 4430 4224 4436 4236
rect 4488 4224 4494 4276
rect 27801 4267 27859 4273
rect 27801 4233 27813 4267
rect 27847 4264 27859 4267
rect 28166 4264 28172 4276
rect 27847 4236 28172 4264
rect 27847 4233 27859 4236
rect 27801 4227 27859 4233
rect 28166 4224 28172 4236
rect 28224 4224 28230 4276
rect 3528 4168 5120 4196
rect 1949 4131 2007 4137
rect 1949 4097 1961 4131
rect 1995 4097 2007 4131
rect 2406 4128 2412 4140
rect 2367 4100 2412 4128
rect 1949 4091 2007 4097
rect 2406 4088 2412 4100
rect 2464 4088 2470 4140
rect 2501 4131 2559 4137
rect 2501 4097 2513 4131
rect 2547 4128 2559 4131
rect 3142 4128 3148 4140
rect 2547 4100 3148 4128
rect 2547 4097 2559 4100
rect 2501 4091 2559 4097
rect 3142 4088 3148 4100
rect 3200 4088 3206 4140
rect 3234 4088 3240 4140
rect 3292 4128 3298 4140
rect 3292 4100 3337 4128
rect 3292 4088 3298 4100
rect 2424 4060 2452 4088
rect 3528 4060 3556 4168
rect 3694 4128 3700 4140
rect 3655 4100 3700 4128
rect 3694 4088 3700 4100
rect 3752 4088 3758 4140
rect 5092 4128 5120 4168
rect 6733 4131 6791 4137
rect 6733 4128 6745 4131
rect 5092 4100 6745 4128
rect 6733 4097 6745 4100
rect 6779 4128 6791 4131
rect 10502 4128 10508 4140
rect 6779 4100 6914 4128
rect 10463 4100 10508 4128
rect 6779 4097 6791 4100
rect 6733 4091 6791 4097
rect 2424 4032 3556 4060
rect 3881 4063 3939 4069
rect 3881 4029 3893 4063
rect 3927 4060 3939 4063
rect 4246 4060 4252 4072
rect 3927 4032 4252 4060
rect 3927 4029 3939 4032
rect 3881 4023 3939 4029
rect 4246 4020 4252 4032
rect 4304 4020 4310 4072
rect 4341 4063 4399 4069
rect 4341 4029 4353 4063
rect 4387 4029 4399 4063
rect 6886 4060 6914 4100
rect 10502 4088 10508 4100
rect 10560 4088 10566 4140
rect 18693 4131 18751 4137
rect 18693 4097 18705 4131
rect 18739 4097 18751 4131
rect 18693 4091 18751 4097
rect 11790 4060 11796 4072
rect 6886 4032 11796 4060
rect 4341 4023 4399 4029
rect 2866 3952 2872 4004
rect 2924 3992 2930 4004
rect 4356 3992 4384 4023
rect 11790 4020 11796 4032
rect 11848 4020 11854 4072
rect 12802 4060 12808 4072
rect 12763 4032 12808 4060
rect 12802 4020 12808 4032
rect 12860 4020 12866 4072
rect 12986 4060 12992 4072
rect 12947 4032 12992 4060
rect 12986 4020 12992 4032
rect 13044 4020 13050 4072
rect 13630 4060 13636 4072
rect 13591 4032 13636 4060
rect 13630 4020 13636 4032
rect 13688 4020 13694 4072
rect 2924 3964 4384 3992
rect 2924 3952 2930 3964
rect 4430 3952 4436 4004
rect 4488 3992 4494 4004
rect 18138 3992 18144 4004
rect 4488 3964 18144 3992
rect 4488 3952 4494 3964
rect 18138 3952 18144 3964
rect 18196 3952 18202 4004
rect 18708 3992 18736 4091
rect 21174 4088 21180 4140
rect 21232 4128 21238 4140
rect 21269 4131 21327 4137
rect 21269 4128 21281 4131
rect 21232 4100 21281 4128
rect 21232 4088 21238 4100
rect 21269 4097 21281 4100
rect 21315 4097 21327 4131
rect 21269 4091 21327 4097
rect 21284 4060 21312 4091
rect 22094 4088 22100 4140
rect 22152 4128 22158 4140
rect 22189 4131 22247 4137
rect 22189 4128 22201 4131
rect 22152 4100 22201 4128
rect 22152 4088 22158 4100
rect 22189 4097 22201 4100
rect 22235 4097 22247 4131
rect 22189 4091 22247 4097
rect 22281 4131 22339 4137
rect 22281 4097 22293 4131
rect 22327 4128 22339 4131
rect 23750 4128 23756 4140
rect 22327 4100 23756 4128
rect 22327 4097 22339 4100
rect 22281 4091 22339 4097
rect 23750 4088 23756 4100
rect 23808 4088 23814 4140
rect 27706 4128 27712 4140
rect 27667 4100 27712 4128
rect 27706 4088 27712 4100
rect 27764 4088 27770 4140
rect 24946 4060 24952 4072
rect 21284 4032 24952 4060
rect 24946 4020 24952 4032
rect 25004 4020 25010 4072
rect 18708 3964 22094 3992
rect 1762 3884 1768 3936
rect 1820 3924 1826 3936
rect 1857 3927 1915 3933
rect 1857 3924 1869 3927
rect 1820 3896 1869 3924
rect 1820 3884 1826 3896
rect 1857 3893 1869 3896
rect 1903 3893 1915 3927
rect 1857 3887 1915 3893
rect 3145 3927 3203 3933
rect 3145 3893 3157 3927
rect 3191 3924 3203 3927
rect 4338 3924 4344 3936
rect 3191 3896 4344 3924
rect 3191 3893 3203 3896
rect 3145 3887 3203 3893
rect 4338 3884 4344 3896
rect 4396 3884 4402 3936
rect 5902 3884 5908 3936
rect 5960 3924 5966 3936
rect 6641 3927 6699 3933
rect 6641 3924 6653 3927
rect 5960 3896 6653 3924
rect 5960 3884 5966 3896
rect 6641 3893 6653 3896
rect 6687 3893 6699 3927
rect 6641 3887 6699 3893
rect 6914 3884 6920 3936
rect 6972 3924 6978 3936
rect 7745 3927 7803 3933
rect 7745 3924 7757 3927
rect 6972 3896 7757 3924
rect 6972 3884 6978 3896
rect 7745 3893 7757 3896
rect 7791 3893 7803 3927
rect 10594 3924 10600 3936
rect 10555 3896 10600 3924
rect 7745 3887 7803 3893
rect 10594 3884 10600 3896
rect 10652 3884 10658 3936
rect 18785 3927 18843 3933
rect 18785 3893 18797 3927
rect 18831 3924 18843 3927
rect 19610 3924 19616 3936
rect 18831 3896 19616 3924
rect 18831 3893 18843 3896
rect 18785 3887 18843 3893
rect 19610 3884 19616 3896
rect 19668 3884 19674 3936
rect 20346 3884 20352 3936
rect 20404 3924 20410 3936
rect 20441 3927 20499 3933
rect 20441 3924 20453 3927
rect 20404 3896 20453 3924
rect 20404 3884 20410 3896
rect 20441 3893 20453 3896
rect 20487 3893 20499 3927
rect 20441 3887 20499 3893
rect 20530 3884 20536 3936
rect 20588 3924 20594 3936
rect 21177 3927 21235 3933
rect 21177 3924 21189 3927
rect 20588 3896 21189 3924
rect 20588 3884 20594 3896
rect 21177 3893 21189 3896
rect 21223 3893 21235 3927
rect 22066 3924 22094 3964
rect 27614 3924 27620 3936
rect 22066 3896 27620 3924
rect 21177 3887 21235 3893
rect 27614 3884 27620 3896
rect 27672 3884 27678 3936
rect 1104 3834 28888 3856
rect 1104 3782 4423 3834
rect 4475 3782 4487 3834
rect 4539 3782 4551 3834
rect 4603 3782 4615 3834
rect 4667 3782 4679 3834
rect 4731 3782 11369 3834
rect 11421 3782 11433 3834
rect 11485 3782 11497 3834
rect 11549 3782 11561 3834
rect 11613 3782 11625 3834
rect 11677 3782 18315 3834
rect 18367 3782 18379 3834
rect 18431 3782 18443 3834
rect 18495 3782 18507 3834
rect 18559 3782 18571 3834
rect 18623 3782 25261 3834
rect 25313 3782 25325 3834
rect 25377 3782 25389 3834
rect 25441 3782 25453 3834
rect 25505 3782 25517 3834
rect 25569 3782 28888 3834
rect 1104 3760 28888 3782
rect 4246 3720 4252 3732
rect 4207 3692 4252 3720
rect 4246 3680 4252 3692
rect 4304 3680 4310 3732
rect 12802 3680 12808 3732
rect 12860 3720 12866 3732
rect 12897 3723 12955 3729
rect 12897 3720 12909 3723
rect 12860 3692 12909 3720
rect 12860 3680 12866 3692
rect 12897 3689 12909 3692
rect 12943 3689 12955 3723
rect 12897 3683 12955 3689
rect 658 3612 664 3664
rect 716 3652 722 3664
rect 716 3624 2084 3652
rect 716 3612 722 3624
rect 1578 3584 1584 3596
rect 1539 3556 1584 3584
rect 1578 3544 1584 3556
rect 1636 3544 1642 3596
rect 1762 3584 1768 3596
rect 1723 3556 1768 3584
rect 1762 3544 1768 3556
rect 1820 3544 1826 3596
rect 2056 3593 2084 3624
rect 3878 3612 3884 3664
rect 3936 3652 3942 3664
rect 5534 3652 5540 3664
rect 3936 3624 5540 3652
rect 3936 3612 3942 3624
rect 5534 3612 5540 3624
rect 5592 3612 5598 3664
rect 21174 3652 21180 3664
rect 8220 3624 21180 3652
rect 2041 3587 2099 3593
rect 2041 3553 2053 3587
rect 2087 3553 2099 3587
rect 5902 3584 5908 3596
rect 5863 3556 5908 3584
rect 2041 3547 2099 3553
rect 5902 3544 5908 3556
rect 5960 3544 5966 3596
rect 6454 3584 6460 3596
rect 6415 3556 6460 3584
rect 6454 3544 6460 3556
rect 6512 3544 6518 3596
rect 3234 3476 3240 3528
rect 3292 3516 3298 3528
rect 8220 3525 8248 3624
rect 21174 3612 21180 3624
rect 21232 3612 21238 3664
rect 10594 3584 10600 3596
rect 10555 3556 10600 3584
rect 10594 3544 10600 3556
rect 10652 3544 10658 3596
rect 10962 3584 10968 3596
rect 10923 3556 10968 3584
rect 10962 3544 10968 3556
rect 11020 3544 11026 3596
rect 11790 3544 11796 3596
rect 11848 3584 11854 3596
rect 20346 3584 20352 3596
rect 11848 3556 16574 3584
rect 11848 3544 11854 3556
rect 4341 3519 4399 3525
rect 4341 3516 4353 3519
rect 3292 3488 4353 3516
rect 3292 3476 3298 3488
rect 4341 3485 4353 3488
rect 4387 3485 4399 3519
rect 4341 3479 4399 3485
rect 5261 3519 5319 3525
rect 5261 3485 5273 3519
rect 5307 3516 5319 3519
rect 5721 3519 5779 3525
rect 5721 3516 5733 3519
rect 5307 3488 5733 3516
rect 5307 3485 5319 3488
rect 5261 3479 5319 3485
rect 5721 3485 5733 3488
rect 5767 3485 5779 3519
rect 5721 3479 5779 3485
rect 8205 3519 8263 3525
rect 8205 3485 8217 3519
rect 8251 3485 8263 3519
rect 8205 3479 8263 3485
rect 4356 3448 4384 3479
rect 8220 3448 8248 3479
rect 9214 3476 9220 3528
rect 9272 3516 9278 3528
rect 9309 3519 9367 3525
rect 9309 3516 9321 3519
rect 9272 3488 9321 3516
rect 9272 3476 9278 3488
rect 9309 3485 9321 3488
rect 9355 3485 9367 3519
rect 9309 3479 9367 3485
rect 9953 3519 10011 3525
rect 9953 3485 9965 3519
rect 9999 3516 10011 3519
rect 10413 3519 10471 3525
rect 10413 3516 10425 3519
rect 9999 3488 10425 3516
rect 9999 3485 10011 3488
rect 9953 3479 10011 3485
rect 10413 3485 10425 3488
rect 10459 3485 10471 3519
rect 13538 3516 13544 3528
rect 13499 3488 13544 3516
rect 10413 3479 10471 3485
rect 13538 3476 13544 3488
rect 13596 3476 13602 3528
rect 13998 3476 14004 3528
rect 14056 3516 14062 3528
rect 14277 3519 14335 3525
rect 14277 3516 14289 3519
rect 14056 3488 14289 3516
rect 14056 3476 14062 3488
rect 14277 3485 14289 3488
rect 14323 3485 14335 3519
rect 16206 3516 16212 3528
rect 16167 3488 16212 3516
rect 14277 3479 14335 3485
rect 16206 3476 16212 3488
rect 16264 3476 16270 3528
rect 16546 3516 16574 3556
rect 16684 3556 19288 3584
rect 20307 3556 20352 3584
rect 16684 3525 16712 3556
rect 16669 3519 16727 3525
rect 16669 3516 16681 3519
rect 16546 3488 16681 3516
rect 16669 3485 16681 3488
rect 16715 3485 16727 3519
rect 16669 3479 16727 3485
rect 17681 3519 17739 3525
rect 17681 3485 17693 3519
rect 17727 3485 17739 3519
rect 18138 3516 18144 3528
rect 18099 3488 18144 3516
rect 17681 3479 17739 3485
rect 4356 3420 8248 3448
rect 17696 3448 17724 3479
rect 18138 3476 18144 3488
rect 18196 3476 18202 3528
rect 19150 3448 19156 3460
rect 17696 3420 19156 3448
rect 19150 3408 19156 3420
rect 19208 3408 19214 3460
rect 19260 3448 19288 3556
rect 20346 3544 20352 3556
rect 20404 3544 20410 3596
rect 20530 3584 20536 3596
rect 20491 3556 20536 3584
rect 20530 3544 20536 3556
rect 20588 3544 20594 3596
rect 21266 3584 21272 3596
rect 21227 3556 21272 3584
rect 21266 3544 21272 3556
rect 21324 3544 21330 3596
rect 27522 3584 27528 3596
rect 27483 3556 27528 3584
rect 27522 3544 27528 3556
rect 27580 3544 27586 3596
rect 19426 3516 19432 3528
rect 19387 3488 19432 3516
rect 19426 3476 19432 3488
rect 19484 3476 19490 3528
rect 26053 3519 26111 3525
rect 26053 3485 26065 3519
rect 26099 3516 26111 3519
rect 26513 3519 26571 3525
rect 26513 3516 26525 3519
rect 26099 3488 26525 3516
rect 26099 3485 26111 3488
rect 26053 3479 26111 3485
rect 26513 3485 26525 3488
rect 26559 3485 26571 3519
rect 26513 3479 26571 3485
rect 22094 3448 22100 3460
rect 19260 3420 22100 3448
rect 22094 3408 22100 3420
rect 22152 3448 22158 3460
rect 23842 3448 23848 3460
rect 22152 3420 23848 3448
rect 22152 3408 22158 3420
rect 23842 3408 23848 3420
rect 23900 3408 23906 3460
rect 26697 3451 26755 3457
rect 26697 3417 26709 3451
rect 26743 3448 26755 3451
rect 27246 3448 27252 3460
rect 26743 3420 27252 3448
rect 26743 3417 26755 3420
rect 26697 3411 26755 3417
rect 27246 3408 27252 3420
rect 27304 3408 27310 3460
rect 7098 3340 7104 3392
rect 7156 3380 7162 3392
rect 8113 3383 8171 3389
rect 8113 3380 8125 3383
rect 7156 3352 8125 3380
rect 7156 3340 7162 3352
rect 8113 3349 8125 3352
rect 8159 3349 8171 3383
rect 8113 3343 8171 3349
rect 13633 3383 13691 3389
rect 13633 3349 13645 3383
rect 13679 3380 13691 3383
rect 14182 3380 14188 3392
rect 13679 3352 14188 3380
rect 13679 3349 13691 3352
rect 13633 3343 13691 3349
rect 14182 3340 14188 3352
rect 14240 3340 14246 3392
rect 16761 3383 16819 3389
rect 16761 3349 16773 3383
rect 16807 3380 16819 3383
rect 17034 3380 17040 3392
rect 16807 3352 17040 3380
rect 16807 3349 16819 3352
rect 16761 3343 16819 3349
rect 17034 3340 17040 3352
rect 17092 3340 17098 3392
rect 18233 3383 18291 3389
rect 18233 3349 18245 3383
rect 18279 3380 18291 3383
rect 19334 3380 19340 3392
rect 18279 3352 19340 3380
rect 18279 3349 18291 3352
rect 18233 3343 18291 3349
rect 19334 3340 19340 3352
rect 19392 3340 19398 3392
rect 1104 3290 29048 3312
rect 1104 3238 7896 3290
rect 7948 3238 7960 3290
rect 8012 3238 8024 3290
rect 8076 3238 8088 3290
rect 8140 3238 8152 3290
rect 8204 3238 14842 3290
rect 14894 3238 14906 3290
rect 14958 3238 14970 3290
rect 15022 3238 15034 3290
rect 15086 3238 15098 3290
rect 15150 3238 21788 3290
rect 21840 3238 21852 3290
rect 21904 3238 21916 3290
rect 21968 3238 21980 3290
rect 22032 3238 22044 3290
rect 22096 3238 28734 3290
rect 28786 3238 28798 3290
rect 28850 3238 28862 3290
rect 28914 3238 28926 3290
rect 28978 3238 28990 3290
rect 29042 3238 29048 3290
rect 1104 3216 29048 3238
rect 2682 3136 2688 3188
rect 2740 3176 2746 3188
rect 4798 3176 4804 3188
rect 2740 3148 4804 3176
rect 2740 3136 2746 3148
rect 4798 3136 4804 3148
rect 4856 3136 4862 3188
rect 12897 3179 12955 3185
rect 12897 3145 12909 3179
rect 12943 3176 12955 3179
rect 12986 3176 12992 3188
rect 12943 3148 12992 3176
rect 12943 3145 12955 3148
rect 12897 3139 12955 3145
rect 12986 3136 12992 3148
rect 13044 3136 13050 3188
rect 27246 3176 27252 3188
rect 27207 3148 27252 3176
rect 27246 3136 27252 3148
rect 27304 3136 27310 3188
rect 1946 3108 1952 3120
rect 1907 3080 1952 3108
rect 1946 3068 1952 3080
rect 2004 3068 2010 3120
rect 4338 3108 4344 3120
rect 4299 3080 4344 3108
rect 4338 3068 4344 3080
rect 4396 3068 4402 3120
rect 7098 3108 7104 3120
rect 7059 3080 7104 3108
rect 7098 3068 7104 3080
rect 7156 3068 7162 3120
rect 9398 3108 9404 3120
rect 9359 3080 9404 3108
rect 9398 3068 9404 3080
rect 9456 3068 9462 3120
rect 14182 3108 14188 3120
rect 14143 3080 14188 3108
rect 14182 3068 14188 3080
rect 14240 3068 14246 3120
rect 17034 3108 17040 3120
rect 16995 3080 17040 3108
rect 17034 3068 17040 3080
rect 17092 3068 17098 3120
rect 19334 3108 19340 3120
rect 19295 3080 19340 3108
rect 19334 3068 19340 3080
rect 19392 3068 19398 3120
rect 26421 3111 26479 3117
rect 26421 3077 26433 3111
rect 26467 3108 26479 3111
rect 27798 3108 27804 3120
rect 26467 3080 27804 3108
rect 26467 3077 26479 3080
rect 26421 3071 26479 3077
rect 27798 3068 27804 3080
rect 27856 3068 27862 3120
rect 4154 3040 4160 3052
rect 4115 3012 4160 3040
rect 4154 3000 4160 3012
rect 4212 3000 4218 3052
rect 9214 3040 9220 3052
rect 9175 3012 9220 3040
rect 9214 3000 9220 3012
rect 9272 3000 9278 3052
rect 12805 3043 12863 3049
rect 12805 3009 12817 3043
rect 12851 3040 12863 3043
rect 13538 3040 13544 3052
rect 12851 3012 13544 3040
rect 12851 3009 12863 3012
rect 12805 3003 12863 3009
rect 13538 3000 13544 3012
rect 13596 3000 13602 3052
rect 13998 3040 14004 3052
rect 13959 3012 14004 3040
rect 13998 3000 14004 3012
rect 14056 3000 14062 3052
rect 16206 3000 16212 3052
rect 16264 3040 16270 3052
rect 16853 3043 16911 3049
rect 16853 3040 16865 3043
rect 16264 3012 16865 3040
rect 16264 3000 16270 3012
rect 16853 3009 16865 3012
rect 16899 3009 16911 3043
rect 19150 3040 19156 3052
rect 19111 3012 19156 3040
rect 16853 3003 16911 3009
rect 19150 3000 19156 3012
rect 19208 3000 19214 3052
rect 26602 3000 26608 3052
rect 26660 3040 26666 3052
rect 27341 3043 27399 3049
rect 26660 3012 26705 3040
rect 26660 3000 26666 3012
rect 27341 3009 27353 3043
rect 27387 3040 27399 3043
rect 27614 3040 27620 3052
rect 27387 3012 27620 3040
rect 27387 3009 27399 3012
rect 27341 3003 27399 3009
rect 27614 3000 27620 3012
rect 27672 3000 27678 3052
rect 28077 3043 28135 3049
rect 28077 3009 28089 3043
rect 28123 3040 28135 3043
rect 28350 3040 28356 3052
rect 28123 3012 28356 3040
rect 28123 3009 28135 3012
rect 28077 3003 28135 3009
rect 28350 3000 28356 3012
rect 28408 3000 28414 3052
rect 1762 2972 1768 2984
rect 1723 2944 1768 2972
rect 1762 2932 1768 2944
rect 1820 2932 1826 2984
rect 2774 2972 2780 2984
rect 2735 2944 2780 2972
rect 2774 2932 2780 2944
rect 2832 2932 2838 2984
rect 4798 2972 4804 2984
rect 4759 2944 4804 2972
rect 4798 2932 4804 2944
rect 4856 2932 4862 2984
rect 6914 2932 6920 2984
rect 6972 2972 6978 2984
rect 8386 2972 8392 2984
rect 6972 2944 7017 2972
rect 8347 2944 8392 2972
rect 6972 2932 6978 2944
rect 8386 2932 8392 2944
rect 8444 2932 8450 2984
rect 9674 2972 9680 2984
rect 9635 2944 9680 2972
rect 9674 2932 9680 2944
rect 9732 2932 9738 2984
rect 14734 2972 14740 2984
rect 14695 2944 14740 2972
rect 14734 2932 14740 2944
rect 14792 2932 14798 2984
rect 16758 2932 16764 2984
rect 16816 2972 16822 2984
rect 17313 2975 17371 2981
rect 17313 2972 17325 2975
rect 16816 2944 17325 2972
rect 16816 2932 16822 2944
rect 17313 2941 17325 2944
rect 17359 2941 17371 2975
rect 17313 2935 17371 2941
rect 19613 2975 19671 2981
rect 19613 2941 19625 2975
rect 19659 2941 19671 2975
rect 26142 2972 26148 2984
rect 26103 2944 26148 2972
rect 19613 2935 19671 2941
rect 18046 2864 18052 2916
rect 18104 2904 18110 2916
rect 19628 2904 19656 2935
rect 26142 2932 26148 2944
rect 26200 2932 26206 2984
rect 18104 2876 19656 2904
rect 18104 2864 18110 2876
rect 1104 2746 28888 2768
rect 1104 2694 4423 2746
rect 4475 2694 4487 2746
rect 4539 2694 4551 2746
rect 4603 2694 4615 2746
rect 4667 2694 4679 2746
rect 4731 2694 11369 2746
rect 11421 2694 11433 2746
rect 11485 2694 11497 2746
rect 11549 2694 11561 2746
rect 11613 2694 11625 2746
rect 11677 2694 18315 2746
rect 18367 2694 18379 2746
rect 18431 2694 18443 2746
rect 18495 2694 18507 2746
rect 18559 2694 18571 2746
rect 18623 2694 25261 2746
rect 25313 2694 25325 2746
rect 25377 2694 25389 2746
rect 25441 2694 25453 2746
rect 25505 2694 25517 2746
rect 25569 2694 28888 2746
rect 1104 2672 28888 2694
rect 1762 2592 1768 2644
rect 1820 2632 1826 2644
rect 1857 2635 1915 2641
rect 1857 2632 1869 2635
rect 1820 2604 1869 2632
rect 1820 2592 1826 2604
rect 1857 2601 1869 2604
rect 1903 2601 1915 2635
rect 17586 2632 17592 2644
rect 17547 2604 17592 2632
rect 1857 2595 1915 2601
rect 17586 2592 17592 2604
rect 17644 2592 17650 2644
rect 25866 2592 25872 2644
rect 25924 2632 25930 2644
rect 26421 2635 26479 2641
rect 26421 2632 26433 2635
rect 25924 2604 26433 2632
rect 25924 2592 25930 2604
rect 26421 2601 26433 2604
rect 26467 2601 26479 2635
rect 27798 2632 27804 2644
rect 27759 2604 27804 2632
rect 26421 2595 26479 2601
rect 27798 2592 27804 2604
rect 27856 2592 27862 2644
rect 15838 2524 15844 2576
rect 15896 2564 15902 2576
rect 16853 2567 16911 2573
rect 16853 2564 16865 2567
rect 15896 2536 16865 2564
rect 15896 2524 15902 2536
rect 16853 2533 16865 2536
rect 16899 2533 16911 2567
rect 16853 2527 16911 2533
rect 3234 2456 3240 2508
rect 3292 2496 3298 2508
rect 4433 2499 4491 2505
rect 4433 2496 4445 2499
rect 3292 2468 4445 2496
rect 3292 2456 3298 2468
rect 4433 2465 4445 2468
rect 4479 2465 4491 2499
rect 4433 2459 4491 2465
rect 9401 2499 9459 2505
rect 9401 2465 9413 2499
rect 9447 2496 9459 2499
rect 9490 2496 9496 2508
rect 9447 2468 9496 2496
rect 9447 2465 9459 2468
rect 9401 2459 9459 2465
rect 9490 2456 9496 2468
rect 9548 2456 9554 2508
rect 19426 2496 19432 2508
rect 19387 2468 19432 2496
rect 19426 2456 19432 2468
rect 19484 2456 19490 2508
rect 19610 2496 19616 2508
rect 19571 2468 19616 2496
rect 19610 2456 19616 2468
rect 19668 2456 19674 2508
rect 19978 2496 19984 2508
rect 19939 2468 19984 2496
rect 19978 2456 19984 2468
rect 20036 2456 20042 2508
rect 2590 2428 2596 2440
rect 2551 2400 2596 2428
rect 2590 2388 2596 2400
rect 2648 2388 2654 2440
rect 3421 2431 3479 2437
rect 3421 2397 3433 2431
rect 3467 2428 3479 2431
rect 3973 2431 4031 2437
rect 3973 2428 3985 2431
rect 3467 2400 3985 2428
rect 3467 2397 3479 2400
rect 3421 2391 3479 2397
rect 3973 2397 3985 2400
rect 4019 2397 4031 2431
rect 3973 2391 4031 2397
rect 9030 2388 9036 2440
rect 9088 2428 9094 2440
rect 9125 2431 9183 2437
rect 9125 2428 9137 2431
rect 9088 2400 9137 2428
rect 9088 2388 9094 2400
rect 9125 2397 9137 2400
rect 9171 2397 9183 2431
rect 9125 2391 9183 2397
rect 17402 2388 17408 2440
rect 17460 2428 17466 2440
rect 17773 2431 17831 2437
rect 17773 2428 17785 2431
rect 17460 2400 17785 2428
rect 17460 2388 17466 2400
rect 17773 2397 17785 2400
rect 17819 2397 17831 2431
rect 17773 2391 17831 2397
rect 26605 2431 26663 2437
rect 26605 2397 26617 2431
rect 26651 2428 26663 2431
rect 27062 2428 27068 2440
rect 26651 2400 27068 2428
rect 26651 2397 26663 2400
rect 26605 2391 26663 2397
rect 27062 2388 27068 2400
rect 27120 2388 27126 2440
rect 27614 2388 27620 2440
rect 27672 2428 27678 2440
rect 27709 2431 27767 2437
rect 27709 2428 27721 2431
rect 27672 2400 27721 2428
rect 27672 2388 27678 2400
rect 27709 2397 27721 2400
rect 27755 2397 27767 2431
rect 27709 2391 27767 2397
rect 2685 2363 2743 2369
rect 2685 2329 2697 2363
rect 2731 2360 2743 2363
rect 4157 2363 4215 2369
rect 4157 2360 4169 2363
rect 2731 2332 4169 2360
rect 2731 2329 2743 2332
rect 2685 2323 2743 2329
rect 4157 2329 4169 2332
rect 4203 2329 4215 2363
rect 4157 2323 4215 2329
rect 16114 2320 16120 2372
rect 16172 2360 16178 2372
rect 17037 2363 17095 2369
rect 17037 2360 17049 2363
rect 16172 2332 17049 2360
rect 16172 2320 16178 2332
rect 17037 2329 17049 2332
rect 17083 2329 17095 2363
rect 17037 2323 17095 2329
rect 3510 2252 3516 2304
rect 3568 2292 3574 2304
rect 8294 2292 8300 2304
rect 3568 2264 8300 2292
rect 3568 2252 3574 2264
rect 8294 2252 8300 2264
rect 8352 2252 8358 2304
rect 1104 2202 29048 2224
rect 1104 2150 7896 2202
rect 7948 2150 7960 2202
rect 8012 2150 8024 2202
rect 8076 2150 8088 2202
rect 8140 2150 8152 2202
rect 8204 2150 14842 2202
rect 14894 2150 14906 2202
rect 14958 2150 14970 2202
rect 15022 2150 15034 2202
rect 15086 2150 15098 2202
rect 15150 2150 21788 2202
rect 21840 2150 21852 2202
rect 21904 2150 21916 2202
rect 21968 2150 21980 2202
rect 22032 2150 22044 2202
rect 22096 2150 28734 2202
rect 28786 2150 28798 2202
rect 28850 2150 28862 2202
rect 28914 2150 28926 2202
rect 28978 2150 28990 2202
rect 29042 2150 29048 2202
rect 1104 2128 29048 2150
<< via1 >>
rect 4423 47302 4475 47354
rect 4487 47302 4539 47354
rect 4551 47302 4603 47354
rect 4615 47302 4667 47354
rect 4679 47302 4731 47354
rect 11369 47302 11421 47354
rect 11433 47302 11485 47354
rect 11497 47302 11549 47354
rect 11561 47302 11613 47354
rect 11625 47302 11677 47354
rect 18315 47302 18367 47354
rect 18379 47302 18431 47354
rect 18443 47302 18495 47354
rect 18507 47302 18559 47354
rect 18571 47302 18623 47354
rect 25261 47302 25313 47354
rect 25325 47302 25377 47354
rect 25389 47302 25441 47354
rect 25453 47302 25505 47354
rect 25517 47302 25569 47354
rect 23756 47132 23808 47184
rect 25044 47132 25096 47184
rect 10324 47107 10376 47116
rect 10324 47073 10333 47107
rect 10333 47073 10367 47107
rect 10367 47073 10376 47107
rect 10324 47064 10376 47073
rect 28356 47064 28408 47116
rect 2228 47039 2280 47048
rect 2228 47005 2237 47039
rect 2237 47005 2271 47039
rect 2271 47005 2280 47039
rect 2228 46996 2280 47005
rect 2872 47039 2924 47048
rect 2872 47005 2881 47039
rect 2881 47005 2915 47039
rect 2915 47005 2924 47039
rect 5816 47039 5868 47048
rect 2872 46996 2924 47005
rect 5816 47005 5825 47039
rect 5825 47005 5859 47039
rect 5859 47005 5868 47039
rect 5816 46996 5868 47005
rect 6460 46996 6512 47048
rect 7012 46996 7064 47048
rect 9312 47039 9364 47048
rect 9312 47005 9321 47039
rect 9321 47005 9355 47039
rect 9355 47005 9364 47039
rect 9312 46996 9364 47005
rect 12900 46996 12952 47048
rect 18236 46996 18288 47048
rect 22836 46996 22888 47048
rect 24032 47039 24084 47048
rect 24032 47005 24041 47039
rect 24041 47005 24075 47039
rect 24075 47005 24084 47039
rect 24032 46996 24084 47005
rect 26608 47039 26660 47048
rect 26608 47005 26617 47039
rect 26617 47005 26651 47039
rect 26651 47005 26660 47039
rect 26608 46996 26660 47005
rect 27344 46996 27396 47048
rect 27896 47039 27948 47048
rect 27896 47005 27905 47039
rect 27905 47005 27939 47039
rect 27939 47005 27948 47039
rect 27896 46996 27948 47005
rect 9220 46928 9272 46980
rect 9496 46971 9548 46980
rect 9496 46937 9505 46971
rect 9505 46937 9539 46971
rect 9539 46937 9548 46971
rect 9496 46928 9548 46937
rect 26424 46971 26476 46980
rect 26424 46937 26433 46971
rect 26433 46937 26467 46971
rect 26467 46937 26476 46971
rect 26424 46928 26476 46937
rect 2780 46903 2832 46912
rect 2780 46869 2789 46903
rect 2789 46869 2823 46903
rect 2823 46869 2832 46903
rect 2780 46860 2832 46869
rect 6000 46903 6052 46912
rect 6000 46869 6009 46903
rect 6009 46869 6043 46903
rect 6043 46869 6052 46903
rect 6000 46860 6052 46869
rect 6736 46903 6788 46912
rect 6736 46869 6745 46903
rect 6745 46869 6779 46903
rect 6779 46869 6788 46903
rect 6736 46860 6788 46869
rect 19984 46860 20036 46912
rect 23480 46860 23532 46912
rect 7896 46758 7948 46810
rect 7960 46758 8012 46810
rect 8024 46758 8076 46810
rect 8088 46758 8140 46810
rect 8152 46758 8204 46810
rect 14842 46758 14894 46810
rect 14906 46758 14958 46810
rect 14970 46758 15022 46810
rect 15034 46758 15086 46810
rect 15098 46758 15150 46810
rect 21788 46758 21840 46810
rect 21852 46758 21904 46810
rect 21916 46758 21968 46810
rect 21980 46758 22032 46810
rect 22044 46758 22096 46810
rect 28734 46758 28786 46810
rect 28798 46758 28850 46810
rect 28862 46758 28914 46810
rect 28926 46758 28978 46810
rect 28990 46758 29042 46810
rect 26424 46699 26476 46708
rect 26424 46665 26433 46699
rect 26433 46665 26467 46699
rect 26467 46665 26476 46699
rect 26424 46656 26476 46665
rect 2780 46588 2832 46640
rect 2228 46520 2280 46572
rect 7012 46563 7064 46572
rect 7012 46529 7021 46563
rect 7021 46529 7055 46563
rect 7055 46529 7064 46563
rect 7012 46520 7064 46529
rect 12900 46563 12952 46572
rect 12900 46529 12909 46563
rect 12909 46529 12943 46563
rect 12943 46529 12952 46563
rect 12900 46520 12952 46529
rect 15844 46563 15896 46572
rect 15844 46529 15853 46563
rect 15853 46529 15887 46563
rect 15887 46529 15896 46563
rect 15844 46520 15896 46529
rect 18236 46563 18288 46572
rect 18236 46529 18245 46563
rect 18245 46529 18279 46563
rect 18279 46529 18288 46563
rect 18236 46520 18288 46529
rect 22836 46563 22888 46572
rect 22836 46529 22845 46563
rect 22845 46529 22879 46563
rect 22879 46529 22888 46563
rect 22836 46520 22888 46529
rect 1952 46452 2004 46504
rect 7932 46452 7984 46504
rect 8392 46495 8444 46504
rect 8392 46461 8401 46495
rect 8401 46461 8435 46495
rect 8435 46461 8444 46495
rect 8392 46452 8444 46461
rect 10140 46452 10192 46504
rect 10968 46495 11020 46504
rect 10968 46461 10977 46495
rect 10977 46461 11011 46495
rect 11011 46461 11020 46495
rect 10968 46452 11020 46461
rect 13084 46495 13136 46504
rect 13084 46461 13093 46495
rect 13093 46461 13127 46495
rect 13127 46461 13136 46495
rect 13084 46452 13136 46461
rect 13544 46495 13596 46504
rect 13544 46461 13553 46495
rect 13553 46461 13587 46495
rect 13587 46461 13596 46495
rect 13544 46452 13596 46461
rect 15936 46452 15988 46504
rect 18144 46452 18196 46504
rect 18696 46495 18748 46504
rect 18696 46461 18705 46495
rect 18705 46461 18739 46495
rect 18739 46461 18748 46495
rect 18696 46452 18748 46461
rect 23112 46452 23164 46504
rect 23204 46452 23256 46504
rect 26608 46452 26660 46504
rect 10416 46384 10468 46436
rect 17224 46384 17276 46436
rect 27436 46520 27488 46572
rect 28540 46384 28592 46436
rect 1676 46359 1728 46368
rect 1676 46325 1685 46359
rect 1685 46325 1719 46359
rect 1719 46325 1728 46359
rect 1676 46316 1728 46325
rect 11704 46359 11756 46368
rect 11704 46325 11713 46359
rect 11713 46325 11747 46359
rect 11747 46325 11756 46359
rect 11704 46316 11756 46325
rect 16120 46316 16172 46368
rect 20260 46316 20312 46368
rect 26516 46316 26568 46368
rect 27252 46316 27304 46368
rect 4423 46214 4475 46266
rect 4487 46214 4539 46266
rect 4551 46214 4603 46266
rect 4615 46214 4667 46266
rect 4679 46214 4731 46266
rect 11369 46214 11421 46266
rect 11433 46214 11485 46266
rect 11497 46214 11549 46266
rect 11561 46214 11613 46266
rect 11625 46214 11677 46266
rect 18315 46214 18367 46266
rect 18379 46214 18431 46266
rect 18443 46214 18495 46266
rect 18507 46214 18559 46266
rect 18571 46214 18623 46266
rect 25261 46214 25313 46266
rect 25325 46214 25377 46266
rect 25389 46214 25441 46266
rect 25453 46214 25505 46266
rect 25517 46214 25569 46266
rect 7932 46155 7984 46164
rect 7932 46121 7941 46155
rect 7941 46121 7975 46155
rect 7975 46121 7984 46155
rect 7932 46112 7984 46121
rect 9496 46155 9548 46164
rect 9496 46121 9505 46155
rect 9505 46121 9539 46155
rect 9539 46121 9548 46155
rect 9496 46112 9548 46121
rect 10140 46155 10192 46164
rect 10140 46121 10149 46155
rect 10149 46121 10183 46155
rect 10183 46121 10192 46155
rect 10140 46112 10192 46121
rect 1032 45976 1084 46028
rect 2596 45976 2648 46028
rect 17224 46112 17276 46164
rect 18144 46112 18196 46164
rect 23112 46155 23164 46164
rect 23112 46121 23121 46155
rect 23121 46121 23155 46155
rect 23155 46121 23164 46155
rect 23112 46112 23164 46121
rect 3424 45951 3476 45960
rect 3424 45917 3433 45951
rect 3433 45917 3467 45951
rect 3467 45917 3476 45951
rect 3976 45951 4028 45960
rect 3424 45908 3476 45917
rect 3976 45917 3985 45951
rect 3985 45917 4019 45951
rect 4019 45917 4028 45951
rect 3976 45908 4028 45917
rect 7748 45908 7800 45960
rect 11704 45976 11756 46028
rect 11796 46019 11848 46028
rect 11796 45985 11805 46019
rect 11805 45985 11839 46019
rect 11839 45985 11848 46019
rect 15936 46019 15988 46028
rect 11796 45976 11848 45985
rect 15936 45985 15945 46019
rect 15945 45985 15979 46019
rect 15979 45985 15988 46019
rect 15936 45976 15988 45985
rect 16120 46019 16172 46028
rect 16120 45985 16129 46019
rect 16129 45985 16163 46019
rect 16163 45985 16172 46019
rect 16120 45976 16172 45985
rect 16764 46019 16816 46028
rect 16764 45985 16773 46019
rect 16773 45985 16807 46019
rect 16807 45985 16816 46019
rect 16764 45976 16816 45985
rect 20260 46019 20312 46028
rect 20260 45985 20269 46019
rect 20269 45985 20303 46019
rect 20303 45985 20312 46019
rect 20260 45976 20312 45985
rect 21272 46019 21324 46028
rect 21272 45985 21281 46019
rect 21281 45985 21315 46019
rect 21315 45985 21324 46019
rect 21272 45976 21324 45985
rect 9220 45908 9272 45960
rect 10692 45951 10744 45960
rect 3240 45883 3292 45892
rect 3240 45849 3249 45883
rect 3249 45849 3283 45883
rect 3283 45849 3292 45883
rect 3240 45840 3292 45849
rect 4160 45883 4212 45892
rect 4160 45849 4169 45883
rect 4169 45849 4203 45883
rect 4203 45849 4212 45883
rect 4160 45840 4212 45849
rect 10692 45917 10701 45951
rect 10701 45917 10735 45951
rect 10735 45917 10744 45951
rect 10692 45908 10744 45917
rect 14188 45908 14240 45960
rect 18328 45951 18380 45960
rect 18328 45917 18337 45951
rect 18337 45917 18371 45951
rect 18371 45917 18380 45951
rect 18328 45908 18380 45917
rect 23204 45951 23256 45960
rect 23204 45917 23213 45951
rect 23213 45917 23247 45951
rect 23247 45917 23256 45951
rect 23204 45908 23256 45917
rect 24952 45908 25004 45960
rect 27436 46044 27488 46096
rect 26516 46019 26568 46028
rect 26516 45985 26525 46019
rect 26525 45985 26559 46019
rect 26559 45985 26568 46019
rect 26516 45976 26568 45985
rect 27712 46019 27764 46028
rect 27712 45985 27721 46019
rect 27721 45985 27755 46019
rect 27755 45985 27764 46019
rect 27712 45976 27764 45985
rect 20444 45883 20496 45892
rect 20444 45849 20453 45883
rect 20453 45849 20487 45883
rect 20487 45849 20496 45883
rect 20444 45840 20496 45849
rect 21272 45840 21324 45892
rect 22560 45840 22612 45892
rect 12716 45772 12768 45824
rect 13268 45772 13320 45824
rect 15844 45772 15896 45824
rect 20352 45772 20404 45824
rect 7896 45670 7948 45722
rect 7960 45670 8012 45722
rect 8024 45670 8076 45722
rect 8088 45670 8140 45722
rect 8152 45670 8204 45722
rect 14842 45670 14894 45722
rect 14906 45670 14958 45722
rect 14970 45670 15022 45722
rect 15034 45670 15086 45722
rect 15098 45670 15150 45722
rect 21788 45670 21840 45722
rect 21852 45670 21904 45722
rect 21916 45670 21968 45722
rect 21980 45670 22032 45722
rect 22044 45670 22096 45722
rect 28734 45670 28786 45722
rect 28798 45670 28850 45722
rect 28862 45670 28914 45722
rect 28926 45670 28978 45722
rect 28990 45670 29042 45722
rect 13084 45568 13136 45620
rect 18328 45568 18380 45620
rect 20444 45611 20496 45620
rect 4160 45500 4212 45552
rect 20444 45577 20453 45611
rect 20453 45577 20487 45611
rect 20487 45577 20496 45611
rect 20444 45568 20496 45577
rect 27712 45568 27764 45620
rect 1676 45475 1728 45484
rect 1676 45441 1685 45475
rect 1685 45441 1719 45475
rect 1719 45441 1728 45475
rect 1676 45432 1728 45441
rect 2044 45364 2096 45416
rect 20 45296 72 45348
rect 2504 45364 2556 45416
rect 9312 45432 9364 45484
rect 10416 45475 10468 45484
rect 10416 45441 10425 45475
rect 10425 45441 10459 45475
rect 10459 45441 10468 45475
rect 10416 45432 10468 45441
rect 13268 45475 13320 45484
rect 13268 45441 13277 45475
rect 13277 45441 13311 45475
rect 13311 45441 13320 45475
rect 27252 45500 27304 45552
rect 14188 45475 14240 45484
rect 13268 45432 13320 45441
rect 14188 45441 14197 45475
rect 14197 45441 14231 45475
rect 14231 45441 14240 45475
rect 14188 45432 14240 45441
rect 20352 45475 20404 45484
rect 20352 45441 20361 45475
rect 20361 45441 20395 45475
rect 20395 45441 20404 45475
rect 20352 45432 20404 45441
rect 27896 45432 27948 45484
rect 14372 45407 14424 45416
rect 14372 45373 14381 45407
rect 14381 45373 14415 45407
rect 14415 45373 14424 45407
rect 14372 45364 14424 45373
rect 15200 45407 15252 45416
rect 15200 45373 15209 45407
rect 15209 45373 15243 45407
rect 15243 45373 15252 45407
rect 15200 45364 15252 45373
rect 26056 45407 26108 45416
rect 26056 45373 26065 45407
rect 26065 45373 26099 45407
rect 26099 45373 26108 45407
rect 26056 45364 26108 45373
rect 27988 45296 28040 45348
rect 20352 45228 20404 45280
rect 21640 45228 21692 45280
rect 27344 45228 27396 45280
rect 28356 45228 28408 45280
rect 4423 45126 4475 45178
rect 4487 45126 4539 45178
rect 4551 45126 4603 45178
rect 4615 45126 4667 45178
rect 4679 45126 4731 45178
rect 11369 45126 11421 45178
rect 11433 45126 11485 45178
rect 11497 45126 11549 45178
rect 11561 45126 11613 45178
rect 11625 45126 11677 45178
rect 18315 45126 18367 45178
rect 18379 45126 18431 45178
rect 18443 45126 18495 45178
rect 18507 45126 18559 45178
rect 18571 45126 18623 45178
rect 25261 45126 25313 45178
rect 25325 45126 25377 45178
rect 25389 45126 25441 45178
rect 25453 45126 25505 45178
rect 25517 45126 25569 45178
rect 2044 45067 2096 45076
rect 2044 45033 2053 45067
rect 2053 45033 2087 45067
rect 2087 45033 2096 45067
rect 2044 45024 2096 45033
rect 3976 45024 4028 45076
rect 27528 44931 27580 44940
rect 27528 44897 27537 44931
rect 27537 44897 27571 44931
rect 27571 44897 27580 44931
rect 27528 44888 27580 44897
rect 28356 44931 28408 44940
rect 28356 44897 28365 44931
rect 28365 44897 28399 44931
rect 28399 44897 28408 44931
rect 28356 44888 28408 44897
rect 2504 44820 2556 44872
rect 5172 44820 5224 44872
rect 23204 44820 23256 44872
rect 26240 44820 26292 44872
rect 27896 44752 27948 44804
rect 7896 44582 7948 44634
rect 7960 44582 8012 44634
rect 8024 44582 8076 44634
rect 8088 44582 8140 44634
rect 8152 44582 8204 44634
rect 14842 44582 14894 44634
rect 14906 44582 14958 44634
rect 14970 44582 15022 44634
rect 15034 44582 15086 44634
rect 15098 44582 15150 44634
rect 21788 44582 21840 44634
rect 21852 44582 21904 44634
rect 21916 44582 21968 44634
rect 21980 44582 22032 44634
rect 22044 44582 22096 44634
rect 28734 44582 28786 44634
rect 28798 44582 28850 44634
rect 28862 44582 28914 44634
rect 28926 44582 28978 44634
rect 28990 44582 29042 44634
rect 3240 44480 3292 44532
rect 14372 44480 14424 44532
rect 27896 44523 27948 44532
rect 27896 44489 27905 44523
rect 27905 44489 27939 44523
rect 27939 44489 27948 44523
rect 27896 44480 27948 44489
rect 25044 44412 25096 44464
rect 4344 44344 4396 44396
rect 5172 44344 5224 44396
rect 14372 44344 14424 44396
rect 19340 44344 19392 44396
rect 27160 44387 27212 44396
rect 27160 44353 27169 44387
rect 27169 44353 27203 44387
rect 27203 44353 27212 44387
rect 27160 44344 27212 44353
rect 27988 44344 28040 44396
rect 24952 44276 25004 44328
rect 26148 44319 26200 44328
rect 26148 44285 26157 44319
rect 26157 44285 26191 44319
rect 26191 44285 26200 44319
rect 26148 44276 26200 44285
rect 2964 44183 3016 44192
rect 2964 44149 2973 44183
rect 2973 44149 3007 44183
rect 3007 44149 3016 44183
rect 2964 44140 3016 44149
rect 26424 44140 26476 44192
rect 4423 44038 4475 44090
rect 4487 44038 4539 44090
rect 4551 44038 4603 44090
rect 4615 44038 4667 44090
rect 4679 44038 4731 44090
rect 11369 44038 11421 44090
rect 11433 44038 11485 44090
rect 11497 44038 11549 44090
rect 11561 44038 11613 44090
rect 11625 44038 11677 44090
rect 18315 44038 18367 44090
rect 18379 44038 18431 44090
rect 18443 44038 18495 44090
rect 18507 44038 18559 44090
rect 18571 44038 18623 44090
rect 25261 44038 25313 44090
rect 25325 44038 25377 44090
rect 25389 44038 25441 44090
rect 25453 44038 25505 44090
rect 25517 44038 25569 44090
rect 3424 43936 3476 43988
rect 21272 43843 21324 43852
rect 21272 43809 21281 43843
rect 21281 43809 21315 43843
rect 21315 43809 21324 43843
rect 21272 43800 21324 43809
rect 26240 43843 26292 43852
rect 26240 43809 26249 43843
rect 26249 43809 26283 43843
rect 26283 43809 26292 43843
rect 26240 43800 26292 43809
rect 26424 43843 26476 43852
rect 26424 43809 26433 43843
rect 26433 43809 26467 43843
rect 26467 43809 26476 43843
rect 28080 43843 28132 43852
rect 26424 43800 26476 43809
rect 28080 43809 28089 43843
rect 28089 43809 28123 43843
rect 28123 43809 28132 43843
rect 28080 43800 28132 43809
rect 1584 43732 1636 43784
rect 5080 43732 5132 43784
rect 10692 43732 10744 43784
rect 19432 43775 19484 43784
rect 19432 43741 19441 43775
rect 19441 43741 19475 43775
rect 19475 43741 19484 43775
rect 19432 43732 19484 43741
rect 19616 43707 19668 43716
rect 19616 43673 19625 43707
rect 19625 43673 19659 43707
rect 19659 43673 19668 43707
rect 19616 43664 19668 43673
rect 3148 43596 3200 43648
rect 7896 43494 7948 43546
rect 7960 43494 8012 43546
rect 8024 43494 8076 43546
rect 8088 43494 8140 43546
rect 8152 43494 8204 43546
rect 14842 43494 14894 43546
rect 14906 43494 14958 43546
rect 14970 43494 15022 43546
rect 15034 43494 15086 43546
rect 15098 43494 15150 43546
rect 21788 43494 21840 43546
rect 21852 43494 21904 43546
rect 21916 43494 21968 43546
rect 21980 43494 22032 43546
rect 22044 43494 22096 43546
rect 28734 43494 28786 43546
rect 28798 43494 28850 43546
rect 28862 43494 28914 43546
rect 28926 43494 28978 43546
rect 28990 43494 29042 43546
rect 3056 43392 3108 43444
rect 15844 43392 15896 43444
rect 19616 43392 19668 43444
rect 3148 43367 3200 43376
rect 3148 43333 3157 43367
rect 3157 43333 3191 43367
rect 3191 43333 3200 43367
rect 3148 43324 3200 43333
rect 2964 43299 3016 43308
rect 2964 43265 2973 43299
rect 2973 43265 3007 43299
rect 3007 43265 3016 43299
rect 2964 43256 3016 43265
rect 19340 43256 19392 43308
rect 27160 43256 27212 43308
rect 4160 43231 4212 43240
rect 4160 43197 4169 43231
rect 4169 43197 4203 43231
rect 4203 43197 4212 43231
rect 4160 43188 4212 43197
rect 3056 43120 3108 43172
rect 1768 43052 1820 43104
rect 26700 43052 26752 43104
rect 27160 43095 27212 43104
rect 27160 43061 27169 43095
rect 27169 43061 27203 43095
rect 27203 43061 27212 43095
rect 27160 43052 27212 43061
rect 28080 43095 28132 43104
rect 28080 43061 28089 43095
rect 28089 43061 28123 43095
rect 28123 43061 28132 43095
rect 28080 43052 28132 43061
rect 4423 42950 4475 43002
rect 4487 42950 4539 43002
rect 4551 42950 4603 43002
rect 4615 42950 4667 43002
rect 4679 42950 4731 43002
rect 11369 42950 11421 43002
rect 11433 42950 11485 43002
rect 11497 42950 11549 43002
rect 11561 42950 11613 43002
rect 11625 42950 11677 43002
rect 18315 42950 18367 43002
rect 18379 42950 18431 43002
rect 18443 42950 18495 43002
rect 18507 42950 18559 43002
rect 18571 42950 18623 43002
rect 25261 42950 25313 43002
rect 25325 42950 25377 43002
rect 25389 42950 25441 43002
rect 25453 42950 25505 43002
rect 25517 42950 25569 43002
rect 1584 42755 1636 42764
rect 1584 42721 1593 42755
rect 1593 42721 1627 42755
rect 1627 42721 1636 42755
rect 1584 42712 1636 42721
rect 1768 42755 1820 42764
rect 1768 42721 1777 42755
rect 1777 42721 1811 42755
rect 1811 42721 1820 42755
rect 1768 42712 1820 42721
rect 2780 42755 2832 42764
rect 2780 42721 2789 42755
rect 2789 42721 2823 42755
rect 2823 42721 2832 42755
rect 2780 42712 2832 42721
rect 27160 42712 27212 42764
rect 28356 42755 28408 42764
rect 28356 42721 28365 42755
rect 28365 42721 28399 42755
rect 28399 42721 28408 42755
rect 28356 42712 28408 42721
rect 26700 42619 26752 42628
rect 26700 42585 26709 42619
rect 26709 42585 26743 42619
rect 26743 42585 26752 42619
rect 26700 42576 26752 42585
rect 7896 42406 7948 42458
rect 7960 42406 8012 42458
rect 8024 42406 8076 42458
rect 8088 42406 8140 42458
rect 8152 42406 8204 42458
rect 14842 42406 14894 42458
rect 14906 42406 14958 42458
rect 14970 42406 15022 42458
rect 15034 42406 15086 42458
rect 15098 42406 15150 42458
rect 21788 42406 21840 42458
rect 21852 42406 21904 42458
rect 21916 42406 21968 42458
rect 21980 42406 22032 42458
rect 22044 42406 22096 42458
rect 28734 42406 28786 42458
rect 28798 42406 28850 42458
rect 28862 42406 28914 42458
rect 28926 42406 28978 42458
rect 28990 42406 29042 42458
rect 2872 42168 2924 42220
rect 27712 42211 27764 42220
rect 27712 42177 27721 42211
rect 27721 42177 27755 42211
rect 27755 42177 27764 42211
rect 27712 42168 27764 42177
rect 1676 42007 1728 42016
rect 1676 41973 1685 42007
rect 1685 41973 1719 42007
rect 1719 41973 1728 42007
rect 1676 41964 1728 41973
rect 3240 41964 3292 42016
rect 3424 41964 3476 42016
rect 28172 41964 28224 42016
rect 4423 41862 4475 41914
rect 4487 41862 4539 41914
rect 4551 41862 4603 41914
rect 4615 41862 4667 41914
rect 4679 41862 4731 41914
rect 11369 41862 11421 41914
rect 11433 41862 11485 41914
rect 11497 41862 11549 41914
rect 11561 41862 11613 41914
rect 11625 41862 11677 41914
rect 18315 41862 18367 41914
rect 18379 41862 18431 41914
rect 18443 41862 18495 41914
rect 18507 41862 18559 41914
rect 18571 41862 18623 41914
rect 25261 41862 25313 41914
rect 25325 41862 25377 41914
rect 25389 41862 25441 41914
rect 25453 41862 25505 41914
rect 25517 41862 25569 41914
rect 28080 41692 28132 41744
rect 3240 41667 3292 41676
rect 3240 41633 3249 41667
rect 3249 41633 3283 41667
rect 3283 41633 3292 41667
rect 3240 41624 3292 41633
rect 3424 41667 3476 41676
rect 3424 41633 3433 41667
rect 3433 41633 3467 41667
rect 3467 41633 3476 41667
rect 3424 41624 3476 41633
rect 27528 41667 27580 41676
rect 27528 41633 27537 41667
rect 27537 41633 27571 41667
rect 27571 41633 27580 41667
rect 27528 41624 27580 41633
rect 28172 41667 28224 41676
rect 28172 41633 28181 41667
rect 28181 41633 28215 41667
rect 28215 41633 28224 41667
rect 28172 41624 28224 41633
rect 1584 41599 1636 41608
rect 1584 41565 1593 41599
rect 1593 41565 1627 41599
rect 1627 41565 1636 41599
rect 1584 41556 1636 41565
rect 7896 41318 7948 41370
rect 7960 41318 8012 41370
rect 8024 41318 8076 41370
rect 8088 41318 8140 41370
rect 8152 41318 8204 41370
rect 14842 41318 14894 41370
rect 14906 41318 14958 41370
rect 14970 41318 15022 41370
rect 15034 41318 15086 41370
rect 15098 41318 15150 41370
rect 21788 41318 21840 41370
rect 21852 41318 21904 41370
rect 21916 41318 21968 41370
rect 21980 41318 22032 41370
rect 22044 41318 22096 41370
rect 28734 41318 28786 41370
rect 28798 41318 28850 41370
rect 28862 41318 28914 41370
rect 28926 41318 28978 41370
rect 28990 41318 29042 41370
rect 1676 41123 1728 41132
rect 1676 41089 1685 41123
rect 1685 41089 1719 41123
rect 1719 41089 1728 41123
rect 1676 41080 1728 41089
rect 27436 41123 27488 41132
rect 27436 41089 27445 41123
rect 27445 41089 27479 41123
rect 27479 41089 27488 41123
rect 27436 41080 27488 41089
rect 2320 41012 2372 41064
rect 2780 41055 2832 41064
rect 2780 41021 2789 41055
rect 2789 41021 2823 41055
rect 2823 41021 2832 41055
rect 2780 41012 2832 41021
rect 28172 40876 28224 40928
rect 28356 40876 28408 40928
rect 4423 40774 4475 40826
rect 4487 40774 4539 40826
rect 4551 40774 4603 40826
rect 4615 40774 4667 40826
rect 4679 40774 4731 40826
rect 11369 40774 11421 40826
rect 11433 40774 11485 40826
rect 11497 40774 11549 40826
rect 11561 40774 11613 40826
rect 11625 40774 11677 40826
rect 18315 40774 18367 40826
rect 18379 40774 18431 40826
rect 18443 40774 18495 40826
rect 18507 40774 18559 40826
rect 18571 40774 18623 40826
rect 25261 40774 25313 40826
rect 25325 40774 25377 40826
rect 25389 40774 25441 40826
rect 25453 40774 25505 40826
rect 25517 40774 25569 40826
rect 27528 40579 27580 40588
rect 27528 40545 27537 40579
rect 27537 40545 27571 40579
rect 27571 40545 27580 40579
rect 27528 40536 27580 40545
rect 28172 40579 28224 40588
rect 28172 40545 28181 40579
rect 28181 40545 28215 40579
rect 28215 40545 28224 40579
rect 28172 40536 28224 40545
rect 28356 40579 28408 40588
rect 28356 40545 28365 40579
rect 28365 40545 28399 40579
rect 28399 40545 28408 40579
rect 28356 40536 28408 40545
rect 1952 40511 2004 40520
rect 1952 40477 1961 40511
rect 1961 40477 1995 40511
rect 1995 40477 2004 40511
rect 1952 40468 2004 40477
rect 2412 40511 2464 40520
rect 2412 40477 2421 40511
rect 2421 40477 2455 40511
rect 2455 40477 2464 40511
rect 2412 40468 2464 40477
rect 17868 40468 17920 40520
rect 18604 40511 18656 40520
rect 18604 40477 18613 40511
rect 18613 40477 18647 40511
rect 18647 40477 18656 40511
rect 18604 40468 18656 40477
rect 18236 40400 18288 40452
rect 1860 40375 1912 40384
rect 1860 40341 1869 40375
rect 1869 40341 1903 40375
rect 1903 40341 1912 40375
rect 1860 40332 1912 40341
rect 17500 40332 17552 40384
rect 18696 40375 18748 40384
rect 18696 40341 18705 40375
rect 18705 40341 18739 40375
rect 18739 40341 18748 40375
rect 18696 40332 18748 40341
rect 7896 40230 7948 40282
rect 7960 40230 8012 40282
rect 8024 40230 8076 40282
rect 8088 40230 8140 40282
rect 8152 40230 8204 40282
rect 14842 40230 14894 40282
rect 14906 40230 14958 40282
rect 14970 40230 15022 40282
rect 15034 40230 15086 40282
rect 15098 40230 15150 40282
rect 21788 40230 21840 40282
rect 21852 40230 21904 40282
rect 21916 40230 21968 40282
rect 21980 40230 22032 40282
rect 22044 40230 22096 40282
rect 28734 40230 28786 40282
rect 28798 40230 28850 40282
rect 28862 40230 28914 40282
rect 28926 40230 28978 40282
rect 28990 40230 29042 40282
rect 18604 40128 18656 40180
rect 19248 40128 19300 40180
rect 1860 40103 1912 40112
rect 1860 40069 1869 40103
rect 1869 40069 1903 40103
rect 1903 40069 1912 40103
rect 1860 40060 1912 40069
rect 3516 40103 3568 40112
rect 3516 40069 3525 40103
rect 3525 40069 3559 40103
rect 3559 40069 3568 40103
rect 3516 40060 3568 40069
rect 17868 40060 17920 40112
rect 17224 40035 17276 40044
rect 17224 40001 17233 40035
rect 17233 40001 17267 40035
rect 17267 40001 17276 40035
rect 17224 39992 17276 40001
rect 17500 40035 17552 40044
rect 17500 40001 17509 40035
rect 17509 40001 17543 40035
rect 17543 40001 17552 40035
rect 17500 39992 17552 40001
rect 18880 39992 18932 40044
rect 19616 40035 19668 40044
rect 19616 40001 19625 40035
rect 19625 40001 19659 40035
rect 19659 40001 19668 40035
rect 19616 39992 19668 40001
rect 2412 39924 2464 39976
rect 16304 39924 16356 39976
rect 17316 39899 17368 39908
rect 17316 39865 17325 39899
rect 17325 39865 17359 39899
rect 17359 39865 17368 39899
rect 17316 39856 17368 39865
rect 20904 39924 20956 39976
rect 17040 39831 17092 39840
rect 17040 39797 17049 39831
rect 17049 39797 17083 39831
rect 17083 39797 17092 39831
rect 17040 39788 17092 39797
rect 18236 39788 18288 39840
rect 19248 39788 19300 39840
rect 26516 39788 26568 39840
rect 27528 39788 27580 39840
rect 4423 39686 4475 39738
rect 4487 39686 4539 39738
rect 4551 39686 4603 39738
rect 4615 39686 4667 39738
rect 4679 39686 4731 39738
rect 11369 39686 11421 39738
rect 11433 39686 11485 39738
rect 11497 39686 11549 39738
rect 11561 39686 11613 39738
rect 11625 39686 11677 39738
rect 18315 39686 18367 39738
rect 18379 39686 18431 39738
rect 18443 39686 18495 39738
rect 18507 39686 18559 39738
rect 18571 39686 18623 39738
rect 25261 39686 25313 39738
rect 25325 39686 25377 39738
rect 25389 39686 25441 39738
rect 25453 39686 25505 39738
rect 25517 39686 25569 39738
rect 2320 39627 2372 39636
rect 2320 39593 2329 39627
rect 2329 39593 2363 39627
rect 2363 39593 2372 39627
rect 2320 39584 2372 39593
rect 17316 39584 17368 39636
rect 1952 39448 2004 39500
rect 18236 39516 18288 39568
rect 18696 39516 18748 39568
rect 18880 39516 18932 39568
rect 19248 39448 19300 39500
rect 18604 39423 18656 39432
rect 2872 39312 2924 39364
rect 17868 39312 17920 39364
rect 18604 39389 18613 39423
rect 18613 39389 18647 39423
rect 18647 39389 18656 39423
rect 18604 39380 18656 39389
rect 18696 39423 18748 39432
rect 18696 39389 18705 39423
rect 18705 39389 18739 39423
rect 18739 39389 18748 39423
rect 18696 39380 18748 39389
rect 18880 39423 18932 39432
rect 18880 39389 18889 39423
rect 18889 39389 18923 39423
rect 18923 39389 18932 39423
rect 18880 39380 18932 39389
rect 19800 39423 19852 39432
rect 19800 39389 19809 39423
rect 19809 39389 19843 39423
rect 19843 39389 19852 39423
rect 26516 39491 26568 39500
rect 26516 39457 26525 39491
rect 26525 39457 26559 39491
rect 26559 39457 26568 39491
rect 26516 39448 26568 39457
rect 28632 39448 28684 39500
rect 19800 39380 19852 39389
rect 20260 39380 20312 39432
rect 20904 39380 20956 39432
rect 3148 39244 3200 39296
rect 17224 39244 17276 39296
rect 18144 39244 18196 39296
rect 19248 39244 19300 39296
rect 27896 39312 27948 39364
rect 19984 39244 20036 39296
rect 20628 39244 20680 39296
rect 7896 39142 7948 39194
rect 7960 39142 8012 39194
rect 8024 39142 8076 39194
rect 8088 39142 8140 39194
rect 8152 39142 8204 39194
rect 14842 39142 14894 39194
rect 14906 39142 14958 39194
rect 14970 39142 15022 39194
rect 15034 39142 15086 39194
rect 15098 39142 15150 39194
rect 21788 39142 21840 39194
rect 21852 39142 21904 39194
rect 21916 39142 21968 39194
rect 21980 39142 22032 39194
rect 22044 39142 22096 39194
rect 28734 39142 28786 39194
rect 28798 39142 28850 39194
rect 28862 39142 28914 39194
rect 28926 39142 28978 39194
rect 28990 39142 29042 39194
rect 18604 39040 18656 39092
rect 18052 38972 18104 39024
rect 18696 38972 18748 39024
rect 18236 38947 18288 38956
rect 18236 38913 18245 38947
rect 18245 38913 18279 38947
rect 18279 38913 18288 38947
rect 19800 39040 19852 39092
rect 18236 38904 18288 38913
rect 19616 38904 19668 38956
rect 20444 38836 20496 38888
rect 3424 38768 3476 38820
rect 3976 38700 4028 38752
rect 18788 38700 18840 38752
rect 20904 38904 20956 38956
rect 27528 38904 27580 38956
rect 27712 38947 27764 38956
rect 27712 38913 27721 38947
rect 27721 38913 27755 38947
rect 27755 38913 27764 38947
rect 27712 38904 27764 38913
rect 28632 38904 28684 38956
rect 22192 38879 22244 38888
rect 22192 38845 22201 38879
rect 22201 38845 22235 38879
rect 22235 38845 22244 38879
rect 22192 38836 22244 38845
rect 23480 38879 23532 38888
rect 23480 38845 23489 38879
rect 23489 38845 23523 38879
rect 23523 38845 23532 38879
rect 23480 38836 23532 38845
rect 26148 38879 26200 38888
rect 26148 38845 26157 38879
rect 26157 38845 26191 38879
rect 26191 38845 26200 38879
rect 26148 38836 26200 38845
rect 23112 38768 23164 38820
rect 4423 38598 4475 38650
rect 4487 38598 4539 38650
rect 4551 38598 4603 38650
rect 4615 38598 4667 38650
rect 4679 38598 4731 38650
rect 11369 38598 11421 38650
rect 11433 38598 11485 38650
rect 11497 38598 11549 38650
rect 11561 38598 11613 38650
rect 11625 38598 11677 38650
rect 18315 38598 18367 38650
rect 18379 38598 18431 38650
rect 18443 38598 18495 38650
rect 18507 38598 18559 38650
rect 18571 38598 18623 38650
rect 25261 38598 25313 38650
rect 25325 38598 25377 38650
rect 25389 38598 25441 38650
rect 25453 38598 25505 38650
rect 25517 38598 25569 38650
rect 15292 38496 15344 38548
rect 16120 38428 16172 38480
rect 15476 38403 15528 38412
rect 15476 38369 15485 38403
rect 15485 38369 15519 38403
rect 15519 38369 15528 38403
rect 15476 38360 15528 38369
rect 15844 38360 15896 38412
rect 1676 38335 1728 38344
rect 1676 38301 1685 38335
rect 1685 38301 1719 38335
rect 1719 38301 1728 38335
rect 1676 38292 1728 38301
rect 5540 38292 5592 38344
rect 16120 38335 16172 38344
rect 16120 38301 16129 38335
rect 16129 38301 16163 38335
rect 16163 38301 16172 38335
rect 16120 38292 16172 38301
rect 22192 38496 22244 38548
rect 15292 38267 15344 38276
rect 15292 38233 15301 38267
rect 15301 38233 15335 38267
rect 15335 38233 15344 38267
rect 15292 38224 15344 38233
rect 17316 38292 17368 38344
rect 3240 38156 3292 38208
rect 16028 38156 16080 38208
rect 17132 38156 17184 38208
rect 17592 38292 17644 38344
rect 17960 38292 18012 38344
rect 21640 38292 21692 38344
rect 27712 38360 27764 38412
rect 28264 38403 28316 38412
rect 28264 38369 28273 38403
rect 28273 38369 28307 38403
rect 28307 38369 28316 38403
rect 28264 38360 28316 38369
rect 26516 38335 26568 38344
rect 26516 38301 26525 38335
rect 26525 38301 26559 38335
rect 26559 38301 26568 38335
rect 26516 38292 26568 38301
rect 18052 38224 18104 38276
rect 26700 38267 26752 38276
rect 26700 38233 26709 38267
rect 26709 38233 26743 38267
rect 26743 38233 26752 38267
rect 26700 38224 26752 38233
rect 17960 38156 18012 38208
rect 18420 38156 18472 38208
rect 7896 38054 7948 38106
rect 7960 38054 8012 38106
rect 8024 38054 8076 38106
rect 8088 38054 8140 38106
rect 8152 38054 8204 38106
rect 14842 38054 14894 38106
rect 14906 38054 14958 38106
rect 14970 38054 15022 38106
rect 15034 38054 15086 38106
rect 15098 38054 15150 38106
rect 21788 38054 21840 38106
rect 21852 38054 21904 38106
rect 21916 38054 21968 38106
rect 21980 38054 22032 38106
rect 22044 38054 22096 38106
rect 28734 38054 28786 38106
rect 28798 38054 28850 38106
rect 28862 38054 28914 38106
rect 28926 38054 28978 38106
rect 28990 38054 29042 38106
rect 15476 37952 15528 38004
rect 27896 37995 27948 38004
rect 27896 37961 27905 37995
rect 27905 37961 27939 37995
rect 27939 37961 27948 37995
rect 27896 37952 27948 37961
rect 3976 37859 4028 37868
rect 3976 37825 3985 37859
rect 3985 37825 4019 37859
rect 4019 37825 4028 37859
rect 3976 37816 4028 37825
rect 4896 37816 4948 37868
rect 16028 37859 16080 37868
rect 16028 37825 16037 37859
rect 16037 37825 16071 37859
rect 16071 37825 16080 37859
rect 16028 37816 16080 37825
rect 16396 37816 16448 37868
rect 2780 37791 2832 37800
rect 2780 37757 2789 37791
rect 2789 37757 2823 37791
rect 2823 37757 2832 37791
rect 2780 37748 2832 37757
rect 16580 37748 16632 37800
rect 17316 37859 17368 37868
rect 17316 37825 17325 37859
rect 17325 37825 17359 37859
rect 17359 37825 17368 37859
rect 18236 37859 18288 37868
rect 17316 37816 17368 37825
rect 18236 37825 18245 37859
rect 18245 37825 18279 37859
rect 18279 37825 18288 37859
rect 18236 37816 18288 37825
rect 18420 37859 18472 37868
rect 18420 37825 18429 37859
rect 18429 37825 18463 37859
rect 18463 37825 18472 37859
rect 18420 37816 18472 37825
rect 18696 37816 18748 37868
rect 19524 37859 19576 37868
rect 17132 37680 17184 37732
rect 18512 37791 18564 37800
rect 18512 37757 18521 37791
rect 18521 37757 18555 37791
rect 18555 37757 18564 37791
rect 18512 37748 18564 37757
rect 19524 37825 19533 37859
rect 19533 37825 19567 37859
rect 19567 37825 19576 37859
rect 19524 37816 19576 37825
rect 26516 37816 26568 37868
rect 27804 37859 27856 37868
rect 27804 37825 27813 37859
rect 27813 37825 27847 37859
rect 27847 37825 27856 37859
rect 27804 37816 27856 37825
rect 20076 37748 20128 37800
rect 16948 37612 17000 37664
rect 17592 37612 17644 37664
rect 18236 37612 18288 37664
rect 19156 37612 19208 37664
rect 19616 37655 19668 37664
rect 19616 37621 19625 37655
rect 19625 37621 19659 37655
rect 19659 37621 19668 37655
rect 19616 37612 19668 37621
rect 4423 37510 4475 37562
rect 4487 37510 4539 37562
rect 4551 37510 4603 37562
rect 4615 37510 4667 37562
rect 4679 37510 4731 37562
rect 11369 37510 11421 37562
rect 11433 37510 11485 37562
rect 11497 37510 11549 37562
rect 11561 37510 11613 37562
rect 11625 37510 11677 37562
rect 18315 37510 18367 37562
rect 18379 37510 18431 37562
rect 18443 37510 18495 37562
rect 18507 37510 18559 37562
rect 18571 37510 18623 37562
rect 25261 37510 25313 37562
rect 25325 37510 25377 37562
rect 25389 37510 25441 37562
rect 25453 37510 25505 37562
rect 25517 37510 25569 37562
rect 17132 37451 17184 37460
rect 17132 37417 17141 37451
rect 17141 37417 17175 37451
rect 17175 37417 17184 37451
rect 17132 37408 17184 37417
rect 17316 37451 17368 37460
rect 17316 37417 17325 37451
rect 17325 37417 17359 37451
rect 17359 37417 17368 37451
rect 17316 37408 17368 37417
rect 16212 37340 16264 37392
rect 18696 37408 18748 37460
rect 20076 37451 20128 37460
rect 20076 37417 20085 37451
rect 20085 37417 20119 37451
rect 20119 37417 20128 37451
rect 20076 37408 20128 37417
rect 20444 37408 20496 37460
rect 20720 37408 20772 37460
rect 24768 37383 24820 37392
rect 3240 37315 3292 37324
rect 3240 37281 3249 37315
rect 3249 37281 3283 37315
rect 3283 37281 3292 37315
rect 3240 37272 3292 37281
rect 15476 37315 15528 37324
rect 15476 37281 15485 37315
rect 15485 37281 15519 37315
rect 15519 37281 15528 37315
rect 15476 37272 15528 37281
rect 1584 37247 1636 37256
rect 1584 37213 1593 37247
rect 1593 37213 1627 37247
rect 1627 37213 1636 37247
rect 1584 37204 1636 37213
rect 3424 37247 3476 37256
rect 3424 37213 3433 37247
rect 3433 37213 3467 37247
rect 3467 37213 3476 37247
rect 3424 37204 3476 37213
rect 20536 37315 20588 37324
rect 3148 37136 3200 37188
rect 4160 37179 4212 37188
rect 4160 37145 4169 37179
rect 4169 37145 4203 37179
rect 4203 37145 4212 37179
rect 4160 37136 4212 37145
rect 18144 37247 18196 37256
rect 18144 37213 18159 37247
rect 18159 37213 18193 37247
rect 18193 37213 18196 37247
rect 18328 37247 18380 37256
rect 18144 37204 18196 37213
rect 18328 37213 18331 37247
rect 18331 37213 18365 37247
rect 18365 37213 18380 37247
rect 18328 37204 18380 37213
rect 16120 37136 16172 37188
rect 16580 37136 16632 37188
rect 17592 37136 17644 37188
rect 20536 37281 20545 37315
rect 20545 37281 20579 37315
rect 20579 37281 20588 37315
rect 20536 37272 20588 37281
rect 22376 37272 22428 37324
rect 24768 37349 24777 37383
rect 24777 37349 24811 37383
rect 24811 37349 24820 37383
rect 24768 37340 24820 37349
rect 26056 37340 26108 37392
rect 26240 37272 26292 37324
rect 20168 37204 20220 37256
rect 20444 37204 20496 37256
rect 20628 37247 20680 37256
rect 20628 37213 20637 37247
rect 20637 37213 20671 37247
rect 20671 37213 20680 37247
rect 20628 37204 20680 37213
rect 20812 37204 20864 37256
rect 21456 37204 21508 37256
rect 23756 37204 23808 37256
rect 24492 37204 24544 37256
rect 24768 37204 24820 37256
rect 28356 37247 28408 37256
rect 28356 37213 28365 37247
rect 28365 37213 28399 37247
rect 28399 37213 28408 37247
rect 28356 37204 28408 37213
rect 26056 37179 26108 37188
rect 6736 37068 6788 37120
rect 16028 37111 16080 37120
rect 16028 37077 16037 37111
rect 16037 37077 16071 37111
rect 16071 37077 16080 37111
rect 16028 37068 16080 37077
rect 18236 37111 18288 37120
rect 18236 37077 18245 37111
rect 18245 37077 18279 37111
rect 18279 37077 18288 37111
rect 18236 37068 18288 37077
rect 19064 37068 19116 37120
rect 21456 37068 21508 37120
rect 22744 37068 22796 37120
rect 23296 37111 23348 37120
rect 23296 37077 23305 37111
rect 23305 37077 23339 37111
rect 23339 37077 23348 37111
rect 23296 37068 23348 37077
rect 26056 37145 26065 37179
rect 26065 37145 26099 37179
rect 26099 37145 26108 37179
rect 26056 37136 26108 37145
rect 26332 37068 26384 37120
rect 28172 37111 28224 37120
rect 28172 37077 28181 37111
rect 28181 37077 28215 37111
rect 28215 37077 28224 37111
rect 28172 37068 28224 37077
rect 7896 36966 7948 37018
rect 7960 36966 8012 37018
rect 8024 36966 8076 37018
rect 8088 36966 8140 37018
rect 8152 36966 8204 37018
rect 14842 36966 14894 37018
rect 14906 36966 14958 37018
rect 14970 36966 15022 37018
rect 15034 36966 15086 37018
rect 15098 36966 15150 37018
rect 21788 36966 21840 37018
rect 21852 36966 21904 37018
rect 21916 36966 21968 37018
rect 21980 36966 22032 37018
rect 22044 36966 22096 37018
rect 28734 36966 28786 37018
rect 28798 36966 28850 37018
rect 28862 36966 28914 37018
rect 28926 36966 28978 37018
rect 28990 36966 29042 37018
rect 4160 36864 4212 36916
rect 17960 36864 18012 36916
rect 19984 36864 20036 36916
rect 20628 36864 20680 36916
rect 20812 36907 20864 36916
rect 20812 36873 20821 36907
rect 20821 36873 20855 36907
rect 20855 36873 20864 36907
rect 20812 36864 20864 36873
rect 23480 36864 23532 36916
rect 23940 36864 23992 36916
rect 26056 36864 26108 36916
rect 26700 36864 26752 36916
rect 3148 36796 3200 36848
rect 4344 36796 4396 36848
rect 4988 36796 5040 36848
rect 20260 36796 20312 36848
rect 20444 36796 20496 36848
rect 21456 36796 21508 36848
rect 4252 36728 4304 36780
rect 2596 36660 2648 36712
rect 4344 36660 4396 36712
rect 6000 36728 6052 36780
rect 19064 36771 19116 36780
rect 19064 36737 19073 36771
rect 19073 36737 19107 36771
rect 19107 36737 19116 36771
rect 19064 36728 19116 36737
rect 19248 36771 19300 36780
rect 19248 36737 19257 36771
rect 19257 36737 19291 36771
rect 19291 36737 19300 36771
rect 19248 36728 19300 36737
rect 20628 36771 20680 36780
rect 20628 36737 20637 36771
rect 20637 36737 20671 36771
rect 20671 36737 20680 36771
rect 20628 36728 20680 36737
rect 21272 36771 21324 36780
rect 21272 36737 21281 36771
rect 21281 36737 21315 36771
rect 21315 36737 21324 36771
rect 21272 36728 21324 36737
rect 23480 36728 23532 36780
rect 25964 36728 26016 36780
rect 27804 36796 27856 36848
rect 26976 36728 27028 36780
rect 16212 36703 16264 36712
rect 16212 36669 16221 36703
rect 16221 36669 16255 36703
rect 16255 36669 16264 36703
rect 16212 36660 16264 36669
rect 20352 36703 20404 36712
rect 20352 36669 20377 36703
rect 20377 36669 20404 36703
rect 20352 36660 20404 36669
rect 20720 36660 20772 36712
rect 4160 36592 4212 36644
rect 20812 36592 20864 36644
rect 1768 36567 1820 36576
rect 1768 36533 1777 36567
rect 1777 36533 1811 36567
rect 1811 36533 1820 36567
rect 1768 36524 1820 36533
rect 15752 36524 15804 36576
rect 19524 36524 19576 36576
rect 27896 36567 27948 36576
rect 27896 36533 27905 36567
rect 27905 36533 27939 36567
rect 27939 36533 27948 36567
rect 27896 36524 27948 36533
rect 4423 36422 4475 36474
rect 4487 36422 4539 36474
rect 4551 36422 4603 36474
rect 4615 36422 4667 36474
rect 4679 36422 4731 36474
rect 11369 36422 11421 36474
rect 11433 36422 11485 36474
rect 11497 36422 11549 36474
rect 11561 36422 11613 36474
rect 11625 36422 11677 36474
rect 18315 36422 18367 36474
rect 18379 36422 18431 36474
rect 18443 36422 18495 36474
rect 18507 36422 18559 36474
rect 18571 36422 18623 36474
rect 25261 36422 25313 36474
rect 25325 36422 25377 36474
rect 25389 36422 25441 36474
rect 25453 36422 25505 36474
rect 25517 36422 25569 36474
rect 4988 36320 5040 36372
rect 1676 36252 1728 36304
rect 19616 36320 19668 36372
rect 20812 36363 20864 36372
rect 20812 36329 20821 36363
rect 20821 36329 20855 36363
rect 20855 36329 20864 36363
rect 20812 36320 20864 36329
rect 27804 36252 27856 36304
rect 1768 36227 1820 36236
rect 1768 36193 1777 36227
rect 1777 36193 1811 36227
rect 1811 36193 1820 36227
rect 1768 36184 1820 36193
rect 2780 36227 2832 36236
rect 2780 36193 2789 36227
rect 2789 36193 2823 36227
rect 2823 36193 2832 36227
rect 2780 36184 2832 36193
rect 4252 36159 4304 36168
rect 4252 36125 4261 36159
rect 4261 36125 4295 36159
rect 4295 36125 4304 36159
rect 4252 36116 4304 36125
rect 18144 36184 18196 36236
rect 19064 36184 19116 36236
rect 17040 36116 17092 36168
rect 20168 36184 20220 36236
rect 23940 36184 23992 36236
rect 27896 36184 27948 36236
rect 4896 36091 4948 36100
rect 4896 36057 4905 36091
rect 4905 36057 4939 36091
rect 4939 36057 4948 36091
rect 4896 36048 4948 36057
rect 12072 36048 12124 36100
rect 19800 36048 19852 36100
rect 20352 36159 20404 36168
rect 20352 36125 20361 36159
rect 20361 36125 20395 36159
rect 20395 36125 20404 36159
rect 20812 36159 20864 36168
rect 20352 36116 20404 36125
rect 20812 36125 20821 36159
rect 20821 36125 20855 36159
rect 20855 36125 20864 36159
rect 20812 36116 20864 36125
rect 21272 36116 21324 36168
rect 22744 36159 22796 36168
rect 22744 36125 22753 36159
rect 22753 36125 22787 36159
rect 22787 36125 22796 36159
rect 22744 36116 22796 36125
rect 28356 36159 28408 36168
rect 28356 36125 28365 36159
rect 28365 36125 28399 36159
rect 28399 36125 28408 36159
rect 28356 36116 28408 36125
rect 20444 36048 20496 36100
rect 23480 36048 23532 36100
rect 24124 36048 24176 36100
rect 26700 36091 26752 36100
rect 26700 36057 26709 36091
rect 26709 36057 26743 36091
rect 26743 36057 26752 36091
rect 26700 36048 26752 36057
rect 17316 35980 17368 36032
rect 23020 35980 23072 36032
rect 7896 35878 7948 35930
rect 7960 35878 8012 35930
rect 8024 35878 8076 35930
rect 8088 35878 8140 35930
rect 8152 35878 8204 35930
rect 14842 35878 14894 35930
rect 14906 35878 14958 35930
rect 14970 35878 15022 35930
rect 15034 35878 15086 35930
rect 15098 35878 15150 35930
rect 21788 35878 21840 35930
rect 21852 35878 21904 35930
rect 21916 35878 21968 35930
rect 21980 35878 22032 35930
rect 22044 35878 22096 35930
rect 28734 35878 28786 35930
rect 28798 35878 28850 35930
rect 28862 35878 28914 35930
rect 28926 35878 28978 35930
rect 28990 35878 29042 35930
rect 2320 35751 2372 35760
rect 2320 35717 2329 35751
rect 2329 35717 2363 35751
rect 2363 35717 2372 35751
rect 2320 35708 2372 35717
rect 2596 35640 2648 35692
rect 4252 35640 4304 35692
rect 12072 35776 12124 35828
rect 12716 35751 12768 35760
rect 12716 35717 12725 35751
rect 12725 35717 12759 35751
rect 12759 35717 12768 35751
rect 12716 35708 12768 35717
rect 15752 35683 15804 35692
rect 15752 35649 15761 35683
rect 15761 35649 15795 35683
rect 15795 35649 15804 35683
rect 15752 35640 15804 35649
rect 18788 35708 18840 35760
rect 26700 35776 26752 35828
rect 26884 35708 26936 35760
rect 18236 35640 18288 35692
rect 23020 35683 23072 35692
rect 23020 35649 23029 35683
rect 23029 35649 23063 35683
rect 23063 35649 23072 35683
rect 23020 35640 23072 35649
rect 27252 35640 27304 35692
rect 28448 35640 28500 35692
rect 4160 35572 4212 35624
rect 4804 35572 4856 35624
rect 5724 35615 5776 35624
rect 5724 35581 5733 35615
rect 5733 35581 5767 35615
rect 5767 35581 5776 35615
rect 5724 35572 5776 35581
rect 15568 35615 15620 35624
rect 15568 35581 15577 35615
rect 15577 35581 15611 35615
rect 15611 35581 15620 35615
rect 15568 35572 15620 35581
rect 25688 35615 25740 35624
rect 25688 35581 25697 35615
rect 25697 35581 25731 35615
rect 25731 35581 25740 35615
rect 25688 35572 25740 35581
rect 19156 35504 19208 35556
rect 17132 35436 17184 35488
rect 22836 35479 22888 35488
rect 22836 35445 22845 35479
rect 22845 35445 22879 35479
rect 22879 35445 22888 35479
rect 22836 35436 22888 35445
rect 24952 35436 25004 35488
rect 26240 35479 26292 35488
rect 26240 35445 26249 35479
rect 26249 35445 26283 35479
rect 26283 35445 26292 35479
rect 27988 35479 28040 35488
rect 26240 35436 26292 35445
rect 27988 35445 27997 35479
rect 27997 35445 28031 35479
rect 28031 35445 28040 35479
rect 27988 35436 28040 35445
rect 4423 35334 4475 35386
rect 4487 35334 4539 35386
rect 4551 35334 4603 35386
rect 4615 35334 4667 35386
rect 4679 35334 4731 35386
rect 11369 35334 11421 35386
rect 11433 35334 11485 35386
rect 11497 35334 11549 35386
rect 11561 35334 11613 35386
rect 11625 35334 11677 35386
rect 18315 35334 18367 35386
rect 18379 35334 18431 35386
rect 18443 35334 18495 35386
rect 18507 35334 18559 35386
rect 18571 35334 18623 35386
rect 25261 35334 25313 35386
rect 25325 35334 25377 35386
rect 25389 35334 25441 35386
rect 25453 35334 25505 35386
rect 25517 35334 25569 35386
rect 12716 35232 12768 35284
rect 17960 35232 18012 35284
rect 20904 35232 20956 35284
rect 21272 35275 21324 35284
rect 21272 35241 21281 35275
rect 21281 35241 21315 35275
rect 21315 35241 21324 35275
rect 21272 35232 21324 35241
rect 28080 35232 28132 35284
rect 2872 35139 2924 35148
rect 2872 35105 2881 35139
rect 2881 35105 2915 35139
rect 2915 35105 2924 35139
rect 2872 35096 2924 35105
rect 4344 35139 4396 35148
rect 4344 35105 4353 35139
rect 4353 35105 4387 35139
rect 4387 35105 4396 35139
rect 4344 35096 4396 35105
rect 1676 35071 1728 35080
rect 1676 35037 1685 35071
rect 1685 35037 1719 35071
rect 1719 35037 1728 35071
rect 1676 35028 1728 35037
rect 4252 35028 4304 35080
rect 17132 35071 17184 35080
rect 17132 35037 17166 35071
rect 17166 35037 17184 35071
rect 4344 34960 4396 35012
rect 14372 34960 14424 35012
rect 17132 35028 17184 35037
rect 18788 35028 18840 35080
rect 19524 35028 19576 35080
rect 22376 35071 22428 35080
rect 22376 35037 22394 35071
rect 22394 35037 22428 35071
rect 22376 35028 22428 35037
rect 17040 34960 17092 35012
rect 20536 34960 20588 35012
rect 23388 34960 23440 35012
rect 25044 34935 25096 34944
rect 25044 34901 25053 34935
rect 25053 34901 25087 34935
rect 25087 34901 25096 34935
rect 25044 34892 25096 34901
rect 26240 34960 26292 35012
rect 28172 34960 28224 35012
rect 26608 34892 26660 34944
rect 27712 34892 27764 34944
rect 7896 34790 7948 34842
rect 7960 34790 8012 34842
rect 8024 34790 8076 34842
rect 8088 34790 8140 34842
rect 8152 34790 8204 34842
rect 14842 34790 14894 34842
rect 14906 34790 14958 34842
rect 14970 34790 15022 34842
rect 15034 34790 15086 34842
rect 15098 34790 15150 34842
rect 21788 34790 21840 34842
rect 21852 34790 21904 34842
rect 21916 34790 21968 34842
rect 21980 34790 22032 34842
rect 22044 34790 22096 34842
rect 28734 34790 28786 34842
rect 28798 34790 28850 34842
rect 28862 34790 28914 34842
rect 28926 34790 28978 34842
rect 28990 34790 29042 34842
rect 15568 34688 15620 34740
rect 1676 34595 1728 34604
rect 1676 34561 1685 34595
rect 1685 34561 1719 34595
rect 1719 34561 1728 34595
rect 1676 34552 1728 34561
rect 4252 34552 4304 34604
rect 7748 34620 7800 34672
rect 16028 34552 16080 34604
rect 17040 34595 17092 34604
rect 17040 34561 17049 34595
rect 17049 34561 17083 34595
rect 17083 34561 17092 34595
rect 17040 34552 17092 34561
rect 17316 34595 17368 34604
rect 17316 34561 17350 34595
rect 17350 34561 17368 34595
rect 17316 34552 17368 34561
rect 17868 34688 17920 34740
rect 21180 34688 21232 34740
rect 23940 34731 23992 34740
rect 23940 34697 23949 34731
rect 23949 34697 23983 34731
rect 23983 34697 23992 34731
rect 23940 34688 23992 34697
rect 24860 34688 24912 34740
rect 25688 34688 25740 34740
rect 21272 34620 21324 34672
rect 22836 34663 22888 34672
rect 22836 34629 22870 34663
rect 22870 34629 22888 34663
rect 22836 34620 22888 34629
rect 20076 34552 20128 34604
rect 26608 34595 26660 34604
rect 26608 34561 26617 34595
rect 26617 34561 26651 34595
rect 26651 34561 26660 34595
rect 26608 34552 26660 34561
rect 27712 34595 27764 34604
rect 27712 34561 27721 34595
rect 27721 34561 27755 34595
rect 27755 34561 27764 34595
rect 27712 34552 27764 34561
rect 1860 34527 1912 34536
rect 1860 34493 1869 34527
rect 1869 34493 1903 34527
rect 1903 34493 1912 34527
rect 1860 34484 1912 34493
rect 2780 34527 2832 34536
rect 2780 34493 2789 34527
rect 2789 34493 2823 34527
rect 2823 34493 2832 34527
rect 2780 34484 2832 34493
rect 5172 34484 5224 34536
rect 5724 34484 5776 34536
rect 8392 34484 8444 34536
rect 12808 34484 12860 34536
rect 20720 34484 20772 34536
rect 22560 34527 22612 34536
rect 22560 34493 22569 34527
rect 22569 34493 22603 34527
rect 22603 34493 22612 34527
rect 22560 34484 22612 34493
rect 27804 34484 27856 34536
rect 28080 34484 28132 34536
rect 16028 34348 16080 34400
rect 20720 34348 20772 34400
rect 4423 34246 4475 34298
rect 4487 34246 4539 34298
rect 4551 34246 4603 34298
rect 4615 34246 4667 34298
rect 4679 34246 4731 34298
rect 11369 34246 11421 34298
rect 11433 34246 11485 34298
rect 11497 34246 11549 34298
rect 11561 34246 11613 34298
rect 11625 34246 11677 34298
rect 18315 34246 18367 34298
rect 18379 34246 18431 34298
rect 18443 34246 18495 34298
rect 18507 34246 18559 34298
rect 18571 34246 18623 34298
rect 25261 34246 25313 34298
rect 25325 34246 25377 34298
rect 25389 34246 25441 34298
rect 25453 34246 25505 34298
rect 25517 34246 25569 34298
rect 1860 34144 1912 34196
rect 20352 34144 20404 34196
rect 23388 34008 23440 34060
rect 27528 34051 27580 34060
rect 27528 34017 27537 34051
rect 27537 34017 27571 34051
rect 27571 34017 27580 34051
rect 27528 34008 27580 34017
rect 27988 34008 28040 34060
rect 2320 33940 2372 33992
rect 2872 33940 2924 33992
rect 4252 33940 4304 33992
rect 16028 33983 16080 33992
rect 16028 33949 16037 33983
rect 16037 33949 16071 33983
rect 16071 33949 16080 33983
rect 16028 33940 16080 33949
rect 20720 33940 20772 33992
rect 21272 33983 21324 33992
rect 21272 33949 21281 33983
rect 21281 33949 21315 33983
rect 21315 33949 21324 33983
rect 21272 33940 21324 33949
rect 23664 33983 23716 33992
rect 23664 33949 23673 33983
rect 23673 33949 23707 33983
rect 23707 33949 23716 33983
rect 23664 33940 23716 33949
rect 23756 33983 23808 33992
rect 23756 33949 23765 33983
rect 23765 33949 23799 33983
rect 23799 33949 23808 33983
rect 23756 33940 23808 33949
rect 4160 33915 4212 33924
rect 4160 33881 4169 33915
rect 4169 33881 4203 33915
rect 4203 33881 4212 33915
rect 4160 33872 4212 33881
rect 5080 33872 5132 33924
rect 21364 33872 21416 33924
rect 24124 33940 24176 33992
rect 24952 33983 25004 33992
rect 24952 33949 24986 33983
rect 24986 33949 25004 33983
rect 24952 33940 25004 33949
rect 16212 33847 16264 33856
rect 16212 33813 16221 33847
rect 16221 33813 16255 33847
rect 16255 33813 16264 33847
rect 16212 33804 16264 33813
rect 20904 33804 20956 33856
rect 23572 33804 23624 33856
rect 25136 33872 25188 33924
rect 28080 33872 28132 33924
rect 25780 33804 25832 33856
rect 25872 33804 25924 33856
rect 7896 33702 7948 33754
rect 7960 33702 8012 33754
rect 8024 33702 8076 33754
rect 8088 33702 8140 33754
rect 8152 33702 8204 33754
rect 14842 33702 14894 33754
rect 14906 33702 14958 33754
rect 14970 33702 15022 33754
rect 15034 33702 15086 33754
rect 15098 33702 15150 33754
rect 21788 33702 21840 33754
rect 21852 33702 21904 33754
rect 21916 33702 21968 33754
rect 21980 33702 22032 33754
rect 22044 33702 22096 33754
rect 28734 33702 28786 33754
rect 28798 33702 28850 33754
rect 28862 33702 28914 33754
rect 28926 33702 28978 33754
rect 28990 33702 29042 33754
rect 16580 33600 16632 33652
rect 21364 33600 21416 33652
rect 25044 33600 25096 33652
rect 16212 33532 16264 33584
rect 24124 33532 24176 33584
rect 27252 33600 27304 33652
rect 28080 33643 28132 33652
rect 28080 33609 28089 33643
rect 28089 33609 28123 33643
rect 28123 33609 28132 33643
rect 28080 33600 28132 33609
rect 15752 33507 15804 33516
rect 15752 33473 15761 33507
rect 15761 33473 15795 33507
rect 15795 33473 15804 33507
rect 15752 33464 15804 33473
rect 15844 33464 15896 33516
rect 16120 33507 16172 33516
rect 16120 33473 16129 33507
rect 16129 33473 16163 33507
rect 16163 33473 16172 33507
rect 16120 33464 16172 33473
rect 20904 33464 20956 33516
rect 21456 33464 21508 33516
rect 23480 33464 23532 33516
rect 18788 33396 18840 33448
rect 21272 33396 21324 33448
rect 22560 33396 22612 33448
rect 23388 33396 23440 33448
rect 26332 33464 26384 33516
rect 28540 33464 28592 33516
rect 28080 33396 28132 33448
rect 3516 33260 3568 33312
rect 13820 33260 13872 33312
rect 16028 33260 16080 33312
rect 23756 33260 23808 33312
rect 4423 33158 4475 33210
rect 4487 33158 4539 33210
rect 4551 33158 4603 33210
rect 4615 33158 4667 33210
rect 4679 33158 4731 33210
rect 11369 33158 11421 33210
rect 11433 33158 11485 33210
rect 11497 33158 11549 33210
rect 11561 33158 11613 33210
rect 11625 33158 11677 33210
rect 18315 33158 18367 33210
rect 18379 33158 18431 33210
rect 18443 33158 18495 33210
rect 18507 33158 18559 33210
rect 18571 33158 18623 33210
rect 25261 33158 25313 33210
rect 25325 33158 25377 33210
rect 25389 33158 25441 33210
rect 25453 33158 25505 33210
rect 25517 33158 25569 33210
rect 16764 33056 16816 33108
rect 23480 33056 23532 33108
rect 24860 33099 24912 33108
rect 24860 33065 24869 33099
rect 24869 33065 24903 33099
rect 24903 33065 24912 33099
rect 24860 33056 24912 33065
rect 15752 32988 15804 33040
rect 16488 32988 16540 33040
rect 20812 32920 20864 32972
rect 23480 32920 23532 32972
rect 23756 32920 23808 32972
rect 27528 32963 27580 32972
rect 16028 32895 16080 32904
rect 16028 32861 16037 32895
rect 16037 32861 16071 32895
rect 16071 32861 16080 32895
rect 16028 32852 16080 32861
rect 16764 32852 16816 32904
rect 17040 32784 17092 32836
rect 19984 32784 20036 32836
rect 20168 32895 20220 32904
rect 20168 32861 20177 32895
rect 20177 32861 20211 32895
rect 20211 32861 20220 32895
rect 20168 32852 20220 32861
rect 20352 32895 20404 32904
rect 20352 32861 20361 32895
rect 20361 32861 20395 32895
rect 20395 32861 20404 32895
rect 20352 32852 20404 32861
rect 23572 32895 23624 32904
rect 20260 32784 20312 32836
rect 23572 32861 23581 32895
rect 23581 32861 23615 32895
rect 23615 32861 23624 32895
rect 23572 32852 23624 32861
rect 23664 32852 23716 32904
rect 27528 32929 27537 32963
rect 27537 32929 27571 32963
rect 27571 32929 27580 32963
rect 27528 32920 27580 32929
rect 25872 32895 25924 32904
rect 16396 32716 16448 32768
rect 18880 32716 18932 32768
rect 25872 32861 25881 32895
rect 25881 32861 25915 32895
rect 25915 32861 25924 32895
rect 25872 32852 25924 32861
rect 28356 32895 28408 32904
rect 28356 32861 28365 32895
rect 28365 32861 28399 32895
rect 28399 32861 28408 32895
rect 28356 32852 28408 32861
rect 25044 32827 25096 32836
rect 25044 32793 25053 32827
rect 25053 32793 25087 32827
rect 25087 32793 25096 32827
rect 25044 32784 25096 32793
rect 28172 32827 28224 32836
rect 28172 32793 28181 32827
rect 28181 32793 28215 32827
rect 28215 32793 28224 32827
rect 28172 32784 28224 32793
rect 24216 32716 24268 32768
rect 7896 32614 7948 32666
rect 7960 32614 8012 32666
rect 8024 32614 8076 32666
rect 8088 32614 8140 32666
rect 8152 32614 8204 32666
rect 14842 32614 14894 32666
rect 14906 32614 14958 32666
rect 14970 32614 15022 32666
rect 15034 32614 15086 32666
rect 15098 32614 15150 32666
rect 21788 32614 21840 32666
rect 21852 32614 21904 32666
rect 21916 32614 21968 32666
rect 21980 32614 22032 32666
rect 22044 32614 22096 32666
rect 28734 32614 28786 32666
rect 28798 32614 28850 32666
rect 28862 32614 28914 32666
rect 28926 32614 28978 32666
rect 28990 32614 29042 32666
rect 17592 32376 17644 32428
rect 20168 32512 20220 32564
rect 21456 32444 21508 32496
rect 18880 32419 18932 32428
rect 18880 32385 18889 32419
rect 18889 32385 18923 32419
rect 18923 32385 18932 32419
rect 18880 32376 18932 32385
rect 21180 32419 21232 32428
rect 21180 32385 21189 32419
rect 21189 32385 21223 32419
rect 21223 32385 21232 32419
rect 21180 32376 21232 32385
rect 23112 32419 23164 32428
rect 12900 32351 12952 32360
rect 12900 32317 12909 32351
rect 12909 32317 12943 32351
rect 12943 32317 12952 32351
rect 12900 32308 12952 32317
rect 13820 32351 13872 32360
rect 13820 32317 13829 32351
rect 13829 32317 13863 32351
rect 13863 32317 13872 32351
rect 13820 32308 13872 32317
rect 23112 32385 23121 32419
rect 23121 32385 23155 32419
rect 23155 32385 23164 32419
rect 23112 32376 23164 32385
rect 25872 32419 25924 32428
rect 25872 32385 25881 32419
rect 25881 32385 25915 32419
rect 25915 32385 25924 32419
rect 25872 32376 25924 32385
rect 28356 32376 28408 32428
rect 13268 32240 13320 32292
rect 18880 32240 18932 32292
rect 20720 32283 20772 32292
rect 20720 32249 20729 32283
rect 20729 32249 20763 32283
rect 20763 32249 20772 32283
rect 20720 32240 20772 32249
rect 23664 32172 23716 32224
rect 25964 32215 26016 32224
rect 25964 32181 25973 32215
rect 25973 32181 26007 32215
rect 26007 32181 26016 32215
rect 25964 32172 26016 32181
rect 26608 32172 26660 32224
rect 4423 32070 4475 32122
rect 4487 32070 4539 32122
rect 4551 32070 4603 32122
rect 4615 32070 4667 32122
rect 4679 32070 4731 32122
rect 11369 32070 11421 32122
rect 11433 32070 11485 32122
rect 11497 32070 11549 32122
rect 11561 32070 11613 32122
rect 11625 32070 11677 32122
rect 18315 32070 18367 32122
rect 18379 32070 18431 32122
rect 18443 32070 18495 32122
rect 18507 32070 18559 32122
rect 18571 32070 18623 32122
rect 25261 32070 25313 32122
rect 25325 32070 25377 32122
rect 25389 32070 25441 32122
rect 25453 32070 25505 32122
rect 25517 32070 25569 32122
rect 12900 32011 12952 32020
rect 12900 31977 12909 32011
rect 12909 31977 12943 32011
rect 12943 31977 12952 32011
rect 12900 31968 12952 31977
rect 16580 31968 16632 32020
rect 19432 32011 19484 32020
rect 12808 31900 12860 31952
rect 19432 31977 19441 32011
rect 19441 31977 19475 32011
rect 19475 31977 19484 32011
rect 19432 31968 19484 31977
rect 16488 31875 16540 31884
rect 16488 31841 16497 31875
rect 16497 31841 16531 31875
rect 16531 31841 16540 31875
rect 16488 31832 16540 31841
rect 16580 31807 16632 31816
rect 16580 31773 16589 31807
rect 16589 31773 16623 31807
rect 16623 31773 16632 31807
rect 16580 31764 16632 31773
rect 17040 31764 17092 31816
rect 18604 31832 18656 31884
rect 20352 31900 20404 31952
rect 20812 31968 20864 32020
rect 22928 31968 22980 32020
rect 23112 31968 23164 32020
rect 25872 31968 25924 32020
rect 27068 31968 27120 32020
rect 28172 32011 28224 32020
rect 28172 31977 28181 32011
rect 28181 31977 28215 32011
rect 28215 31977 28224 32011
rect 28172 31968 28224 31977
rect 17592 31807 17644 31816
rect 17592 31773 17601 31807
rect 17601 31773 17635 31807
rect 17635 31773 17644 31807
rect 17592 31764 17644 31773
rect 16856 31696 16908 31748
rect 19616 31696 19668 31748
rect 19892 31807 19944 31816
rect 19892 31773 19901 31807
rect 19901 31773 19935 31807
rect 19935 31773 19944 31807
rect 19892 31764 19944 31773
rect 20076 31807 20128 31816
rect 20076 31773 20085 31807
rect 20085 31773 20119 31807
rect 20119 31773 20128 31807
rect 20076 31764 20128 31773
rect 20352 31764 20404 31816
rect 21272 31764 21324 31816
rect 22192 31764 22244 31816
rect 24308 31900 24360 31952
rect 23664 31875 23716 31884
rect 23664 31841 23673 31875
rect 23673 31841 23707 31875
rect 23707 31841 23716 31875
rect 23664 31832 23716 31841
rect 25780 31875 25832 31884
rect 25780 31841 25789 31875
rect 25789 31841 25823 31875
rect 25823 31841 25832 31875
rect 25780 31832 25832 31841
rect 25964 31875 26016 31884
rect 25964 31841 25973 31875
rect 25973 31841 26007 31875
rect 26007 31841 26016 31875
rect 25964 31832 26016 31841
rect 27528 31875 27580 31884
rect 27528 31841 27537 31875
rect 27537 31841 27571 31875
rect 27571 31841 27580 31875
rect 27528 31832 27580 31841
rect 23572 31807 23624 31816
rect 23572 31773 23581 31807
rect 23581 31773 23615 31807
rect 23615 31773 23624 31807
rect 23572 31764 23624 31773
rect 27896 31764 27948 31816
rect 28172 31764 28224 31816
rect 23940 31696 23992 31748
rect 24952 31739 25004 31748
rect 24952 31705 24961 31739
rect 24961 31705 24995 31739
rect 24995 31705 25004 31739
rect 24952 31696 25004 31705
rect 22560 31628 22612 31680
rect 23204 31671 23256 31680
rect 23204 31637 23213 31671
rect 23213 31637 23247 31671
rect 23247 31637 23256 31671
rect 23204 31628 23256 31637
rect 7896 31526 7948 31578
rect 7960 31526 8012 31578
rect 8024 31526 8076 31578
rect 8088 31526 8140 31578
rect 8152 31526 8204 31578
rect 14842 31526 14894 31578
rect 14906 31526 14958 31578
rect 14970 31526 15022 31578
rect 15034 31526 15086 31578
rect 15098 31526 15150 31578
rect 21788 31526 21840 31578
rect 21852 31526 21904 31578
rect 21916 31526 21968 31578
rect 21980 31526 22032 31578
rect 22044 31526 22096 31578
rect 28734 31526 28786 31578
rect 28798 31526 28850 31578
rect 28862 31526 28914 31578
rect 28926 31526 28978 31578
rect 28990 31526 29042 31578
rect 16212 31424 16264 31476
rect 16672 31424 16724 31476
rect 22192 31424 22244 31476
rect 23204 31467 23256 31476
rect 23204 31433 23213 31467
rect 23213 31433 23247 31467
rect 23247 31433 23256 31467
rect 23204 31424 23256 31433
rect 23572 31424 23624 31476
rect 18604 31399 18656 31408
rect 18604 31365 18622 31399
rect 18622 31365 18656 31399
rect 18604 31356 18656 31365
rect 22468 31356 22520 31408
rect 22928 31399 22980 31408
rect 22928 31365 22937 31399
rect 22937 31365 22971 31399
rect 22971 31365 22980 31399
rect 22928 31356 22980 31365
rect 24216 31399 24268 31408
rect 24216 31365 24225 31399
rect 24225 31365 24259 31399
rect 24259 31365 24268 31399
rect 24216 31356 24268 31365
rect 16764 31288 16816 31340
rect 17224 31288 17276 31340
rect 21088 31288 21140 31340
rect 21640 31288 21692 31340
rect 22560 31288 22612 31340
rect 22836 31331 22888 31340
rect 18880 31263 18932 31272
rect 16580 31152 16632 31204
rect 18880 31229 18889 31263
rect 18889 31229 18923 31263
rect 18923 31229 18932 31263
rect 18880 31220 18932 31229
rect 22836 31297 22845 31331
rect 22845 31297 22879 31331
rect 22879 31297 22888 31331
rect 22836 31288 22888 31297
rect 23112 31288 23164 31340
rect 23940 31288 23992 31340
rect 26608 31331 26660 31340
rect 26608 31297 26617 31331
rect 26617 31297 26651 31331
rect 26651 31297 26660 31331
rect 26608 31288 26660 31297
rect 27620 31288 27672 31340
rect 23388 31220 23440 31272
rect 26148 31263 26200 31272
rect 26148 31229 26157 31263
rect 26157 31229 26191 31263
rect 26191 31229 26200 31263
rect 26148 31220 26200 31229
rect 16672 31084 16724 31136
rect 19892 31084 19944 31136
rect 20076 31084 20128 31136
rect 4423 30982 4475 31034
rect 4487 30982 4539 31034
rect 4551 30982 4603 31034
rect 4615 30982 4667 31034
rect 4679 30982 4731 31034
rect 11369 30982 11421 31034
rect 11433 30982 11485 31034
rect 11497 30982 11549 31034
rect 11561 30982 11613 31034
rect 11625 30982 11677 31034
rect 18315 30982 18367 31034
rect 18379 30982 18431 31034
rect 18443 30982 18495 31034
rect 18507 30982 18559 31034
rect 18571 30982 18623 31034
rect 25261 30982 25313 31034
rect 25325 30982 25377 31034
rect 25389 30982 25441 31034
rect 25453 30982 25505 31034
rect 25517 30982 25569 31034
rect 15844 30880 15896 30932
rect 22836 30880 22888 30932
rect 23112 30923 23164 30932
rect 23112 30889 23121 30923
rect 23121 30889 23155 30923
rect 23155 30889 23164 30923
rect 23112 30880 23164 30889
rect 24952 30880 25004 30932
rect 16304 30744 16356 30796
rect 16672 30719 16724 30728
rect 16672 30685 16681 30719
rect 16681 30685 16715 30719
rect 16715 30685 16724 30719
rect 16672 30676 16724 30685
rect 19340 30676 19392 30728
rect 22468 30719 22520 30728
rect 22468 30685 22477 30719
rect 22477 30685 22511 30719
rect 22511 30685 22520 30719
rect 22468 30676 22520 30685
rect 23940 30744 23992 30796
rect 28264 30787 28316 30796
rect 28264 30753 28273 30787
rect 28273 30753 28307 30787
rect 28307 30753 28316 30787
rect 28264 30744 28316 30753
rect 23388 30719 23440 30728
rect 23388 30685 23397 30719
rect 23397 30685 23431 30719
rect 23431 30685 23440 30719
rect 23388 30676 23440 30685
rect 23572 30676 23624 30728
rect 24860 30719 24912 30728
rect 24860 30685 24869 30719
rect 24869 30685 24903 30719
rect 24903 30685 24912 30719
rect 24860 30676 24912 30685
rect 26332 30676 26384 30728
rect 21640 30608 21692 30660
rect 23664 30651 23716 30660
rect 23664 30617 23673 30651
rect 23673 30617 23707 30651
rect 23707 30617 23716 30651
rect 23664 30608 23716 30617
rect 23756 30651 23808 30660
rect 23756 30617 23765 30651
rect 23765 30617 23799 30651
rect 23799 30617 23808 30651
rect 23756 30608 23808 30617
rect 17224 30540 17276 30592
rect 23112 30540 23164 30592
rect 25136 30608 25188 30660
rect 26608 30651 26660 30660
rect 24584 30583 24636 30592
rect 24584 30549 24593 30583
rect 24593 30549 24627 30583
rect 24627 30549 24636 30583
rect 24584 30540 24636 30549
rect 24768 30540 24820 30592
rect 26608 30617 26617 30651
rect 26617 30617 26651 30651
rect 26651 30617 26660 30651
rect 26608 30608 26660 30617
rect 7896 30438 7948 30490
rect 7960 30438 8012 30490
rect 8024 30438 8076 30490
rect 8088 30438 8140 30490
rect 8152 30438 8204 30490
rect 14842 30438 14894 30490
rect 14906 30438 14958 30490
rect 14970 30438 15022 30490
rect 15034 30438 15086 30490
rect 15098 30438 15150 30490
rect 21788 30438 21840 30490
rect 21852 30438 21904 30490
rect 21916 30438 21968 30490
rect 21980 30438 22032 30490
rect 22044 30438 22096 30490
rect 28734 30438 28786 30490
rect 28798 30438 28850 30490
rect 28862 30438 28914 30490
rect 28926 30438 28978 30490
rect 28990 30438 29042 30490
rect 19340 30336 19392 30388
rect 16672 30268 16724 30320
rect 16856 30268 16908 30320
rect 19892 30268 19944 30320
rect 16304 30243 16356 30252
rect 16304 30209 16313 30243
rect 16313 30209 16347 30243
rect 16347 30209 16356 30243
rect 16304 30200 16356 30209
rect 17040 30243 17092 30252
rect 17040 30209 17049 30243
rect 17049 30209 17083 30243
rect 17083 30209 17092 30243
rect 17040 30200 17092 30209
rect 17224 30243 17276 30252
rect 17224 30209 17233 30243
rect 17233 30209 17267 30243
rect 17267 30209 17276 30243
rect 17224 30200 17276 30209
rect 17500 30243 17552 30252
rect 17500 30209 17509 30243
rect 17509 30209 17543 30243
rect 17543 30209 17552 30243
rect 17500 30200 17552 30209
rect 21088 30336 21140 30388
rect 24216 30336 24268 30388
rect 21640 30268 21692 30320
rect 23296 30268 23348 30320
rect 24860 30268 24912 30320
rect 1584 30175 1636 30184
rect 1584 30141 1593 30175
rect 1593 30141 1627 30175
rect 1627 30141 1636 30175
rect 1584 30132 1636 30141
rect 1860 30175 1912 30184
rect 1860 30141 1869 30175
rect 1869 30141 1903 30175
rect 1903 30141 1912 30175
rect 1860 30132 1912 30141
rect 15844 30132 15896 30184
rect 20076 30200 20128 30252
rect 22284 30243 22336 30252
rect 22284 30209 22293 30243
rect 22293 30209 22327 30243
rect 22327 30209 22336 30243
rect 22284 30200 22336 30209
rect 22468 30200 22520 30252
rect 24216 30200 24268 30252
rect 24584 30200 24636 30252
rect 25964 30200 26016 30252
rect 26148 30243 26200 30252
rect 26148 30209 26157 30243
rect 26157 30209 26191 30243
rect 26191 30209 26200 30243
rect 26608 30336 26660 30388
rect 26148 30200 26200 30209
rect 26976 30200 27028 30252
rect 27160 30200 27212 30252
rect 28356 30243 28408 30252
rect 28356 30209 28365 30243
rect 28365 30209 28399 30243
rect 28399 30209 28408 30243
rect 28356 30200 28408 30209
rect 23204 30132 23256 30184
rect 22744 30064 22796 30116
rect 23664 30064 23716 30116
rect 24308 30107 24360 30116
rect 16856 30039 16908 30048
rect 16856 30005 16865 30039
rect 16865 30005 16899 30039
rect 16899 30005 16908 30039
rect 16856 29996 16908 30005
rect 19524 29996 19576 30048
rect 22008 30039 22060 30048
rect 22008 30005 22017 30039
rect 22017 30005 22051 30039
rect 22051 30005 22060 30039
rect 22008 29996 22060 30005
rect 23296 30039 23348 30048
rect 23296 30005 23305 30039
rect 23305 30005 23339 30039
rect 23339 30005 23348 30039
rect 23296 29996 23348 30005
rect 23756 29996 23808 30048
rect 24308 30073 24317 30107
rect 24317 30073 24351 30107
rect 24351 30073 24360 30107
rect 24308 30064 24360 30073
rect 24768 30132 24820 30184
rect 26516 30132 26568 30184
rect 26056 30064 26108 30116
rect 28080 30064 28132 30116
rect 24952 30039 25004 30048
rect 24952 30005 24961 30039
rect 24961 30005 24995 30039
rect 24995 30005 25004 30039
rect 24952 29996 25004 30005
rect 26240 29996 26292 30048
rect 4423 29894 4475 29946
rect 4487 29894 4539 29946
rect 4551 29894 4603 29946
rect 4615 29894 4667 29946
rect 4679 29894 4731 29946
rect 11369 29894 11421 29946
rect 11433 29894 11485 29946
rect 11497 29894 11549 29946
rect 11561 29894 11613 29946
rect 11625 29894 11677 29946
rect 18315 29894 18367 29946
rect 18379 29894 18431 29946
rect 18443 29894 18495 29946
rect 18507 29894 18559 29946
rect 18571 29894 18623 29946
rect 25261 29894 25313 29946
rect 25325 29894 25377 29946
rect 25389 29894 25441 29946
rect 25453 29894 25505 29946
rect 25517 29894 25569 29946
rect 16672 29792 16724 29844
rect 17500 29792 17552 29844
rect 17776 29792 17828 29844
rect 20352 29792 20404 29844
rect 21088 29792 21140 29844
rect 24952 29835 25004 29844
rect 24952 29801 24961 29835
rect 24961 29801 24995 29835
rect 24995 29801 25004 29835
rect 24952 29792 25004 29801
rect 26516 29792 26568 29844
rect 23756 29724 23808 29776
rect 26148 29724 26200 29776
rect 17592 29656 17644 29708
rect 24032 29656 24084 29708
rect 27528 29699 27580 29708
rect 27528 29665 27537 29699
rect 27537 29665 27571 29699
rect 27571 29665 27580 29699
rect 27528 29656 27580 29665
rect 16856 29631 16908 29640
rect 16856 29597 16865 29631
rect 16865 29597 16899 29631
rect 16899 29597 16908 29631
rect 16856 29588 16908 29597
rect 18880 29588 18932 29640
rect 19524 29588 19576 29640
rect 21180 29588 21232 29640
rect 22652 29631 22704 29640
rect 22652 29597 22661 29631
rect 22661 29597 22695 29631
rect 22695 29597 22704 29631
rect 22652 29588 22704 29597
rect 24584 29631 24636 29640
rect 24584 29597 24593 29631
rect 24593 29597 24627 29631
rect 24627 29597 24636 29631
rect 24584 29588 24636 29597
rect 25872 29631 25924 29640
rect 25872 29597 25881 29631
rect 25881 29597 25915 29631
rect 25915 29597 25924 29631
rect 25872 29588 25924 29597
rect 26056 29631 26108 29640
rect 26056 29597 26065 29631
rect 26065 29597 26099 29631
rect 26099 29597 26108 29631
rect 26516 29631 26568 29640
rect 26056 29588 26108 29597
rect 26516 29597 26525 29631
rect 26525 29597 26559 29631
rect 26559 29597 26568 29631
rect 26516 29588 26568 29597
rect 22008 29520 22060 29572
rect 21272 29495 21324 29504
rect 21272 29461 21281 29495
rect 21281 29461 21315 29495
rect 21315 29461 21324 29495
rect 21272 29452 21324 29461
rect 22192 29452 22244 29504
rect 25044 29452 25096 29504
rect 27344 29520 27396 29572
rect 27068 29452 27120 29504
rect 7896 29350 7948 29402
rect 7960 29350 8012 29402
rect 8024 29350 8076 29402
rect 8088 29350 8140 29402
rect 8152 29350 8204 29402
rect 14842 29350 14894 29402
rect 14906 29350 14958 29402
rect 14970 29350 15022 29402
rect 15034 29350 15086 29402
rect 15098 29350 15150 29402
rect 21788 29350 21840 29402
rect 21852 29350 21904 29402
rect 21916 29350 21968 29402
rect 21980 29350 22032 29402
rect 22044 29350 22096 29402
rect 28734 29350 28786 29402
rect 28798 29350 28850 29402
rect 28862 29350 28914 29402
rect 28926 29350 28978 29402
rect 28990 29350 29042 29402
rect 20260 29248 20312 29300
rect 22284 29248 22336 29300
rect 23204 29291 23256 29300
rect 23204 29257 23213 29291
rect 23213 29257 23247 29291
rect 23247 29257 23256 29291
rect 23204 29248 23256 29257
rect 23664 29248 23716 29300
rect 25964 29291 26016 29300
rect 25964 29257 25973 29291
rect 25973 29257 26007 29291
rect 26007 29257 26016 29291
rect 25964 29248 26016 29257
rect 27344 29291 27396 29300
rect 27344 29257 27353 29291
rect 27353 29257 27387 29291
rect 27387 29257 27396 29291
rect 27344 29248 27396 29257
rect 4804 29180 4856 29232
rect 20812 29180 20864 29232
rect 20076 29112 20128 29164
rect 21272 29044 21324 29096
rect 22192 29112 22244 29164
rect 22284 29112 22336 29164
rect 23204 29112 23256 29164
rect 23480 29112 23532 29164
rect 22744 29044 22796 29096
rect 22192 28976 22244 29028
rect 24952 29112 25004 29164
rect 26608 29112 26660 29164
rect 27068 29112 27120 29164
rect 18880 28908 18932 28960
rect 23756 28908 23808 28960
rect 25872 29044 25924 29096
rect 26056 28976 26108 29028
rect 26516 28976 26568 29028
rect 4423 28806 4475 28858
rect 4487 28806 4539 28858
rect 4551 28806 4603 28858
rect 4615 28806 4667 28858
rect 4679 28806 4731 28858
rect 11369 28806 11421 28858
rect 11433 28806 11485 28858
rect 11497 28806 11549 28858
rect 11561 28806 11613 28858
rect 11625 28806 11677 28858
rect 18315 28806 18367 28858
rect 18379 28806 18431 28858
rect 18443 28806 18495 28858
rect 18507 28806 18559 28858
rect 18571 28806 18623 28858
rect 25261 28806 25313 28858
rect 25325 28806 25377 28858
rect 25389 28806 25441 28858
rect 25453 28806 25505 28858
rect 25517 28806 25569 28858
rect 16028 28704 16080 28756
rect 24676 28747 24728 28756
rect 24676 28713 24685 28747
rect 24685 28713 24719 28747
rect 24719 28713 24728 28747
rect 24676 28704 24728 28713
rect 22652 28568 22704 28620
rect 25136 28568 25188 28620
rect 26516 28611 26568 28620
rect 26516 28577 26525 28611
rect 26525 28577 26559 28611
rect 26559 28577 26568 28611
rect 26516 28568 26568 28577
rect 27436 28611 27488 28620
rect 27436 28577 27445 28611
rect 27445 28577 27479 28611
rect 27479 28577 27488 28611
rect 27436 28568 27488 28577
rect 18880 28500 18932 28552
rect 20812 28543 20864 28552
rect 20812 28509 20821 28543
rect 20821 28509 20855 28543
rect 20855 28509 20864 28543
rect 20812 28500 20864 28509
rect 22560 28500 22612 28552
rect 23388 28500 23440 28552
rect 15660 28475 15712 28484
rect 15660 28441 15669 28475
rect 15669 28441 15703 28475
rect 15703 28441 15712 28475
rect 15660 28432 15712 28441
rect 15752 28432 15804 28484
rect 16764 28364 16816 28416
rect 17040 28432 17092 28484
rect 22468 28432 22520 28484
rect 23940 28432 23992 28484
rect 27344 28432 27396 28484
rect 19340 28364 19392 28416
rect 22652 28364 22704 28416
rect 23204 28407 23256 28416
rect 23204 28373 23213 28407
rect 23213 28373 23247 28407
rect 23247 28373 23256 28407
rect 23204 28364 23256 28373
rect 24492 28364 24544 28416
rect 7896 28262 7948 28314
rect 7960 28262 8012 28314
rect 8024 28262 8076 28314
rect 8088 28262 8140 28314
rect 8152 28262 8204 28314
rect 14842 28262 14894 28314
rect 14906 28262 14958 28314
rect 14970 28262 15022 28314
rect 15034 28262 15086 28314
rect 15098 28262 15150 28314
rect 21788 28262 21840 28314
rect 21852 28262 21904 28314
rect 21916 28262 21968 28314
rect 21980 28262 22032 28314
rect 22044 28262 22096 28314
rect 28734 28262 28786 28314
rect 28798 28262 28850 28314
rect 28862 28262 28914 28314
rect 28926 28262 28978 28314
rect 28990 28262 29042 28314
rect 17040 28203 17092 28212
rect 17040 28169 17049 28203
rect 17049 28169 17083 28203
rect 17083 28169 17092 28203
rect 17040 28160 17092 28169
rect 22468 28203 22520 28212
rect 22468 28169 22477 28203
rect 22477 28169 22511 28203
rect 22511 28169 22520 28203
rect 22468 28160 22520 28169
rect 23388 28203 23440 28212
rect 23388 28169 23397 28203
rect 23397 28169 23431 28203
rect 23431 28169 23440 28203
rect 23388 28160 23440 28169
rect 27344 28203 27396 28212
rect 27344 28169 27353 28203
rect 27353 28169 27387 28203
rect 27387 28169 27396 28203
rect 27344 28160 27396 28169
rect 23664 28092 23716 28144
rect 23756 28135 23808 28144
rect 23756 28101 23765 28135
rect 23765 28101 23799 28135
rect 23799 28101 23808 28135
rect 23756 28092 23808 28101
rect 1584 28067 1636 28076
rect 1584 28033 1593 28067
rect 1593 28033 1627 28067
rect 1627 28033 1636 28067
rect 1584 28024 1636 28033
rect 16764 28024 16816 28076
rect 19340 28024 19392 28076
rect 22192 28067 22244 28076
rect 2964 27956 3016 28008
rect 15200 27956 15252 28008
rect 20260 27956 20312 28008
rect 22192 28033 22201 28067
rect 22201 28033 22235 28067
rect 22235 28033 22244 28067
rect 22192 28024 22244 28033
rect 22284 28067 22336 28076
rect 22284 28033 22293 28067
rect 22293 28033 22327 28067
rect 22327 28033 22336 28067
rect 22284 28024 22336 28033
rect 24124 28024 24176 28076
rect 24492 28067 24544 28076
rect 24492 28033 24501 28067
rect 24501 28033 24535 28067
rect 24535 28033 24544 28067
rect 24492 28024 24544 28033
rect 26240 28092 26292 28144
rect 25780 28024 25832 28076
rect 27252 28024 27304 28076
rect 27988 28024 28040 28076
rect 24400 27999 24452 28008
rect 24400 27965 24409 27999
rect 24409 27965 24443 27999
rect 24443 27965 24452 27999
rect 24400 27956 24452 27965
rect 25136 27956 25188 28008
rect 1768 27863 1820 27872
rect 1768 27829 1777 27863
rect 1777 27829 1811 27863
rect 1811 27829 1820 27863
rect 1768 27820 1820 27829
rect 24492 27820 24544 27872
rect 24768 27863 24820 27872
rect 24768 27829 24777 27863
rect 24777 27829 24811 27863
rect 24811 27829 24820 27863
rect 24768 27820 24820 27829
rect 25596 27820 25648 27872
rect 26608 27863 26660 27872
rect 26608 27829 26617 27863
rect 26617 27829 26651 27863
rect 26651 27829 26660 27863
rect 26608 27820 26660 27829
rect 28080 27863 28132 27872
rect 28080 27829 28089 27863
rect 28089 27829 28123 27863
rect 28123 27829 28132 27863
rect 28080 27820 28132 27829
rect 4423 27718 4475 27770
rect 4487 27718 4539 27770
rect 4551 27718 4603 27770
rect 4615 27718 4667 27770
rect 4679 27718 4731 27770
rect 11369 27718 11421 27770
rect 11433 27718 11485 27770
rect 11497 27718 11549 27770
rect 11561 27718 11613 27770
rect 11625 27718 11677 27770
rect 18315 27718 18367 27770
rect 18379 27718 18431 27770
rect 18443 27718 18495 27770
rect 18507 27718 18559 27770
rect 18571 27718 18623 27770
rect 25261 27718 25313 27770
rect 25325 27718 25377 27770
rect 25389 27718 25441 27770
rect 25453 27718 25505 27770
rect 25517 27718 25569 27770
rect 15660 27616 15712 27668
rect 24492 27616 24544 27668
rect 25780 27659 25832 27668
rect 2596 27548 2648 27600
rect 4988 27548 5040 27600
rect 15200 27548 15252 27600
rect 21456 27548 21508 27600
rect 22192 27548 22244 27600
rect 25136 27548 25188 27600
rect 25780 27625 25789 27659
rect 25789 27625 25823 27659
rect 25823 27625 25832 27659
rect 25780 27616 25832 27625
rect 26608 27616 26660 27668
rect 15844 27480 15896 27532
rect 27528 27523 27580 27532
rect 14372 27455 14424 27464
rect 14372 27421 14381 27455
rect 14381 27421 14415 27455
rect 14415 27421 14424 27455
rect 14372 27412 14424 27421
rect 16028 27412 16080 27464
rect 16304 27412 16356 27464
rect 18880 27412 18932 27464
rect 24952 27412 25004 27464
rect 27528 27489 27537 27523
rect 27537 27489 27571 27523
rect 27571 27489 27580 27523
rect 27528 27480 27580 27489
rect 28080 27480 28132 27532
rect 1768 27344 1820 27396
rect 19800 27344 19852 27396
rect 23204 27344 23256 27396
rect 25044 27344 25096 27396
rect 25596 27344 25648 27396
rect 27804 27344 27856 27396
rect 17132 27276 17184 27328
rect 21088 27276 21140 27328
rect 22284 27276 22336 27328
rect 7896 27174 7948 27226
rect 7960 27174 8012 27226
rect 8024 27174 8076 27226
rect 8088 27174 8140 27226
rect 8152 27174 8204 27226
rect 14842 27174 14894 27226
rect 14906 27174 14958 27226
rect 14970 27174 15022 27226
rect 15034 27174 15086 27226
rect 15098 27174 15150 27226
rect 21788 27174 21840 27226
rect 21852 27174 21904 27226
rect 21916 27174 21968 27226
rect 21980 27174 22032 27226
rect 22044 27174 22096 27226
rect 28734 27174 28786 27226
rect 28798 27174 28850 27226
rect 28862 27174 28914 27226
rect 28926 27174 28978 27226
rect 28990 27174 29042 27226
rect 16304 27115 16356 27124
rect 16304 27081 16313 27115
rect 16313 27081 16347 27115
rect 16347 27081 16356 27115
rect 16304 27072 16356 27081
rect 20260 27115 20312 27124
rect 20260 27081 20269 27115
rect 20269 27081 20303 27115
rect 20303 27081 20312 27115
rect 20260 27072 20312 27081
rect 15936 26979 15988 26988
rect 15936 26945 15945 26979
rect 15945 26945 15979 26979
rect 15979 26945 15988 26979
rect 15936 26936 15988 26945
rect 16764 26868 16816 26920
rect 16856 26868 16908 26920
rect 17132 26936 17184 26988
rect 20720 27004 20772 27056
rect 21640 27072 21692 27124
rect 23204 27115 23256 27124
rect 23204 27081 23213 27115
rect 23213 27081 23247 27115
rect 23247 27081 23256 27115
rect 23204 27072 23256 27081
rect 24492 27115 24544 27124
rect 24492 27081 24501 27115
rect 24501 27081 24535 27115
rect 24535 27081 24544 27115
rect 24492 27072 24544 27081
rect 27804 27115 27856 27124
rect 27804 27081 27813 27115
rect 27813 27081 27847 27115
rect 27847 27081 27856 27115
rect 27804 27072 27856 27081
rect 22928 27004 22980 27056
rect 23756 27004 23808 27056
rect 18880 26979 18932 26988
rect 18880 26945 18889 26979
rect 18889 26945 18923 26979
rect 18923 26945 18932 26979
rect 18880 26936 18932 26945
rect 18972 26936 19024 26988
rect 23296 26979 23348 26988
rect 22008 26911 22060 26920
rect 22008 26877 22017 26911
rect 22017 26877 22051 26911
rect 22051 26877 22060 26911
rect 22008 26868 22060 26877
rect 22376 26911 22428 26920
rect 22376 26877 22385 26911
rect 22385 26877 22419 26911
rect 22419 26877 22428 26911
rect 22376 26868 22428 26877
rect 22744 26868 22796 26920
rect 22192 26800 22244 26852
rect 23296 26945 23305 26979
rect 23305 26945 23339 26979
rect 23339 26945 23348 26979
rect 23296 26936 23348 26945
rect 23664 26936 23716 26988
rect 24124 26936 24176 26988
rect 24492 26936 24544 26988
rect 27712 26979 27764 26988
rect 27712 26945 27721 26979
rect 27721 26945 27755 26979
rect 27755 26945 27764 26979
rect 27712 26936 27764 26945
rect 28264 26936 28316 26988
rect 24676 26843 24728 26852
rect 24676 26809 24685 26843
rect 24685 26809 24719 26843
rect 24719 26809 24728 26843
rect 24676 26800 24728 26809
rect 18236 26732 18288 26784
rect 19616 26732 19668 26784
rect 21180 26775 21232 26784
rect 21180 26741 21189 26775
rect 21189 26741 21223 26775
rect 21223 26741 21232 26775
rect 21180 26732 21232 26741
rect 4423 26630 4475 26682
rect 4487 26630 4539 26682
rect 4551 26630 4603 26682
rect 4615 26630 4667 26682
rect 4679 26630 4731 26682
rect 11369 26630 11421 26682
rect 11433 26630 11485 26682
rect 11497 26630 11549 26682
rect 11561 26630 11613 26682
rect 11625 26630 11677 26682
rect 18315 26630 18367 26682
rect 18379 26630 18431 26682
rect 18443 26630 18495 26682
rect 18507 26630 18559 26682
rect 18571 26630 18623 26682
rect 25261 26630 25313 26682
rect 25325 26630 25377 26682
rect 25389 26630 25441 26682
rect 25453 26630 25505 26682
rect 25517 26630 25569 26682
rect 15936 26528 15988 26580
rect 19800 26571 19852 26580
rect 19800 26537 19809 26571
rect 19809 26537 19843 26571
rect 19843 26537 19852 26571
rect 19800 26528 19852 26537
rect 20904 26528 20956 26580
rect 22008 26571 22060 26580
rect 22008 26537 22017 26571
rect 22017 26537 22051 26571
rect 22051 26537 22060 26571
rect 22008 26528 22060 26537
rect 24032 26571 24084 26580
rect 24032 26537 24041 26571
rect 24041 26537 24075 26571
rect 24075 26537 24084 26571
rect 24032 26528 24084 26537
rect 24676 26528 24728 26580
rect 24124 26460 24176 26512
rect 15476 26392 15528 26444
rect 18880 26392 18932 26444
rect 2596 26324 2648 26376
rect 18236 26324 18288 26376
rect 19984 26367 20036 26376
rect 19984 26333 19993 26367
rect 19993 26333 20027 26367
rect 20027 26333 20036 26367
rect 19984 26324 20036 26333
rect 21180 26324 21232 26376
rect 23940 26324 23992 26376
rect 24124 26324 24176 26376
rect 25136 26324 25188 26376
rect 15752 26299 15804 26308
rect 15752 26265 15761 26299
rect 15761 26265 15795 26299
rect 15795 26265 15804 26299
rect 15752 26256 15804 26265
rect 26240 26256 26292 26308
rect 1860 26188 1912 26240
rect 25504 26188 25556 26240
rect 25964 26231 26016 26240
rect 25964 26197 25973 26231
rect 25973 26197 26007 26231
rect 26007 26197 26016 26231
rect 25964 26188 26016 26197
rect 7896 26086 7948 26138
rect 7960 26086 8012 26138
rect 8024 26086 8076 26138
rect 8088 26086 8140 26138
rect 8152 26086 8204 26138
rect 14842 26086 14894 26138
rect 14906 26086 14958 26138
rect 14970 26086 15022 26138
rect 15034 26086 15086 26138
rect 15098 26086 15150 26138
rect 21788 26086 21840 26138
rect 21852 26086 21904 26138
rect 21916 26086 21968 26138
rect 21980 26086 22032 26138
rect 22044 26086 22096 26138
rect 28734 26086 28786 26138
rect 28798 26086 28850 26138
rect 28862 26086 28914 26138
rect 28926 26086 28978 26138
rect 28990 26086 29042 26138
rect 1860 25959 1912 25968
rect 1860 25925 1869 25959
rect 1869 25925 1903 25959
rect 1903 25925 1912 25959
rect 1860 25916 1912 25925
rect 16488 25984 16540 26036
rect 19708 25984 19760 26036
rect 19984 25984 20036 26036
rect 22928 26027 22980 26036
rect 22928 25993 22937 26027
rect 22937 25993 22971 26027
rect 22971 25993 22980 26027
rect 22928 25984 22980 25993
rect 25596 25984 25648 26036
rect 27068 25984 27120 26036
rect 27436 25984 27488 26036
rect 16120 25891 16172 25900
rect 16120 25857 16129 25891
rect 16129 25857 16163 25891
rect 16163 25857 16172 25891
rect 16120 25848 16172 25857
rect 19984 25891 20036 25900
rect 19984 25857 19993 25891
rect 19993 25857 20027 25891
rect 20027 25857 20036 25891
rect 19984 25848 20036 25857
rect 20168 25891 20220 25900
rect 20168 25857 20177 25891
rect 20177 25857 20211 25891
rect 20211 25857 20220 25891
rect 20168 25848 20220 25857
rect 22652 25848 22704 25900
rect 26056 25916 26108 25968
rect 25504 25891 25556 25900
rect 1676 25823 1728 25832
rect 1676 25789 1685 25823
rect 1685 25789 1719 25823
rect 1719 25789 1728 25823
rect 1676 25780 1728 25789
rect 2780 25823 2832 25832
rect 2780 25789 2789 25823
rect 2789 25789 2823 25823
rect 2823 25789 2832 25823
rect 2780 25780 2832 25789
rect 16856 25823 16908 25832
rect 16856 25789 16865 25823
rect 16865 25789 16899 25823
rect 16899 25789 16908 25823
rect 16856 25780 16908 25789
rect 25504 25857 25513 25891
rect 25513 25857 25547 25891
rect 25547 25857 25556 25891
rect 25504 25848 25556 25857
rect 25964 25848 26016 25900
rect 26976 25848 27028 25900
rect 21732 25644 21784 25696
rect 23664 25712 23716 25764
rect 26148 25823 26200 25832
rect 26148 25789 26157 25823
rect 26157 25789 26191 25823
rect 26191 25789 26200 25823
rect 26148 25780 26200 25789
rect 25872 25712 25924 25764
rect 25688 25644 25740 25696
rect 25780 25644 25832 25696
rect 4423 25542 4475 25594
rect 4487 25542 4539 25594
rect 4551 25542 4603 25594
rect 4615 25542 4667 25594
rect 4679 25542 4731 25594
rect 11369 25542 11421 25594
rect 11433 25542 11485 25594
rect 11497 25542 11549 25594
rect 11561 25542 11613 25594
rect 11625 25542 11677 25594
rect 18315 25542 18367 25594
rect 18379 25542 18431 25594
rect 18443 25542 18495 25594
rect 18507 25542 18559 25594
rect 18571 25542 18623 25594
rect 25261 25542 25313 25594
rect 25325 25542 25377 25594
rect 25389 25542 25441 25594
rect 25453 25542 25505 25594
rect 25517 25542 25569 25594
rect 1676 25483 1728 25492
rect 1676 25449 1685 25483
rect 1685 25449 1719 25483
rect 1719 25449 1728 25483
rect 1676 25440 1728 25449
rect 16120 25440 16172 25492
rect 18972 25440 19024 25492
rect 26240 25440 26292 25492
rect 22376 25372 22428 25424
rect 15476 25304 15528 25356
rect 24952 25304 25004 25356
rect 25688 25304 25740 25356
rect 27712 25304 27764 25356
rect 16488 25236 16540 25288
rect 18236 25236 18288 25288
rect 9496 25100 9548 25152
rect 16764 25168 16816 25220
rect 17132 25168 17184 25220
rect 20720 25236 20772 25288
rect 21456 25236 21508 25288
rect 21732 25279 21784 25288
rect 21732 25245 21741 25279
rect 21741 25245 21775 25279
rect 21775 25245 21784 25279
rect 21732 25236 21784 25245
rect 22836 25236 22888 25288
rect 24860 25236 24912 25288
rect 25044 25279 25096 25288
rect 25044 25245 25053 25279
rect 25053 25245 25087 25279
rect 25087 25245 25096 25279
rect 25044 25236 25096 25245
rect 25228 25279 25280 25288
rect 25228 25245 25237 25279
rect 25237 25245 25271 25279
rect 25271 25245 25280 25279
rect 25228 25236 25280 25245
rect 25596 25279 25648 25288
rect 25596 25245 25605 25279
rect 25605 25245 25639 25279
rect 25639 25245 25648 25279
rect 25596 25236 25648 25245
rect 25964 25236 26016 25288
rect 24216 25168 24268 25220
rect 26700 25211 26752 25220
rect 26700 25177 26709 25211
rect 26709 25177 26743 25211
rect 26743 25177 26752 25211
rect 26700 25168 26752 25177
rect 28356 25211 28408 25220
rect 28356 25177 28365 25211
rect 28365 25177 28399 25211
rect 28399 25177 28408 25211
rect 28356 25168 28408 25177
rect 22560 25143 22612 25152
rect 22560 25109 22569 25143
rect 22569 25109 22603 25143
rect 22603 25109 22612 25143
rect 22560 25100 22612 25109
rect 7896 24998 7948 25050
rect 7960 24998 8012 25050
rect 8024 24998 8076 25050
rect 8088 24998 8140 25050
rect 8152 24998 8204 25050
rect 14842 24998 14894 25050
rect 14906 24998 14958 25050
rect 14970 24998 15022 25050
rect 15034 24998 15086 25050
rect 15098 24998 15150 25050
rect 21788 24998 21840 25050
rect 21852 24998 21904 25050
rect 21916 24998 21968 25050
rect 21980 24998 22032 25050
rect 22044 24998 22096 25050
rect 28734 24998 28786 25050
rect 28798 24998 28850 25050
rect 28862 24998 28914 25050
rect 28926 24998 28978 25050
rect 28990 24998 29042 25050
rect 19984 24896 20036 24948
rect 25228 24896 25280 24948
rect 26700 24896 26752 24948
rect 21088 24828 21140 24880
rect 21548 24828 21600 24880
rect 1584 24803 1636 24812
rect 1584 24769 1593 24803
rect 1593 24769 1627 24803
rect 1627 24769 1636 24803
rect 1584 24760 1636 24769
rect 16856 24760 16908 24812
rect 17500 24760 17552 24812
rect 20444 24760 20496 24812
rect 21640 24760 21692 24812
rect 22468 24760 22520 24812
rect 22836 24803 22888 24812
rect 22836 24769 22845 24803
rect 22845 24769 22879 24803
rect 22879 24769 22888 24803
rect 22836 24760 22888 24769
rect 24032 24760 24084 24812
rect 25596 24803 25648 24812
rect 25596 24769 25605 24803
rect 25605 24769 25639 24803
rect 25639 24769 25648 24803
rect 25596 24760 25648 24769
rect 26148 24828 26200 24880
rect 25872 24803 25924 24812
rect 25872 24769 25881 24803
rect 25881 24769 25915 24803
rect 25915 24769 25924 24803
rect 25872 24760 25924 24769
rect 26884 24760 26936 24812
rect 27068 24760 27120 24812
rect 27712 24760 27764 24812
rect 20168 24692 20220 24744
rect 21180 24735 21232 24744
rect 21180 24701 21189 24735
rect 21189 24701 21223 24735
rect 21223 24701 21232 24735
rect 21180 24692 21232 24701
rect 22744 24692 22796 24744
rect 24676 24692 24728 24744
rect 25780 24735 25832 24744
rect 25780 24701 25789 24735
rect 25789 24701 25823 24735
rect 25823 24701 25832 24735
rect 25780 24692 25832 24701
rect 18788 24667 18840 24676
rect 18788 24633 18797 24667
rect 18797 24633 18831 24667
rect 18831 24633 18840 24667
rect 18788 24624 18840 24633
rect 24124 24624 24176 24676
rect 15752 24556 15804 24608
rect 19892 24556 19944 24608
rect 24676 24599 24728 24608
rect 24676 24565 24685 24599
rect 24685 24565 24719 24599
rect 24719 24565 24728 24599
rect 24676 24556 24728 24565
rect 4423 24454 4475 24506
rect 4487 24454 4539 24506
rect 4551 24454 4603 24506
rect 4615 24454 4667 24506
rect 4679 24454 4731 24506
rect 11369 24454 11421 24506
rect 11433 24454 11485 24506
rect 11497 24454 11549 24506
rect 11561 24454 11613 24506
rect 11625 24454 11677 24506
rect 18315 24454 18367 24506
rect 18379 24454 18431 24506
rect 18443 24454 18495 24506
rect 18507 24454 18559 24506
rect 18571 24454 18623 24506
rect 25261 24454 25313 24506
rect 25325 24454 25377 24506
rect 25389 24454 25441 24506
rect 25453 24454 25505 24506
rect 25517 24454 25569 24506
rect 17500 24352 17552 24404
rect 21640 24395 21692 24404
rect 21640 24361 21649 24395
rect 21649 24361 21683 24395
rect 21683 24361 21692 24395
rect 21640 24352 21692 24361
rect 23756 24352 23808 24404
rect 24952 24352 25004 24404
rect 28356 24259 28408 24268
rect 28356 24225 28365 24259
rect 28365 24225 28399 24259
rect 28399 24225 28408 24259
rect 28356 24216 28408 24225
rect 17132 24191 17184 24200
rect 17132 24157 17141 24191
rect 17141 24157 17175 24191
rect 17175 24157 17184 24191
rect 17132 24148 17184 24157
rect 17316 24191 17368 24200
rect 17316 24157 17325 24191
rect 17325 24157 17359 24191
rect 17359 24157 17368 24191
rect 17316 24148 17368 24157
rect 19432 24191 19484 24200
rect 19432 24157 19441 24191
rect 19441 24157 19475 24191
rect 19475 24157 19484 24191
rect 19432 24148 19484 24157
rect 22376 24148 22428 24200
rect 23388 24148 23440 24200
rect 24676 24191 24728 24200
rect 24676 24157 24685 24191
rect 24685 24157 24719 24191
rect 24719 24157 24728 24191
rect 24676 24148 24728 24157
rect 24860 24191 24912 24200
rect 24860 24157 24869 24191
rect 24869 24157 24903 24191
rect 24903 24157 24912 24191
rect 24860 24148 24912 24157
rect 25688 24148 25740 24200
rect 26516 24191 26568 24200
rect 26516 24157 26525 24191
rect 26525 24157 26559 24191
rect 26559 24157 26568 24191
rect 26516 24148 26568 24157
rect 19708 24123 19760 24132
rect 19708 24089 19742 24123
rect 19742 24089 19760 24123
rect 23480 24123 23532 24132
rect 19708 24080 19760 24089
rect 23480 24089 23489 24123
rect 23489 24089 23523 24123
rect 23523 24089 23532 24123
rect 23480 24080 23532 24089
rect 23664 24123 23716 24132
rect 23664 24089 23689 24123
rect 23689 24089 23716 24123
rect 23664 24080 23716 24089
rect 27344 24080 27396 24132
rect 20996 24012 21048 24064
rect 24032 24012 24084 24064
rect 7896 23910 7948 23962
rect 7960 23910 8012 23962
rect 8024 23910 8076 23962
rect 8088 23910 8140 23962
rect 8152 23910 8204 23962
rect 14842 23910 14894 23962
rect 14906 23910 14958 23962
rect 14970 23910 15022 23962
rect 15034 23910 15086 23962
rect 15098 23910 15150 23962
rect 21788 23910 21840 23962
rect 21852 23910 21904 23962
rect 21916 23910 21968 23962
rect 21980 23910 22032 23962
rect 22044 23910 22096 23962
rect 28734 23910 28786 23962
rect 28798 23910 28850 23962
rect 28862 23910 28914 23962
rect 28926 23910 28978 23962
rect 28990 23910 29042 23962
rect 19708 23851 19760 23860
rect 19708 23817 19717 23851
rect 19717 23817 19751 23851
rect 19751 23817 19760 23851
rect 19708 23808 19760 23817
rect 20444 23851 20496 23860
rect 20444 23817 20453 23851
rect 20453 23817 20487 23851
rect 20487 23817 20496 23851
rect 20444 23808 20496 23817
rect 20904 23851 20956 23860
rect 20904 23817 20913 23851
rect 20913 23817 20947 23851
rect 20947 23817 20956 23851
rect 20904 23808 20956 23817
rect 27344 23851 27396 23860
rect 27344 23817 27353 23851
rect 27353 23817 27387 23851
rect 27387 23817 27396 23851
rect 27344 23808 27396 23817
rect 16580 23740 16632 23792
rect 18696 23672 18748 23724
rect 19800 23740 19852 23792
rect 20260 23740 20312 23792
rect 20996 23740 21048 23792
rect 26516 23740 26568 23792
rect 19892 23715 19944 23724
rect 19892 23681 19901 23715
rect 19901 23681 19935 23715
rect 19935 23681 19944 23715
rect 19892 23672 19944 23681
rect 26884 23672 26936 23724
rect 27620 23672 27672 23724
rect 21180 23604 21232 23656
rect 21640 23604 21692 23656
rect 17592 23536 17644 23588
rect 16396 23468 16448 23520
rect 17684 23468 17736 23520
rect 18880 23468 18932 23520
rect 26516 23468 26568 23520
rect 4423 23366 4475 23418
rect 4487 23366 4539 23418
rect 4551 23366 4603 23418
rect 4615 23366 4667 23418
rect 4679 23366 4731 23418
rect 11369 23366 11421 23418
rect 11433 23366 11485 23418
rect 11497 23366 11549 23418
rect 11561 23366 11613 23418
rect 11625 23366 11677 23418
rect 18315 23366 18367 23418
rect 18379 23366 18431 23418
rect 18443 23366 18495 23418
rect 18507 23366 18559 23418
rect 18571 23366 18623 23418
rect 25261 23366 25313 23418
rect 25325 23366 25377 23418
rect 25389 23366 25441 23418
rect 25453 23366 25505 23418
rect 25517 23366 25569 23418
rect 17316 23264 17368 23316
rect 23572 23196 23624 23248
rect 16396 23103 16448 23112
rect 16396 23069 16405 23103
rect 16405 23069 16439 23103
rect 16439 23069 16448 23103
rect 16396 23060 16448 23069
rect 17224 23128 17276 23180
rect 17684 23171 17736 23180
rect 17684 23137 17693 23171
rect 17693 23137 17727 23171
rect 17727 23137 17736 23171
rect 17684 23128 17736 23137
rect 19800 23171 19852 23180
rect 16580 23060 16632 23112
rect 17040 23060 17092 23112
rect 17592 23103 17644 23112
rect 17592 23069 17601 23103
rect 17601 23069 17635 23103
rect 17635 23069 17644 23103
rect 17592 23060 17644 23069
rect 17868 23103 17920 23112
rect 17868 23069 17877 23103
rect 17877 23069 17911 23103
rect 17911 23069 17920 23103
rect 17868 23060 17920 23069
rect 16212 22992 16264 23044
rect 17224 22992 17276 23044
rect 18696 23060 18748 23112
rect 19800 23137 19809 23171
rect 19809 23137 19843 23171
rect 19843 23137 19852 23171
rect 19800 23128 19852 23137
rect 20168 23128 20220 23180
rect 20536 23171 20588 23180
rect 20536 23137 20545 23171
rect 20545 23137 20579 23171
rect 20579 23137 20588 23171
rect 20536 23128 20588 23137
rect 25044 23128 25096 23180
rect 25780 23128 25832 23180
rect 26516 23171 26568 23180
rect 26516 23137 26525 23171
rect 26525 23137 26559 23171
rect 26559 23137 26568 23171
rect 26516 23128 26568 23137
rect 29920 23128 29972 23180
rect 20720 23103 20772 23112
rect 20720 23069 20729 23103
rect 20729 23069 20763 23103
rect 20763 23069 20772 23103
rect 20720 23060 20772 23069
rect 23664 23060 23716 23112
rect 24676 23060 24728 23112
rect 23756 23035 23808 23044
rect 23756 23001 23765 23035
rect 23765 23001 23799 23035
rect 23799 23001 23808 23035
rect 23756 22992 23808 23001
rect 26148 22992 26200 23044
rect 27252 22992 27304 23044
rect 15752 22967 15804 22976
rect 15752 22933 15761 22967
rect 15761 22933 15795 22967
rect 15795 22933 15804 22967
rect 15752 22924 15804 22933
rect 19984 22924 20036 22976
rect 20904 22967 20956 22976
rect 20904 22933 20913 22967
rect 20913 22933 20947 22967
rect 20947 22933 20956 22967
rect 20904 22924 20956 22933
rect 23480 22924 23532 22976
rect 24676 22924 24728 22976
rect 25596 22924 25648 22976
rect 7896 22822 7948 22874
rect 7960 22822 8012 22874
rect 8024 22822 8076 22874
rect 8088 22822 8140 22874
rect 8152 22822 8204 22874
rect 14842 22822 14894 22874
rect 14906 22822 14958 22874
rect 14970 22822 15022 22874
rect 15034 22822 15086 22874
rect 15098 22822 15150 22874
rect 21788 22822 21840 22874
rect 21852 22822 21904 22874
rect 21916 22822 21968 22874
rect 21980 22822 22032 22874
rect 22044 22822 22096 22874
rect 28734 22822 28786 22874
rect 28798 22822 28850 22874
rect 28862 22822 28914 22874
rect 28926 22822 28978 22874
rect 28990 22822 29042 22874
rect 17040 22720 17092 22772
rect 15752 22652 15804 22704
rect 17040 22627 17092 22636
rect 17040 22593 17049 22627
rect 17049 22593 17083 22627
rect 17083 22593 17092 22627
rect 17040 22584 17092 22593
rect 17224 22627 17276 22636
rect 17224 22593 17233 22627
rect 17233 22593 17267 22627
rect 17267 22593 17276 22627
rect 17224 22584 17276 22593
rect 17776 22584 17828 22636
rect 18236 22720 18288 22772
rect 20720 22763 20772 22772
rect 20720 22729 20729 22763
rect 20729 22729 20763 22763
rect 20763 22729 20772 22763
rect 20720 22720 20772 22729
rect 21180 22763 21232 22772
rect 21180 22729 21189 22763
rect 21189 22729 21223 22763
rect 21223 22729 21232 22763
rect 21180 22720 21232 22729
rect 26148 22720 26200 22772
rect 27252 22763 27304 22772
rect 27252 22729 27261 22763
rect 27261 22729 27295 22763
rect 27295 22729 27304 22763
rect 27252 22720 27304 22729
rect 21272 22652 21324 22704
rect 23388 22652 23440 22704
rect 18696 22627 18748 22636
rect 18696 22593 18705 22627
rect 18705 22593 18739 22627
rect 18739 22593 18748 22627
rect 18696 22584 18748 22593
rect 18880 22627 18932 22636
rect 18880 22593 18889 22627
rect 18889 22593 18923 22627
rect 18923 22593 18932 22627
rect 18880 22584 18932 22593
rect 18972 22627 19024 22636
rect 18972 22593 18980 22627
rect 18980 22593 19014 22627
rect 19014 22593 19024 22627
rect 18972 22584 19024 22593
rect 19800 22627 19852 22636
rect 17316 22559 17368 22568
rect 17316 22525 17325 22559
rect 17325 22525 17359 22559
rect 17359 22525 17368 22559
rect 19800 22593 19809 22627
rect 19809 22593 19843 22627
rect 19843 22593 19852 22627
rect 19800 22584 19852 22593
rect 22652 22584 22704 22636
rect 23756 22584 23808 22636
rect 23940 22584 23992 22636
rect 24032 22627 24084 22636
rect 24032 22593 24041 22627
rect 24041 22593 24075 22627
rect 24075 22593 24084 22627
rect 24308 22627 24360 22636
rect 24032 22584 24084 22593
rect 24308 22593 24317 22627
rect 24317 22593 24351 22627
rect 24351 22593 24360 22627
rect 24308 22584 24360 22593
rect 25228 22584 25280 22636
rect 28632 22584 28684 22636
rect 17316 22516 17368 22525
rect 21640 22516 21692 22568
rect 24124 22559 24176 22568
rect 24124 22525 24133 22559
rect 24133 22525 24167 22559
rect 24167 22525 24176 22559
rect 24124 22516 24176 22525
rect 19984 22448 20036 22500
rect 23572 22448 23624 22500
rect 16856 22423 16908 22432
rect 16856 22389 16865 22423
rect 16865 22389 16899 22423
rect 16899 22389 16908 22423
rect 16856 22380 16908 22389
rect 19064 22380 19116 22432
rect 22468 22380 22520 22432
rect 23848 22380 23900 22432
rect 28080 22423 28132 22432
rect 28080 22389 28089 22423
rect 28089 22389 28123 22423
rect 28123 22389 28132 22423
rect 28080 22380 28132 22389
rect 4423 22278 4475 22330
rect 4487 22278 4539 22330
rect 4551 22278 4603 22330
rect 4615 22278 4667 22330
rect 4679 22278 4731 22330
rect 11369 22278 11421 22330
rect 11433 22278 11485 22330
rect 11497 22278 11549 22330
rect 11561 22278 11613 22330
rect 11625 22278 11677 22330
rect 18315 22278 18367 22330
rect 18379 22278 18431 22330
rect 18443 22278 18495 22330
rect 18507 22278 18559 22330
rect 18571 22278 18623 22330
rect 25261 22278 25313 22330
rect 25325 22278 25377 22330
rect 25389 22278 25441 22330
rect 25453 22278 25505 22330
rect 25517 22278 25569 22330
rect 18696 22176 18748 22228
rect 23940 22176 23992 22228
rect 24400 22176 24452 22228
rect 25136 22176 25188 22228
rect 17132 22040 17184 22092
rect 27528 22083 27580 22092
rect 16856 21972 16908 22024
rect 18236 21972 18288 22024
rect 19432 21972 19484 22024
rect 21456 21972 21508 22024
rect 22468 22015 22520 22024
rect 22468 21981 22477 22015
rect 22477 21981 22511 22015
rect 22511 21981 22520 22015
rect 22468 21972 22520 21981
rect 22928 21972 22980 22024
rect 23848 22015 23900 22024
rect 23848 21981 23857 22015
rect 23857 21981 23891 22015
rect 23891 21981 23900 22015
rect 23848 21972 23900 21981
rect 19708 21904 19760 21956
rect 20720 21947 20772 21956
rect 20720 21913 20754 21947
rect 20754 21913 20772 21947
rect 20720 21904 20772 21913
rect 16120 21879 16172 21888
rect 16120 21845 16129 21879
rect 16129 21845 16163 21879
rect 16163 21845 16172 21879
rect 16120 21836 16172 21845
rect 21272 21836 21324 21888
rect 23112 21836 23164 21888
rect 24216 21972 24268 22024
rect 24676 21972 24728 22024
rect 27528 22049 27537 22083
rect 27537 22049 27571 22083
rect 27571 22049 27580 22083
rect 27528 22040 27580 22049
rect 28080 22040 28132 22092
rect 26148 21972 26200 22024
rect 27896 21904 27948 21956
rect 24860 21836 24912 21888
rect 7896 21734 7948 21786
rect 7960 21734 8012 21786
rect 8024 21734 8076 21786
rect 8088 21734 8140 21786
rect 8152 21734 8204 21786
rect 14842 21734 14894 21786
rect 14906 21734 14958 21786
rect 14970 21734 15022 21786
rect 15034 21734 15086 21786
rect 15098 21734 15150 21786
rect 21788 21734 21840 21786
rect 21852 21734 21904 21786
rect 21916 21734 21968 21786
rect 21980 21734 22032 21786
rect 22044 21734 22096 21786
rect 28734 21734 28786 21786
rect 28798 21734 28850 21786
rect 28862 21734 28914 21786
rect 28926 21734 28978 21786
rect 28990 21734 29042 21786
rect 16212 21632 16264 21684
rect 20720 21675 20772 21684
rect 20720 21641 20729 21675
rect 20729 21641 20763 21675
rect 20763 21641 20772 21675
rect 20720 21632 20772 21641
rect 22928 21675 22980 21684
rect 22928 21641 22937 21675
rect 22937 21641 22971 21675
rect 22971 21641 22980 21675
rect 22928 21632 22980 21641
rect 27896 21675 27948 21684
rect 27896 21641 27905 21675
rect 27905 21641 27939 21675
rect 27939 21641 27948 21675
rect 27896 21632 27948 21641
rect 16120 21564 16172 21616
rect 24400 21564 24452 21616
rect 19708 21496 19760 21548
rect 20904 21539 20956 21548
rect 20904 21505 20913 21539
rect 20913 21505 20947 21539
rect 20947 21505 20956 21539
rect 20904 21496 20956 21505
rect 22376 21496 22428 21548
rect 23664 21496 23716 21548
rect 24124 21496 24176 21548
rect 22008 21428 22060 21480
rect 22744 21471 22796 21480
rect 22744 21437 22753 21471
rect 22753 21437 22787 21471
rect 22787 21437 22796 21471
rect 22744 21428 22796 21437
rect 18236 21292 18288 21344
rect 24308 21428 24360 21480
rect 24860 21496 24912 21548
rect 25044 21496 25096 21548
rect 25596 21564 25648 21616
rect 25320 21496 25372 21548
rect 25688 21496 25740 21548
rect 27436 21496 27488 21548
rect 27804 21539 27856 21548
rect 27804 21505 27813 21539
rect 27813 21505 27847 21539
rect 27847 21505 27856 21539
rect 27804 21496 27856 21505
rect 28172 21496 28224 21548
rect 26976 21428 27028 21480
rect 25320 21360 25372 21412
rect 24032 21292 24084 21344
rect 25136 21292 25188 21344
rect 26700 21292 26752 21344
rect 4423 21190 4475 21242
rect 4487 21190 4539 21242
rect 4551 21190 4603 21242
rect 4615 21190 4667 21242
rect 4679 21190 4731 21242
rect 11369 21190 11421 21242
rect 11433 21190 11485 21242
rect 11497 21190 11549 21242
rect 11561 21190 11613 21242
rect 11625 21190 11677 21242
rect 18315 21190 18367 21242
rect 18379 21190 18431 21242
rect 18443 21190 18495 21242
rect 18507 21190 18559 21242
rect 18571 21190 18623 21242
rect 25261 21190 25313 21242
rect 25325 21190 25377 21242
rect 25389 21190 25441 21242
rect 25453 21190 25505 21242
rect 25517 21190 25569 21242
rect 16028 20927 16080 20936
rect 16028 20893 16037 20927
rect 16037 20893 16071 20927
rect 16071 20893 16080 20927
rect 16028 20884 16080 20893
rect 21640 20952 21692 21004
rect 23388 20995 23440 21004
rect 23388 20961 23397 20995
rect 23397 20961 23431 20995
rect 23431 20961 23440 20995
rect 23388 20952 23440 20961
rect 27712 20952 27764 21004
rect 28356 20995 28408 21004
rect 28356 20961 28365 20995
rect 28365 20961 28399 20995
rect 28399 20961 28408 20995
rect 28356 20952 28408 20961
rect 19340 20816 19392 20868
rect 20536 20884 20588 20936
rect 23112 20927 23164 20936
rect 23112 20893 23130 20927
rect 23130 20893 23164 20927
rect 23112 20884 23164 20893
rect 27344 20816 27396 20868
rect 16948 20748 17000 20800
rect 19524 20748 19576 20800
rect 20352 20748 20404 20800
rect 22008 20791 22060 20800
rect 22008 20757 22017 20791
rect 22017 20757 22051 20791
rect 22051 20757 22060 20791
rect 22008 20748 22060 20757
rect 7896 20646 7948 20698
rect 7960 20646 8012 20698
rect 8024 20646 8076 20698
rect 8088 20646 8140 20698
rect 8152 20646 8204 20698
rect 14842 20646 14894 20698
rect 14906 20646 14958 20698
rect 14970 20646 15022 20698
rect 15034 20646 15086 20698
rect 15098 20646 15150 20698
rect 21788 20646 21840 20698
rect 21852 20646 21904 20698
rect 21916 20646 21968 20698
rect 21980 20646 22032 20698
rect 22044 20646 22096 20698
rect 28734 20646 28786 20698
rect 28798 20646 28850 20698
rect 28862 20646 28914 20698
rect 28926 20646 28978 20698
rect 28990 20646 29042 20698
rect 16028 20544 16080 20596
rect 25688 20544 25740 20596
rect 2044 20408 2096 20460
rect 15200 20408 15252 20460
rect 15660 20451 15712 20460
rect 15660 20417 15669 20451
rect 15669 20417 15703 20451
rect 15703 20417 15712 20451
rect 15660 20408 15712 20417
rect 15844 20408 15896 20460
rect 18236 20476 18288 20528
rect 19524 20519 19576 20528
rect 19524 20485 19558 20519
rect 19558 20485 19576 20519
rect 19524 20476 19576 20485
rect 25596 20476 25648 20528
rect 16948 20408 17000 20460
rect 23480 20340 23532 20392
rect 1768 20204 1820 20256
rect 15292 20204 15344 20256
rect 20352 20204 20404 20256
rect 27896 20247 27948 20256
rect 27896 20213 27905 20247
rect 27905 20213 27939 20247
rect 27939 20213 27948 20247
rect 27896 20204 27948 20213
rect 4423 20102 4475 20154
rect 4487 20102 4539 20154
rect 4551 20102 4603 20154
rect 4615 20102 4667 20154
rect 4679 20102 4731 20154
rect 11369 20102 11421 20154
rect 11433 20102 11485 20154
rect 11497 20102 11549 20154
rect 11561 20102 11613 20154
rect 11625 20102 11677 20154
rect 18315 20102 18367 20154
rect 18379 20102 18431 20154
rect 18443 20102 18495 20154
rect 18507 20102 18559 20154
rect 18571 20102 18623 20154
rect 25261 20102 25313 20154
rect 25325 20102 25377 20154
rect 25389 20102 25441 20154
rect 25453 20102 25505 20154
rect 25517 20102 25569 20154
rect 15200 20043 15252 20052
rect 15200 20009 15209 20043
rect 15209 20009 15243 20043
rect 15243 20009 15252 20043
rect 15200 20000 15252 20009
rect 1768 19907 1820 19916
rect 1768 19873 1777 19907
rect 1777 19873 1811 19907
rect 1811 19873 1820 19907
rect 1768 19864 1820 19873
rect 2780 19907 2832 19916
rect 2780 19873 2789 19907
rect 2789 19873 2823 19907
rect 2823 19873 2832 19907
rect 2780 19864 2832 19873
rect 15476 19864 15528 19916
rect 1584 19839 1636 19848
rect 1584 19805 1593 19839
rect 1593 19805 1627 19839
rect 1627 19805 1636 19839
rect 1584 19796 1636 19805
rect 15292 19796 15344 19848
rect 21456 19839 21508 19848
rect 21456 19805 21465 19839
rect 21465 19805 21499 19839
rect 21499 19805 21508 19839
rect 21456 19796 21508 19805
rect 24676 19932 24728 19984
rect 24492 19864 24544 19916
rect 27896 19864 27948 19916
rect 28356 19907 28408 19916
rect 28356 19873 28365 19907
rect 28365 19873 28399 19907
rect 28399 19873 28408 19907
rect 28356 19864 28408 19873
rect 14372 19728 14424 19780
rect 21180 19728 21232 19780
rect 21824 19839 21876 19848
rect 21824 19805 21833 19839
rect 21833 19805 21867 19839
rect 21867 19805 21876 19839
rect 21824 19796 21876 19805
rect 22468 19796 22520 19848
rect 24768 19839 24820 19848
rect 24768 19805 24777 19839
rect 24777 19805 24811 19839
rect 24811 19805 24820 19839
rect 24768 19796 24820 19805
rect 25044 19839 25096 19848
rect 25044 19805 25053 19839
rect 25053 19805 25087 19839
rect 25087 19805 25096 19839
rect 25044 19796 25096 19805
rect 25228 19839 25280 19848
rect 25228 19805 25237 19839
rect 25237 19805 25271 19839
rect 25271 19805 25280 19839
rect 25228 19796 25280 19805
rect 22376 19728 22428 19780
rect 26700 19771 26752 19780
rect 26700 19737 26709 19771
rect 26709 19737 26743 19771
rect 26743 19737 26752 19771
rect 26700 19728 26752 19737
rect 15660 19703 15712 19712
rect 15660 19669 15669 19703
rect 15669 19669 15703 19703
rect 15703 19669 15712 19703
rect 15660 19660 15712 19669
rect 23204 19660 23256 19712
rect 24860 19660 24912 19712
rect 7896 19558 7948 19610
rect 7960 19558 8012 19610
rect 8024 19558 8076 19610
rect 8088 19558 8140 19610
rect 8152 19558 8204 19610
rect 14842 19558 14894 19610
rect 14906 19558 14958 19610
rect 14970 19558 15022 19610
rect 15034 19558 15086 19610
rect 15098 19558 15150 19610
rect 21788 19558 21840 19610
rect 21852 19558 21904 19610
rect 21916 19558 21968 19610
rect 21980 19558 22032 19610
rect 22044 19558 22096 19610
rect 28734 19558 28786 19610
rect 28798 19558 28850 19610
rect 28862 19558 28914 19610
rect 28926 19558 28978 19610
rect 28990 19558 29042 19610
rect 16672 19456 16724 19508
rect 22468 19456 22520 19508
rect 25596 19499 25648 19508
rect 25596 19465 25605 19499
rect 25605 19465 25639 19499
rect 25639 19465 25648 19499
rect 25596 19456 25648 19465
rect 27344 19499 27396 19508
rect 27344 19465 27353 19499
rect 27353 19465 27387 19499
rect 27387 19465 27396 19499
rect 27344 19456 27396 19465
rect 17224 19388 17276 19440
rect 18880 19388 18932 19440
rect 1584 19320 1636 19372
rect 16120 19363 16172 19372
rect 16120 19329 16129 19363
rect 16129 19329 16163 19363
rect 16163 19329 16172 19363
rect 16120 19320 16172 19329
rect 16856 19363 16908 19372
rect 16856 19329 16865 19363
rect 16865 19329 16899 19363
rect 16899 19329 16908 19363
rect 16856 19320 16908 19329
rect 17408 19320 17460 19372
rect 18972 19363 19024 19372
rect 18972 19329 18981 19363
rect 18981 19329 19015 19363
rect 19015 19329 19024 19363
rect 18972 19320 19024 19329
rect 19708 19363 19760 19372
rect 18696 19184 18748 19236
rect 18788 19184 18840 19236
rect 19156 19295 19208 19304
rect 19156 19261 19165 19295
rect 19165 19261 19199 19295
rect 19199 19261 19208 19295
rect 19708 19329 19717 19363
rect 19717 19329 19751 19363
rect 19751 19329 19760 19363
rect 19708 19320 19760 19329
rect 20720 19320 20772 19372
rect 22284 19388 22336 19440
rect 23204 19431 23256 19440
rect 23204 19397 23222 19431
rect 23222 19397 23256 19431
rect 23204 19388 23256 19397
rect 25044 19388 25096 19440
rect 21180 19320 21232 19372
rect 22100 19320 22152 19372
rect 23480 19363 23532 19372
rect 23480 19329 23489 19363
rect 23489 19329 23523 19363
rect 23523 19329 23532 19363
rect 23480 19320 23532 19329
rect 24676 19320 24728 19372
rect 25136 19363 25188 19372
rect 25136 19329 25145 19363
rect 25145 19329 25179 19363
rect 25179 19329 25188 19363
rect 25136 19320 25188 19329
rect 25688 19320 25740 19372
rect 27252 19320 27304 19372
rect 27804 19320 27856 19372
rect 19156 19252 19208 19261
rect 19616 19252 19668 19304
rect 19800 19252 19852 19304
rect 20076 19295 20128 19304
rect 20076 19261 20085 19295
rect 20085 19261 20119 19295
rect 20119 19261 20128 19295
rect 20076 19252 20128 19261
rect 27712 19252 27764 19304
rect 18144 19116 18196 19168
rect 19156 19116 19208 19168
rect 19248 19116 19300 19168
rect 19984 19116 20036 19168
rect 4423 19014 4475 19066
rect 4487 19014 4539 19066
rect 4551 19014 4603 19066
rect 4615 19014 4667 19066
rect 4679 19014 4731 19066
rect 11369 19014 11421 19066
rect 11433 19014 11485 19066
rect 11497 19014 11549 19066
rect 11561 19014 11613 19066
rect 11625 19014 11677 19066
rect 18315 19014 18367 19066
rect 18379 19014 18431 19066
rect 18443 19014 18495 19066
rect 18507 19014 18559 19066
rect 18571 19014 18623 19066
rect 25261 19014 25313 19066
rect 25325 19014 25377 19066
rect 25389 19014 25441 19066
rect 25453 19014 25505 19066
rect 25517 19014 25569 19066
rect 1584 18751 1636 18760
rect 1584 18717 1593 18751
rect 1593 18717 1627 18751
rect 1627 18717 1636 18751
rect 1584 18708 1636 18717
rect 18052 18912 18104 18964
rect 18788 18912 18840 18964
rect 19248 18912 19300 18964
rect 19708 18912 19760 18964
rect 27528 18912 27580 18964
rect 17960 18776 18012 18828
rect 17224 18708 17276 18760
rect 17684 18708 17736 18760
rect 18052 18751 18104 18760
rect 18052 18717 18061 18751
rect 18061 18717 18095 18751
rect 18095 18717 18104 18751
rect 18052 18708 18104 18717
rect 23296 18844 23348 18896
rect 19340 18776 19392 18828
rect 19800 18776 19852 18828
rect 22100 18819 22152 18828
rect 22100 18785 22109 18819
rect 22109 18785 22143 18819
rect 22143 18785 22152 18819
rect 22100 18776 22152 18785
rect 22284 18819 22336 18828
rect 22284 18785 22293 18819
rect 22293 18785 22327 18819
rect 22327 18785 22336 18819
rect 22284 18776 22336 18785
rect 23204 18776 23256 18828
rect 24584 18776 24636 18828
rect 18972 18708 19024 18760
rect 19616 18751 19668 18760
rect 19616 18717 19625 18751
rect 19625 18717 19659 18751
rect 19659 18717 19668 18751
rect 19616 18708 19668 18717
rect 3332 18640 3384 18692
rect 20720 18640 20772 18692
rect 24952 18708 25004 18760
rect 28356 18751 28408 18760
rect 28356 18717 28365 18751
rect 28365 18717 28399 18751
rect 28399 18717 28408 18751
rect 28356 18708 28408 18717
rect 22376 18640 22428 18692
rect 23388 18640 23440 18692
rect 27988 18640 28040 18692
rect 15660 18572 15712 18624
rect 17224 18572 17276 18624
rect 17500 18572 17552 18624
rect 18512 18615 18564 18624
rect 18512 18581 18521 18615
rect 18521 18581 18555 18615
rect 18555 18581 18564 18615
rect 18512 18572 18564 18581
rect 23664 18572 23716 18624
rect 7896 18470 7948 18522
rect 7960 18470 8012 18522
rect 8024 18470 8076 18522
rect 8088 18470 8140 18522
rect 8152 18470 8204 18522
rect 14842 18470 14894 18522
rect 14906 18470 14958 18522
rect 14970 18470 15022 18522
rect 15034 18470 15086 18522
rect 15098 18470 15150 18522
rect 21788 18470 21840 18522
rect 21852 18470 21904 18522
rect 21916 18470 21968 18522
rect 21980 18470 22032 18522
rect 22044 18470 22096 18522
rect 28734 18470 28786 18522
rect 28798 18470 28850 18522
rect 28862 18470 28914 18522
rect 28926 18470 28978 18522
rect 28990 18470 29042 18522
rect 16856 18411 16908 18420
rect 16856 18377 16865 18411
rect 16865 18377 16899 18411
rect 16899 18377 16908 18411
rect 16856 18368 16908 18377
rect 17224 18411 17276 18420
rect 17224 18377 17233 18411
rect 17233 18377 17267 18411
rect 17267 18377 17276 18411
rect 17224 18368 17276 18377
rect 21456 18368 21508 18420
rect 23480 18368 23532 18420
rect 24584 18368 24636 18420
rect 27988 18411 28040 18420
rect 27988 18377 27997 18411
rect 27997 18377 28031 18411
rect 28031 18377 28040 18411
rect 27988 18368 28040 18377
rect 18512 18300 18564 18352
rect 22560 18300 22612 18352
rect 15660 18275 15712 18284
rect 15660 18241 15669 18275
rect 15669 18241 15703 18275
rect 15703 18241 15712 18275
rect 15660 18232 15712 18241
rect 15844 18275 15896 18284
rect 15844 18241 15853 18275
rect 15853 18241 15887 18275
rect 15887 18241 15896 18275
rect 17132 18275 17184 18284
rect 15844 18232 15896 18241
rect 17132 18241 17141 18275
rect 17141 18241 17175 18275
rect 17175 18241 17184 18275
rect 17132 18232 17184 18241
rect 17316 18275 17368 18284
rect 17316 18241 17325 18275
rect 17325 18241 17359 18275
rect 17359 18241 17368 18275
rect 17316 18232 17368 18241
rect 17500 18275 17552 18284
rect 17500 18241 17509 18275
rect 17509 18241 17543 18275
rect 17543 18241 17552 18275
rect 17500 18232 17552 18241
rect 20720 18232 20772 18284
rect 16212 18164 16264 18216
rect 18236 18207 18288 18216
rect 18236 18173 18245 18207
rect 18245 18173 18279 18207
rect 18279 18173 18288 18207
rect 18236 18164 18288 18173
rect 22192 18232 22244 18284
rect 23848 18232 23900 18284
rect 27344 18275 27396 18284
rect 27344 18241 27353 18275
rect 27353 18241 27387 18275
rect 27387 18241 27396 18275
rect 27344 18232 27396 18241
rect 22284 18164 22336 18216
rect 26516 18164 26568 18216
rect 23940 18096 23992 18148
rect 1584 18028 1636 18080
rect 16856 18028 16908 18080
rect 23664 18028 23716 18080
rect 4423 17926 4475 17978
rect 4487 17926 4539 17978
rect 4551 17926 4603 17978
rect 4615 17926 4667 17978
rect 4679 17926 4731 17978
rect 11369 17926 11421 17978
rect 11433 17926 11485 17978
rect 11497 17926 11549 17978
rect 11561 17926 11613 17978
rect 11625 17926 11677 17978
rect 18315 17926 18367 17978
rect 18379 17926 18431 17978
rect 18443 17926 18495 17978
rect 18507 17926 18559 17978
rect 18571 17926 18623 17978
rect 25261 17926 25313 17978
rect 25325 17926 25377 17978
rect 25389 17926 25441 17978
rect 25453 17926 25505 17978
rect 25517 17926 25569 17978
rect 2228 17824 2280 17876
rect 5172 17824 5224 17876
rect 15660 17824 15712 17876
rect 17132 17824 17184 17876
rect 17408 17867 17460 17876
rect 17408 17833 17417 17867
rect 17417 17833 17451 17867
rect 17451 17833 17460 17867
rect 17408 17824 17460 17833
rect 1860 17756 1912 17808
rect 1584 17731 1636 17740
rect 1584 17697 1593 17731
rect 1593 17697 1627 17731
rect 1627 17697 1636 17731
rect 1584 17688 1636 17697
rect 2780 17731 2832 17740
rect 2780 17697 2789 17731
rect 2789 17697 2823 17731
rect 2823 17697 2832 17731
rect 2780 17688 2832 17697
rect 15936 17731 15988 17740
rect 15936 17697 15945 17731
rect 15945 17697 15979 17731
rect 15979 17697 15988 17731
rect 15936 17688 15988 17697
rect 17224 17688 17276 17740
rect 19616 17824 19668 17876
rect 24584 17731 24636 17740
rect 18696 17620 18748 17672
rect 24584 17697 24593 17731
rect 24593 17697 24627 17731
rect 24627 17697 24636 17731
rect 24584 17688 24636 17697
rect 26148 17688 26200 17740
rect 28356 17731 28408 17740
rect 28356 17697 28365 17731
rect 28365 17697 28399 17731
rect 28399 17697 28408 17731
rect 28356 17688 28408 17697
rect 1952 17552 2004 17604
rect 17316 17552 17368 17604
rect 19892 17620 19944 17672
rect 23204 17620 23256 17672
rect 23388 17620 23440 17672
rect 24860 17663 24912 17672
rect 24860 17629 24894 17663
rect 24894 17629 24912 17663
rect 24860 17620 24912 17629
rect 17960 17484 18012 17536
rect 21456 17552 21508 17604
rect 28172 17595 28224 17604
rect 28172 17561 28181 17595
rect 28181 17561 28215 17595
rect 28215 17561 28224 17595
rect 28172 17552 28224 17561
rect 18420 17527 18472 17536
rect 18420 17493 18429 17527
rect 18429 17493 18463 17527
rect 18463 17493 18472 17527
rect 18420 17484 18472 17493
rect 22284 17484 22336 17536
rect 24124 17484 24176 17536
rect 25044 17484 25096 17536
rect 7896 17382 7948 17434
rect 7960 17382 8012 17434
rect 8024 17382 8076 17434
rect 8088 17382 8140 17434
rect 8152 17382 8204 17434
rect 14842 17382 14894 17434
rect 14906 17382 14958 17434
rect 14970 17382 15022 17434
rect 15034 17382 15086 17434
rect 15098 17382 15150 17434
rect 21788 17382 21840 17434
rect 21852 17382 21904 17434
rect 21916 17382 21968 17434
rect 21980 17382 22032 17434
rect 22044 17382 22096 17434
rect 28734 17382 28786 17434
rect 28798 17382 28850 17434
rect 28862 17382 28914 17434
rect 28926 17382 28978 17434
rect 28990 17382 29042 17434
rect 1952 17323 2004 17332
rect 1952 17289 1961 17323
rect 1961 17289 1995 17323
rect 1995 17289 2004 17323
rect 1952 17280 2004 17289
rect 18420 17280 18472 17332
rect 19892 17323 19944 17332
rect 19892 17289 19901 17323
rect 19901 17289 19935 17323
rect 19935 17289 19944 17323
rect 19892 17280 19944 17289
rect 15476 17212 15528 17264
rect 17316 17212 17368 17264
rect 2044 17187 2096 17196
rect 2044 17153 2053 17187
rect 2053 17153 2087 17187
rect 2087 17153 2096 17187
rect 2044 17144 2096 17153
rect 15844 17144 15896 17196
rect 16856 17187 16908 17196
rect 16856 17153 16865 17187
rect 16865 17153 16899 17187
rect 16899 17153 16908 17187
rect 16856 17144 16908 17153
rect 17868 17144 17920 17196
rect 19064 17212 19116 17264
rect 24676 17280 24728 17332
rect 27344 17280 27396 17332
rect 27528 17323 27580 17332
rect 27528 17289 27537 17323
rect 27537 17289 27571 17323
rect 27571 17289 27580 17323
rect 27528 17280 27580 17289
rect 18788 17144 18840 17196
rect 19616 17144 19668 17196
rect 23940 17212 23992 17264
rect 22192 17187 22244 17196
rect 22192 17153 22201 17187
rect 22201 17153 22235 17187
rect 22235 17153 22244 17187
rect 22192 17144 22244 17153
rect 23480 17144 23532 17196
rect 23664 17144 23716 17196
rect 26424 17187 26476 17196
rect 26424 17153 26433 17187
rect 26433 17153 26467 17187
rect 26467 17153 26476 17187
rect 26424 17144 26476 17153
rect 18696 17008 18748 17060
rect 19340 17076 19392 17128
rect 27620 17119 27672 17128
rect 27620 17085 27629 17119
rect 27629 17085 27663 17119
rect 27663 17085 27672 17119
rect 27620 17076 27672 17085
rect 25872 17008 25924 17060
rect 17132 16940 17184 16992
rect 17316 16940 17368 16992
rect 17868 16940 17920 16992
rect 23020 16983 23072 16992
rect 23020 16949 23029 16983
rect 23029 16949 23063 16983
rect 23063 16949 23072 16983
rect 23020 16940 23072 16949
rect 24952 16983 25004 16992
rect 24952 16949 24961 16983
rect 24961 16949 24995 16983
rect 24995 16949 25004 16983
rect 24952 16940 25004 16949
rect 26516 16983 26568 16992
rect 26516 16949 26525 16983
rect 26525 16949 26559 16983
rect 26559 16949 26568 16983
rect 26516 16940 26568 16949
rect 4423 16838 4475 16890
rect 4487 16838 4539 16890
rect 4551 16838 4603 16890
rect 4615 16838 4667 16890
rect 4679 16838 4731 16890
rect 11369 16838 11421 16890
rect 11433 16838 11485 16890
rect 11497 16838 11549 16890
rect 11561 16838 11613 16890
rect 11625 16838 11677 16890
rect 18315 16838 18367 16890
rect 18379 16838 18431 16890
rect 18443 16838 18495 16890
rect 18507 16838 18559 16890
rect 18571 16838 18623 16890
rect 25261 16838 25313 16890
rect 25325 16838 25377 16890
rect 25389 16838 25441 16890
rect 25453 16838 25505 16890
rect 25517 16838 25569 16890
rect 13268 16779 13320 16788
rect 13268 16745 13277 16779
rect 13277 16745 13311 16779
rect 13311 16745 13320 16779
rect 13268 16736 13320 16745
rect 2228 16600 2280 16652
rect 18236 16736 18288 16788
rect 18788 16779 18840 16788
rect 18788 16745 18797 16779
rect 18797 16745 18831 16779
rect 18831 16745 18840 16779
rect 18788 16736 18840 16745
rect 17868 16668 17920 16720
rect 25872 16736 25924 16788
rect 26424 16736 26476 16788
rect 28172 16736 28224 16788
rect 13452 16575 13504 16584
rect 13452 16541 13461 16575
rect 13461 16541 13495 16575
rect 13495 16541 13504 16575
rect 13452 16532 13504 16541
rect 13728 16575 13780 16584
rect 13728 16541 13737 16575
rect 13737 16541 13771 16575
rect 13771 16541 13780 16575
rect 13728 16532 13780 16541
rect 17132 16575 17184 16584
rect 17132 16541 17166 16575
rect 17166 16541 17184 16575
rect 17132 16532 17184 16541
rect 20444 16600 20496 16652
rect 21272 16643 21324 16652
rect 21272 16609 21281 16643
rect 21281 16609 21315 16643
rect 21315 16609 21324 16643
rect 21272 16600 21324 16609
rect 23480 16600 23532 16652
rect 18972 16532 19024 16584
rect 16028 16464 16080 16516
rect 20812 16532 20864 16584
rect 23020 16575 23072 16584
rect 23020 16541 23038 16575
rect 23038 16541 23072 16575
rect 23756 16575 23808 16584
rect 23020 16532 23072 16541
rect 23756 16541 23765 16575
rect 23765 16541 23799 16575
rect 23799 16541 23808 16575
rect 23756 16532 23808 16541
rect 24032 16600 24084 16652
rect 26516 16600 26568 16652
rect 23848 16507 23900 16516
rect 1860 16396 1912 16448
rect 13820 16396 13872 16448
rect 17960 16396 18012 16448
rect 19432 16396 19484 16448
rect 22376 16396 22428 16448
rect 23848 16473 23857 16507
rect 23857 16473 23891 16507
rect 23891 16473 23900 16507
rect 23848 16464 23900 16473
rect 25596 16575 25648 16584
rect 25596 16541 25605 16575
rect 25605 16541 25639 16575
rect 25639 16541 25648 16575
rect 25596 16532 25648 16541
rect 27344 16575 27396 16584
rect 27344 16541 27353 16575
rect 27353 16541 27387 16575
rect 27387 16541 27396 16575
rect 27344 16532 27396 16541
rect 27896 16600 27948 16652
rect 24676 16439 24728 16448
rect 24676 16405 24685 16439
rect 24685 16405 24719 16439
rect 24719 16405 24728 16439
rect 24676 16396 24728 16405
rect 24860 16396 24912 16448
rect 7896 16294 7948 16346
rect 7960 16294 8012 16346
rect 8024 16294 8076 16346
rect 8088 16294 8140 16346
rect 8152 16294 8204 16346
rect 14842 16294 14894 16346
rect 14906 16294 14958 16346
rect 14970 16294 15022 16346
rect 15034 16294 15086 16346
rect 15098 16294 15150 16346
rect 21788 16294 21840 16346
rect 21852 16294 21904 16346
rect 21916 16294 21968 16346
rect 21980 16294 22032 16346
rect 22044 16294 22096 16346
rect 28734 16294 28786 16346
rect 28798 16294 28850 16346
rect 28862 16294 28914 16346
rect 28926 16294 28978 16346
rect 28990 16294 29042 16346
rect 13728 16192 13780 16244
rect 20352 16235 20404 16244
rect 20352 16201 20361 16235
rect 20361 16201 20395 16235
rect 20395 16201 20404 16235
rect 20352 16192 20404 16201
rect 22192 16192 22244 16244
rect 22376 16235 22428 16244
rect 22376 16201 22385 16235
rect 22385 16201 22419 16235
rect 22419 16201 22428 16235
rect 22376 16192 22428 16201
rect 1860 16167 1912 16176
rect 1860 16133 1869 16167
rect 1869 16133 1903 16167
rect 1903 16133 1912 16167
rect 1860 16124 1912 16133
rect 16028 16124 16080 16176
rect 24492 16124 24544 16176
rect 1676 16031 1728 16040
rect 1676 15997 1685 16031
rect 1685 15997 1719 16031
rect 1719 15997 1728 16031
rect 1676 15988 1728 15997
rect 2780 16031 2832 16040
rect 2780 15997 2789 16031
rect 2789 15997 2823 16031
rect 2823 15997 2832 16031
rect 2780 15988 2832 15997
rect 14280 16056 14332 16108
rect 15200 16056 15252 16108
rect 15844 16056 15896 16108
rect 20812 16056 20864 16108
rect 24860 16056 24912 16108
rect 27160 16056 27212 16108
rect 20720 15988 20772 16040
rect 22560 16031 22612 16040
rect 22560 15997 22569 16031
rect 22569 15997 22603 16031
rect 22603 15997 22612 16031
rect 22560 15988 22612 15997
rect 23480 15988 23532 16040
rect 23848 15988 23900 16040
rect 22836 15920 22888 15972
rect 14648 15852 14700 15904
rect 16304 15852 16356 15904
rect 26608 15895 26660 15904
rect 26608 15861 26617 15895
rect 26617 15861 26651 15895
rect 26651 15861 26660 15895
rect 26608 15852 26660 15861
rect 28172 15852 28224 15904
rect 28356 15852 28408 15904
rect 4423 15750 4475 15802
rect 4487 15750 4539 15802
rect 4551 15750 4603 15802
rect 4615 15750 4667 15802
rect 4679 15750 4731 15802
rect 11369 15750 11421 15802
rect 11433 15750 11485 15802
rect 11497 15750 11549 15802
rect 11561 15750 11613 15802
rect 11625 15750 11677 15802
rect 18315 15750 18367 15802
rect 18379 15750 18431 15802
rect 18443 15750 18495 15802
rect 18507 15750 18559 15802
rect 18571 15750 18623 15802
rect 25261 15750 25313 15802
rect 25325 15750 25377 15802
rect 25389 15750 25441 15802
rect 25453 15750 25505 15802
rect 25517 15750 25569 15802
rect 1676 15691 1728 15700
rect 1676 15657 1685 15691
rect 1685 15657 1719 15691
rect 1719 15657 1728 15691
rect 1676 15648 1728 15657
rect 13820 15648 13872 15700
rect 15752 15691 15804 15700
rect 15752 15657 15761 15691
rect 15761 15657 15795 15691
rect 15795 15657 15804 15691
rect 15752 15648 15804 15657
rect 20444 15648 20496 15700
rect 19616 15580 19668 15632
rect 12900 15444 12952 15496
rect 13728 15487 13780 15496
rect 13728 15453 13737 15487
rect 13737 15453 13771 15487
rect 13771 15453 13780 15487
rect 13728 15444 13780 15453
rect 14372 15444 14424 15496
rect 14648 15487 14700 15496
rect 14648 15453 14657 15487
rect 14657 15453 14691 15487
rect 14691 15453 14700 15487
rect 14648 15444 14700 15453
rect 15292 15444 15344 15496
rect 20996 15512 21048 15564
rect 20720 15487 20772 15496
rect 20720 15453 20729 15487
rect 20729 15453 20763 15487
rect 20763 15453 20772 15487
rect 20720 15444 20772 15453
rect 21548 15444 21600 15496
rect 25596 15648 25648 15700
rect 25872 15555 25924 15564
rect 25872 15521 25881 15555
rect 25881 15521 25915 15555
rect 25915 15521 25924 15555
rect 25872 15512 25924 15521
rect 27528 15555 27580 15564
rect 27528 15521 27537 15555
rect 27537 15521 27571 15555
rect 27571 15521 27580 15555
rect 27528 15512 27580 15521
rect 28172 15555 28224 15564
rect 28172 15521 28181 15555
rect 28181 15521 28215 15555
rect 28215 15521 28224 15555
rect 28172 15512 28224 15521
rect 28356 15555 28408 15564
rect 28356 15521 28365 15555
rect 28365 15521 28399 15555
rect 28399 15521 28408 15555
rect 28356 15512 28408 15521
rect 26608 15444 26660 15496
rect 15476 15308 15528 15360
rect 16120 15308 16172 15360
rect 20536 15308 20588 15360
rect 22652 15308 22704 15360
rect 25872 15308 25924 15360
rect 7896 15206 7948 15258
rect 7960 15206 8012 15258
rect 8024 15206 8076 15258
rect 8088 15206 8140 15258
rect 8152 15206 8204 15258
rect 14842 15206 14894 15258
rect 14906 15206 14958 15258
rect 14970 15206 15022 15258
rect 15034 15206 15086 15258
rect 15098 15206 15150 15258
rect 21788 15206 21840 15258
rect 21852 15206 21904 15258
rect 21916 15206 21968 15258
rect 21980 15206 22032 15258
rect 22044 15206 22096 15258
rect 28734 15206 28786 15258
rect 28798 15206 28850 15258
rect 28862 15206 28914 15258
rect 28926 15206 28978 15258
rect 28990 15206 29042 15258
rect 13452 15104 13504 15156
rect 14372 15147 14424 15156
rect 14372 15113 14381 15147
rect 14381 15113 14415 15147
rect 14415 15113 14424 15147
rect 14372 15104 14424 15113
rect 15752 15104 15804 15156
rect 16304 15147 16356 15156
rect 16304 15113 16313 15147
rect 16313 15113 16347 15147
rect 16347 15113 16356 15147
rect 16304 15104 16356 15113
rect 13728 15036 13780 15088
rect 2044 15011 2096 15020
rect 2044 14977 2053 15011
rect 2053 14977 2087 15011
rect 2087 14977 2096 15011
rect 2044 14968 2096 14977
rect 2504 14968 2556 15020
rect 13360 14968 13412 15020
rect 12900 14900 12952 14952
rect 14280 14968 14332 15020
rect 19616 15036 19668 15088
rect 19340 15011 19392 15020
rect 19340 14977 19374 15011
rect 19374 14977 19392 15011
rect 12624 14832 12676 14884
rect 14648 14832 14700 14884
rect 19340 14968 19392 14977
rect 23112 14968 23164 15020
rect 23848 15011 23900 15020
rect 23848 14977 23857 15011
rect 23857 14977 23891 15011
rect 23891 14977 23900 15011
rect 23848 14968 23900 14977
rect 26884 14968 26936 15020
rect 27528 14968 27580 15020
rect 15200 14875 15252 14884
rect 1768 14764 1820 14816
rect 14740 14764 14792 14816
rect 15200 14841 15209 14875
rect 15209 14841 15243 14875
rect 15243 14841 15252 14875
rect 15200 14832 15252 14841
rect 16120 14900 16172 14952
rect 19064 14943 19116 14952
rect 19064 14909 19073 14943
rect 19073 14909 19107 14943
rect 19107 14909 19116 14943
rect 19064 14900 19116 14909
rect 16028 14832 16080 14884
rect 15292 14764 15344 14816
rect 15568 14764 15620 14816
rect 20444 14807 20496 14816
rect 20444 14773 20453 14807
rect 20453 14773 20487 14807
rect 20487 14773 20496 14807
rect 20444 14764 20496 14773
rect 22376 14764 22428 14816
rect 26700 14764 26752 14816
rect 27896 14807 27948 14816
rect 27896 14773 27905 14807
rect 27905 14773 27939 14807
rect 27939 14773 27948 14807
rect 27896 14764 27948 14773
rect 4423 14662 4475 14714
rect 4487 14662 4539 14714
rect 4551 14662 4603 14714
rect 4615 14662 4667 14714
rect 4679 14662 4731 14714
rect 11369 14662 11421 14714
rect 11433 14662 11485 14714
rect 11497 14662 11549 14714
rect 11561 14662 11613 14714
rect 11625 14662 11677 14714
rect 18315 14662 18367 14714
rect 18379 14662 18431 14714
rect 18443 14662 18495 14714
rect 18507 14662 18559 14714
rect 18571 14662 18623 14714
rect 25261 14662 25313 14714
rect 25325 14662 25377 14714
rect 25389 14662 25441 14714
rect 25453 14662 25505 14714
rect 25517 14662 25569 14714
rect 1768 14467 1820 14476
rect 1768 14433 1777 14467
rect 1777 14433 1811 14467
rect 1811 14433 1820 14467
rect 1768 14424 1820 14433
rect 2780 14467 2832 14476
rect 2780 14433 2789 14467
rect 2789 14433 2823 14467
rect 2823 14433 2832 14467
rect 2780 14424 2832 14433
rect 9680 14467 9732 14476
rect 9680 14433 9689 14467
rect 9689 14433 9723 14467
rect 9723 14433 9732 14467
rect 9680 14424 9732 14433
rect 20812 14603 20864 14612
rect 1584 14399 1636 14408
rect 1584 14365 1593 14399
rect 1593 14365 1627 14399
rect 1627 14365 1636 14399
rect 1584 14356 1636 14365
rect 8392 14399 8444 14408
rect 8392 14365 8401 14399
rect 8401 14365 8435 14399
rect 8435 14365 8444 14399
rect 8392 14356 8444 14365
rect 12624 14424 12676 14476
rect 12900 14467 12952 14476
rect 12900 14433 12909 14467
rect 12909 14433 12943 14467
rect 12943 14433 12952 14467
rect 12900 14424 12952 14433
rect 13084 14492 13136 14544
rect 14832 14492 14884 14544
rect 16028 14492 16080 14544
rect 18052 14492 18104 14544
rect 20812 14569 20821 14603
rect 20821 14569 20855 14603
rect 20855 14569 20864 14603
rect 20812 14560 20864 14569
rect 26332 14560 26384 14612
rect 14280 14424 14332 14476
rect 13360 14399 13412 14408
rect 10968 14288 11020 14340
rect 11244 14331 11296 14340
rect 11244 14297 11253 14331
rect 11253 14297 11287 14331
rect 11287 14297 11296 14331
rect 11244 14288 11296 14297
rect 12900 14288 12952 14340
rect 13360 14365 13369 14399
rect 13369 14365 13403 14399
rect 13403 14365 13412 14399
rect 13360 14356 13412 14365
rect 18144 14424 18196 14476
rect 14832 14399 14884 14408
rect 14832 14365 14840 14399
rect 14840 14365 14874 14399
rect 14874 14365 14884 14399
rect 14832 14356 14884 14365
rect 15476 14399 15528 14408
rect 13820 14288 13872 14340
rect 14648 14331 14700 14340
rect 14648 14297 14657 14331
rect 14657 14297 14691 14331
rect 14691 14297 14700 14331
rect 14648 14288 14700 14297
rect 15476 14365 15485 14399
rect 15485 14365 15519 14399
rect 15519 14365 15528 14399
rect 15476 14356 15528 14365
rect 15568 14399 15620 14408
rect 15568 14365 15577 14399
rect 15577 14365 15611 14399
rect 15611 14365 15620 14399
rect 15568 14356 15620 14365
rect 15844 14356 15896 14408
rect 18236 14356 18288 14408
rect 23848 14424 23900 14476
rect 24216 14424 24268 14476
rect 27896 14492 27948 14544
rect 26700 14467 26752 14476
rect 26700 14433 26709 14467
rect 26709 14433 26743 14467
rect 26743 14433 26752 14467
rect 26700 14424 26752 14433
rect 19064 14356 19116 14408
rect 21272 14399 21324 14408
rect 21272 14365 21281 14399
rect 21281 14365 21315 14399
rect 21315 14365 21324 14399
rect 21272 14356 21324 14365
rect 28356 14399 28408 14408
rect 28356 14365 28365 14399
rect 28365 14365 28399 14399
rect 28399 14365 28408 14399
rect 28356 14356 28408 14365
rect 9956 14220 10008 14272
rect 13084 14263 13136 14272
rect 13084 14229 13093 14263
rect 13093 14229 13127 14263
rect 13127 14229 13136 14263
rect 13084 14220 13136 14229
rect 13452 14220 13504 14272
rect 16304 14288 16356 14340
rect 19708 14331 19760 14340
rect 19708 14297 19742 14331
rect 19742 14297 19760 14331
rect 19708 14288 19760 14297
rect 21548 14331 21600 14340
rect 21548 14297 21582 14331
rect 21582 14297 21600 14331
rect 21548 14288 21600 14297
rect 24584 14288 24636 14340
rect 18512 14220 18564 14272
rect 22652 14263 22704 14272
rect 22652 14229 22661 14263
rect 22661 14229 22695 14263
rect 22695 14229 22704 14263
rect 22652 14220 22704 14229
rect 25964 14263 26016 14272
rect 25964 14229 25973 14263
rect 25973 14229 26007 14263
rect 26007 14229 26016 14263
rect 25964 14220 26016 14229
rect 7896 14118 7948 14170
rect 7960 14118 8012 14170
rect 8024 14118 8076 14170
rect 8088 14118 8140 14170
rect 8152 14118 8204 14170
rect 14842 14118 14894 14170
rect 14906 14118 14958 14170
rect 14970 14118 15022 14170
rect 15034 14118 15086 14170
rect 15098 14118 15150 14170
rect 21788 14118 21840 14170
rect 21852 14118 21904 14170
rect 21916 14118 21968 14170
rect 21980 14118 22032 14170
rect 22044 14118 22096 14170
rect 28734 14118 28786 14170
rect 28798 14118 28850 14170
rect 28862 14118 28914 14170
rect 28926 14118 28978 14170
rect 28990 14118 29042 14170
rect 9956 13991 10008 14000
rect 9956 13957 9965 13991
rect 9965 13957 9999 13991
rect 9999 13957 10008 13991
rect 9956 13948 10008 13957
rect 1584 13880 1636 13932
rect 3700 13880 3752 13932
rect 13084 14016 13136 14068
rect 15292 14059 15344 14068
rect 15292 14025 15301 14059
rect 15301 14025 15335 14059
rect 15335 14025 15344 14059
rect 15292 14016 15344 14025
rect 16120 14016 16172 14068
rect 16304 14059 16356 14068
rect 16304 14025 16313 14059
rect 16313 14025 16347 14059
rect 16347 14025 16356 14059
rect 16304 14016 16356 14025
rect 18052 14016 18104 14068
rect 19524 14016 19576 14068
rect 27620 14016 27672 14068
rect 3424 13812 3476 13864
rect 8300 13855 8352 13864
rect 8300 13821 8309 13855
rect 8309 13821 8343 13855
rect 8343 13821 8352 13855
rect 8300 13812 8352 13821
rect 10968 13923 11020 13932
rect 10968 13889 10977 13923
rect 10977 13889 11011 13923
rect 11011 13889 11020 13923
rect 10968 13880 11020 13889
rect 14464 13855 14516 13864
rect 14464 13821 14473 13855
rect 14473 13821 14507 13855
rect 14507 13821 14516 13855
rect 14464 13812 14516 13821
rect 15016 13880 15068 13932
rect 15108 13880 15160 13932
rect 16028 13948 16080 14000
rect 16580 13880 16632 13932
rect 17592 13880 17644 13932
rect 18236 13923 18288 13932
rect 18236 13889 18245 13923
rect 18245 13889 18279 13923
rect 18279 13889 18288 13923
rect 19064 13948 19116 14000
rect 21640 13948 21692 14000
rect 18512 13923 18564 13932
rect 18236 13880 18288 13889
rect 18512 13889 18546 13923
rect 18546 13889 18564 13923
rect 18512 13880 18564 13889
rect 21272 13880 21324 13932
rect 24216 13923 24268 13932
rect 24216 13889 24225 13923
rect 24225 13889 24259 13923
rect 24259 13889 24268 13923
rect 24216 13880 24268 13889
rect 24768 13880 24820 13932
rect 27160 13880 27212 13932
rect 28448 13880 28500 13932
rect 14648 13855 14700 13864
rect 14648 13821 14657 13855
rect 14657 13821 14691 13855
rect 14691 13821 14700 13855
rect 14648 13812 14700 13821
rect 17316 13744 17368 13796
rect 16764 13676 16816 13728
rect 23388 13719 23440 13728
rect 23388 13685 23397 13719
rect 23397 13685 23431 13719
rect 23431 13685 23440 13719
rect 23388 13676 23440 13685
rect 25596 13719 25648 13728
rect 25596 13685 25605 13719
rect 25605 13685 25639 13719
rect 25639 13685 25648 13719
rect 25596 13676 25648 13685
rect 26700 13676 26752 13728
rect 4423 13574 4475 13626
rect 4487 13574 4539 13626
rect 4551 13574 4603 13626
rect 4615 13574 4667 13626
rect 4679 13574 4731 13626
rect 11369 13574 11421 13626
rect 11433 13574 11485 13626
rect 11497 13574 11549 13626
rect 11561 13574 11613 13626
rect 11625 13574 11677 13626
rect 18315 13574 18367 13626
rect 18379 13574 18431 13626
rect 18443 13574 18495 13626
rect 18507 13574 18559 13626
rect 18571 13574 18623 13626
rect 25261 13574 25313 13626
rect 25325 13574 25377 13626
rect 25389 13574 25441 13626
rect 25453 13574 25505 13626
rect 25517 13574 25569 13626
rect 11244 13472 11296 13524
rect 14464 13472 14516 13524
rect 16580 13515 16632 13524
rect 16580 13481 16589 13515
rect 16589 13481 16623 13515
rect 16623 13481 16632 13515
rect 16580 13472 16632 13481
rect 19432 13472 19484 13524
rect 19800 13472 19852 13524
rect 1584 13379 1636 13388
rect 1584 13345 1593 13379
rect 1593 13345 1627 13379
rect 1627 13345 1636 13379
rect 1584 13336 1636 13345
rect 3424 13379 3476 13388
rect 3424 13345 3433 13379
rect 3433 13345 3467 13379
rect 3467 13345 3476 13379
rect 3424 13336 3476 13345
rect 26700 13379 26752 13388
rect 26700 13345 26709 13379
rect 26709 13345 26743 13379
rect 26743 13345 26752 13379
rect 26700 13336 26752 13345
rect 28080 13379 28132 13388
rect 28080 13345 28089 13379
rect 28089 13345 28123 13379
rect 28123 13345 28132 13379
rect 28080 13336 28132 13345
rect 9772 13268 9824 13320
rect 13544 13268 13596 13320
rect 14372 13268 14424 13320
rect 14556 13268 14608 13320
rect 14740 13268 14792 13320
rect 15108 13311 15160 13320
rect 15108 13277 15117 13311
rect 15117 13277 15151 13311
rect 15151 13277 15160 13311
rect 15108 13268 15160 13277
rect 16764 13311 16816 13320
rect 16764 13277 16773 13311
rect 16773 13277 16807 13311
rect 16807 13277 16816 13311
rect 16764 13268 16816 13277
rect 2044 13200 2096 13252
rect 15016 13243 15068 13252
rect 15016 13209 15025 13243
rect 15025 13209 15059 13243
rect 15059 13209 15068 13243
rect 15016 13200 15068 13209
rect 7896 13030 7948 13082
rect 7960 13030 8012 13082
rect 8024 13030 8076 13082
rect 8088 13030 8140 13082
rect 8152 13030 8204 13082
rect 14842 13030 14894 13082
rect 14906 13030 14958 13082
rect 14970 13030 15022 13082
rect 15034 13030 15086 13082
rect 15098 13030 15150 13082
rect 21788 13030 21840 13082
rect 21852 13030 21904 13082
rect 21916 13030 21968 13082
rect 21980 13030 22032 13082
rect 22044 13030 22096 13082
rect 28734 13030 28786 13082
rect 28798 13030 28850 13082
rect 28862 13030 28914 13082
rect 28926 13030 28978 13082
rect 28990 13030 29042 13082
rect 2044 12971 2096 12980
rect 2044 12937 2053 12971
rect 2053 12937 2087 12971
rect 2087 12937 2096 12971
rect 2044 12928 2096 12937
rect 19340 12928 19392 12980
rect 24768 12971 24820 12980
rect 24768 12937 24777 12971
rect 24777 12937 24811 12971
rect 24811 12937 24820 12971
rect 24768 12928 24820 12937
rect 2136 12835 2188 12844
rect 2136 12801 2145 12835
rect 2145 12801 2179 12835
rect 2179 12801 2188 12835
rect 2136 12792 2188 12801
rect 19616 12835 19668 12844
rect 19616 12801 19625 12835
rect 19625 12801 19659 12835
rect 19659 12801 19668 12835
rect 19616 12792 19668 12801
rect 22284 12792 22336 12844
rect 22744 12835 22796 12844
rect 22744 12801 22753 12835
rect 22753 12801 22787 12835
rect 22787 12801 22796 12835
rect 22744 12792 22796 12801
rect 24676 12860 24728 12912
rect 24308 12835 24360 12844
rect 24308 12801 24317 12835
rect 24317 12801 24351 12835
rect 24351 12801 24360 12835
rect 24308 12792 24360 12801
rect 24216 12724 24268 12776
rect 24492 12835 24544 12844
rect 24492 12801 24501 12835
rect 24501 12801 24535 12835
rect 24535 12801 24544 12835
rect 24492 12792 24544 12801
rect 27252 12792 27304 12844
rect 25688 12724 25740 12776
rect 26516 12656 26568 12708
rect 23480 12588 23532 12640
rect 23848 12588 23900 12640
rect 24492 12588 24544 12640
rect 26700 12588 26752 12640
rect 4423 12486 4475 12538
rect 4487 12486 4539 12538
rect 4551 12486 4603 12538
rect 4615 12486 4667 12538
rect 4679 12486 4731 12538
rect 11369 12486 11421 12538
rect 11433 12486 11485 12538
rect 11497 12486 11549 12538
rect 11561 12486 11613 12538
rect 11625 12486 11677 12538
rect 18315 12486 18367 12538
rect 18379 12486 18431 12538
rect 18443 12486 18495 12538
rect 18507 12486 18559 12538
rect 18571 12486 18623 12538
rect 25261 12486 25313 12538
rect 25325 12486 25377 12538
rect 25389 12486 25441 12538
rect 25453 12486 25505 12538
rect 25517 12486 25569 12538
rect 3608 12384 3660 12436
rect 9680 12384 9732 12436
rect 19708 12384 19760 12436
rect 21548 12427 21600 12436
rect 21548 12393 21557 12427
rect 21557 12393 21591 12427
rect 21591 12393 21600 12427
rect 21548 12384 21600 12393
rect 23572 12384 23624 12436
rect 24584 12427 24636 12436
rect 24584 12393 24593 12427
rect 24593 12393 24627 12427
rect 24627 12393 24636 12427
rect 24584 12384 24636 12393
rect 25688 12427 25740 12436
rect 25688 12393 25697 12427
rect 25697 12393 25731 12427
rect 25731 12393 25740 12427
rect 25688 12384 25740 12393
rect 20996 12291 21048 12300
rect 20996 12257 21005 12291
rect 21005 12257 21039 12291
rect 21039 12257 21048 12291
rect 20996 12248 21048 12257
rect 22560 12248 22612 12300
rect 19432 12223 19484 12232
rect 19432 12189 19441 12223
rect 19441 12189 19475 12223
rect 19475 12189 19484 12223
rect 19432 12180 19484 12189
rect 20812 12180 20864 12232
rect 21088 12180 21140 12232
rect 22284 12180 22336 12232
rect 22468 12223 22520 12232
rect 22468 12189 22477 12223
rect 22477 12189 22511 12223
rect 22511 12189 22520 12223
rect 23388 12316 23440 12368
rect 22744 12248 22796 12300
rect 23756 12316 23808 12368
rect 24400 12316 24452 12368
rect 24032 12248 24084 12300
rect 24492 12248 24544 12300
rect 26516 12291 26568 12300
rect 22468 12180 22520 12189
rect 22928 12180 22980 12232
rect 23388 12180 23440 12232
rect 23664 12223 23716 12232
rect 23664 12189 23673 12223
rect 23673 12189 23707 12223
rect 23707 12189 23716 12223
rect 23664 12180 23716 12189
rect 24860 12223 24912 12232
rect 20352 12087 20404 12096
rect 20352 12053 20361 12087
rect 20361 12053 20395 12087
rect 20395 12053 20404 12087
rect 20352 12044 20404 12053
rect 22192 12087 22244 12096
rect 22192 12053 22201 12087
rect 22201 12053 22235 12087
rect 22235 12053 22244 12087
rect 22192 12044 22244 12053
rect 22376 12044 22428 12096
rect 22560 12087 22612 12096
rect 22560 12053 22569 12087
rect 22569 12053 22603 12087
rect 22603 12053 22612 12087
rect 22560 12044 22612 12053
rect 23020 12044 23072 12096
rect 23296 12087 23348 12096
rect 23296 12053 23305 12087
rect 23305 12053 23339 12087
rect 23339 12053 23348 12087
rect 23296 12044 23348 12053
rect 23572 12112 23624 12164
rect 24860 12189 24869 12223
rect 24869 12189 24903 12223
rect 24903 12189 24912 12223
rect 24860 12180 24912 12189
rect 26516 12257 26525 12291
rect 26525 12257 26559 12291
rect 26559 12257 26568 12291
rect 26516 12248 26568 12257
rect 26700 12291 26752 12300
rect 26700 12257 26709 12291
rect 26709 12257 26743 12291
rect 26743 12257 26752 12291
rect 26700 12248 26752 12257
rect 28356 12291 28408 12300
rect 28356 12257 28365 12291
rect 28365 12257 28399 12291
rect 28399 12257 28408 12291
rect 28356 12248 28408 12257
rect 25136 12180 25188 12232
rect 24216 12112 24268 12164
rect 25596 12180 25648 12232
rect 25964 12223 26016 12232
rect 25964 12189 25973 12223
rect 25973 12189 26007 12223
rect 26007 12189 26016 12223
rect 25964 12180 26016 12189
rect 7896 11942 7948 11994
rect 7960 11942 8012 11994
rect 8024 11942 8076 11994
rect 8088 11942 8140 11994
rect 8152 11942 8204 11994
rect 14842 11942 14894 11994
rect 14906 11942 14958 11994
rect 14970 11942 15022 11994
rect 15034 11942 15086 11994
rect 15098 11942 15150 11994
rect 21788 11942 21840 11994
rect 21852 11942 21904 11994
rect 21916 11942 21968 11994
rect 21980 11942 22032 11994
rect 22044 11942 22096 11994
rect 28734 11942 28786 11994
rect 28798 11942 28850 11994
rect 28862 11942 28914 11994
rect 28926 11942 28978 11994
rect 28990 11942 29042 11994
rect 19432 11883 19484 11892
rect 19432 11849 19441 11883
rect 19441 11849 19475 11883
rect 19475 11849 19484 11883
rect 19432 11840 19484 11849
rect 20444 11840 20496 11892
rect 21640 11840 21692 11892
rect 22376 11840 22428 11892
rect 23112 11883 23164 11892
rect 23112 11849 23121 11883
rect 23121 11849 23155 11883
rect 23155 11849 23164 11883
rect 23112 11840 23164 11849
rect 23204 11840 23256 11892
rect 20352 11704 20404 11756
rect 23296 11772 23348 11824
rect 24308 11840 24360 11892
rect 24860 11840 24912 11892
rect 23848 11772 23900 11824
rect 24032 11772 24084 11824
rect 1676 11679 1728 11688
rect 1676 11645 1685 11679
rect 1685 11645 1719 11679
rect 1719 11645 1728 11679
rect 1676 11636 1728 11645
rect 2412 11636 2464 11688
rect 2780 11679 2832 11688
rect 2780 11645 2789 11679
rect 2789 11645 2823 11679
rect 2823 11645 2832 11679
rect 2780 11636 2832 11645
rect 19800 11679 19852 11688
rect 19800 11645 19809 11679
rect 19809 11645 19843 11679
rect 19843 11645 19852 11679
rect 19800 11636 19852 11645
rect 20996 11679 21048 11688
rect 20996 11645 21005 11679
rect 21005 11645 21039 11679
rect 21039 11645 21048 11679
rect 20996 11636 21048 11645
rect 19708 11500 19760 11552
rect 23204 11568 23256 11620
rect 23480 11713 23489 11722
rect 23489 11713 23523 11722
rect 23523 11713 23532 11722
rect 23480 11670 23532 11713
rect 23572 11747 23624 11756
rect 23572 11713 23581 11747
rect 23581 11713 23615 11747
rect 23615 11713 23624 11747
rect 23572 11704 23624 11713
rect 24216 11704 24268 11756
rect 24860 11704 24912 11756
rect 25964 11704 26016 11756
rect 24400 11679 24452 11688
rect 24400 11645 24409 11679
rect 24409 11645 24443 11679
rect 24443 11645 24452 11679
rect 24400 11636 24452 11645
rect 24768 11568 24820 11620
rect 23112 11500 23164 11552
rect 25596 11636 25648 11688
rect 4423 11398 4475 11450
rect 4487 11398 4539 11450
rect 4551 11398 4603 11450
rect 4615 11398 4667 11450
rect 4679 11398 4731 11450
rect 11369 11398 11421 11450
rect 11433 11398 11485 11450
rect 11497 11398 11549 11450
rect 11561 11398 11613 11450
rect 11625 11398 11677 11450
rect 18315 11398 18367 11450
rect 18379 11398 18431 11450
rect 18443 11398 18495 11450
rect 18507 11398 18559 11450
rect 18571 11398 18623 11450
rect 25261 11398 25313 11450
rect 25325 11398 25377 11450
rect 25389 11398 25441 11450
rect 25453 11398 25505 11450
rect 25517 11398 25569 11450
rect 1676 11339 1728 11348
rect 1676 11305 1685 11339
rect 1685 11305 1719 11339
rect 1719 11305 1728 11339
rect 1676 11296 1728 11305
rect 2412 11339 2464 11348
rect 2412 11305 2421 11339
rect 2421 11305 2455 11339
rect 2455 11305 2464 11339
rect 2412 11296 2464 11305
rect 19616 11296 19668 11348
rect 22376 11339 22428 11348
rect 22376 11305 22385 11339
rect 22385 11305 22419 11339
rect 22419 11305 22428 11339
rect 22376 11296 22428 11305
rect 23388 11296 23440 11348
rect 23572 11339 23624 11348
rect 23572 11305 23581 11339
rect 23581 11305 23615 11339
rect 23615 11305 23624 11339
rect 23572 11296 23624 11305
rect 25136 11339 25188 11348
rect 25136 11305 25145 11339
rect 25145 11305 25179 11339
rect 25179 11305 25188 11339
rect 25136 11296 25188 11305
rect 23112 11228 23164 11280
rect 20996 11160 21048 11212
rect 2228 11092 2280 11144
rect 9772 11092 9824 11144
rect 19708 11135 19760 11144
rect 19708 11101 19717 11135
rect 19717 11101 19751 11135
rect 19751 11101 19760 11135
rect 19708 11092 19760 11101
rect 19800 11092 19852 11144
rect 20720 11092 20772 11144
rect 22468 11160 22520 11212
rect 23388 11203 23440 11212
rect 23388 11169 23397 11203
rect 23397 11169 23431 11203
rect 23431 11169 23440 11203
rect 24860 11228 24912 11280
rect 24952 11228 25004 11280
rect 23388 11160 23440 11169
rect 25596 11160 25648 11212
rect 27528 11203 27580 11212
rect 27528 11169 27537 11203
rect 27537 11169 27571 11203
rect 27571 11169 27580 11203
rect 27528 11160 27580 11169
rect 22192 11092 22244 11144
rect 24400 11092 24452 11144
rect 22652 11024 22704 11076
rect 23664 11024 23716 11076
rect 24952 11135 25004 11144
rect 24952 11101 24961 11135
rect 24961 11101 24995 11135
rect 24995 11101 25004 11135
rect 24952 11092 25004 11101
rect 28356 11135 28408 11144
rect 28356 11101 28365 11135
rect 28365 11101 28399 11135
rect 28399 11101 28408 11135
rect 28356 11092 28408 11101
rect 27712 11024 27764 11076
rect 20904 10956 20956 11008
rect 23296 10956 23348 11008
rect 7896 10854 7948 10906
rect 7960 10854 8012 10906
rect 8024 10854 8076 10906
rect 8088 10854 8140 10906
rect 8152 10854 8204 10906
rect 14842 10854 14894 10906
rect 14906 10854 14958 10906
rect 14970 10854 15022 10906
rect 15034 10854 15086 10906
rect 15098 10854 15150 10906
rect 21788 10854 21840 10906
rect 21852 10854 21904 10906
rect 21916 10854 21968 10906
rect 21980 10854 22032 10906
rect 22044 10854 22096 10906
rect 28734 10854 28786 10906
rect 28798 10854 28850 10906
rect 28862 10854 28914 10906
rect 28926 10854 28978 10906
rect 28990 10854 29042 10906
rect 21088 10795 21140 10804
rect 21088 10761 21097 10795
rect 21097 10761 21131 10795
rect 21131 10761 21140 10795
rect 21088 10752 21140 10761
rect 22744 10795 22796 10804
rect 22744 10761 22753 10795
rect 22753 10761 22787 10795
rect 22787 10761 22796 10795
rect 22744 10752 22796 10761
rect 13544 10684 13596 10736
rect 22376 10727 22428 10736
rect 20720 10659 20772 10668
rect 20720 10625 20729 10659
rect 20729 10625 20763 10659
rect 20763 10625 20772 10659
rect 20720 10616 20772 10625
rect 20904 10659 20956 10668
rect 20904 10625 20913 10659
rect 20913 10625 20947 10659
rect 20947 10625 20956 10659
rect 20904 10616 20956 10625
rect 22376 10693 22385 10727
rect 22385 10693 22419 10727
rect 22419 10693 22428 10727
rect 22376 10684 22428 10693
rect 23296 10684 23348 10736
rect 28356 10616 28408 10668
rect 22376 10548 22428 10600
rect 22560 10548 22612 10600
rect 23388 10548 23440 10600
rect 23112 10412 23164 10464
rect 26700 10412 26752 10464
rect 27160 10455 27212 10464
rect 27160 10421 27169 10455
rect 27169 10421 27203 10455
rect 27203 10421 27212 10455
rect 27160 10412 27212 10421
rect 4423 10310 4475 10362
rect 4487 10310 4539 10362
rect 4551 10310 4603 10362
rect 4615 10310 4667 10362
rect 4679 10310 4731 10362
rect 11369 10310 11421 10362
rect 11433 10310 11485 10362
rect 11497 10310 11549 10362
rect 11561 10310 11613 10362
rect 11625 10310 11677 10362
rect 18315 10310 18367 10362
rect 18379 10310 18431 10362
rect 18443 10310 18495 10362
rect 18507 10310 18559 10362
rect 18571 10310 18623 10362
rect 25261 10310 25313 10362
rect 25325 10310 25377 10362
rect 25389 10310 25441 10362
rect 25453 10310 25505 10362
rect 25517 10310 25569 10362
rect 27160 10140 27212 10192
rect 26700 10115 26752 10124
rect 26700 10081 26709 10115
rect 26709 10081 26743 10115
rect 26743 10081 26752 10115
rect 26700 10072 26752 10081
rect 29920 10072 29972 10124
rect 1676 10004 1728 10056
rect 3056 10047 3108 10056
rect 3056 10013 3065 10047
rect 3065 10013 3099 10047
rect 3099 10013 3108 10047
rect 3056 10004 3108 10013
rect 7896 9766 7948 9818
rect 7960 9766 8012 9818
rect 8024 9766 8076 9818
rect 8088 9766 8140 9818
rect 8152 9766 8204 9818
rect 14842 9766 14894 9818
rect 14906 9766 14958 9818
rect 14970 9766 15022 9818
rect 15034 9766 15086 9818
rect 15098 9766 15150 9818
rect 21788 9766 21840 9818
rect 21852 9766 21904 9818
rect 21916 9766 21968 9818
rect 21980 9766 22032 9818
rect 22044 9766 22096 9818
rect 28734 9766 28786 9818
rect 28798 9766 28850 9818
rect 28862 9766 28914 9818
rect 28926 9766 28978 9818
rect 28990 9766 29042 9818
rect 2504 9571 2556 9580
rect 2504 9537 2513 9571
rect 2513 9537 2547 9571
rect 2547 9537 2556 9571
rect 25688 9596 25740 9648
rect 27712 9639 27764 9648
rect 27712 9605 27721 9639
rect 27721 9605 27755 9639
rect 27755 9605 27764 9639
rect 27712 9596 27764 9605
rect 3056 9571 3108 9580
rect 2504 9528 2556 9537
rect 3056 9537 3065 9571
rect 3065 9537 3099 9571
rect 3099 9537 3108 9571
rect 3056 9528 3108 9537
rect 21364 9528 21416 9580
rect 27620 9571 27672 9580
rect 27620 9537 27629 9571
rect 27629 9537 27663 9571
rect 27663 9537 27672 9571
rect 27620 9528 27672 9537
rect 4068 9460 4120 9512
rect 4160 9503 4212 9512
rect 4160 9469 4169 9503
rect 4169 9469 4203 9503
rect 4203 9469 4212 9503
rect 4160 9460 4212 9469
rect 1584 9324 1636 9376
rect 1768 9324 1820 9376
rect 25780 9324 25832 9376
rect 4423 9222 4475 9274
rect 4487 9222 4539 9274
rect 4551 9222 4603 9274
rect 4615 9222 4667 9274
rect 4679 9222 4731 9274
rect 11369 9222 11421 9274
rect 11433 9222 11485 9274
rect 11497 9222 11549 9274
rect 11561 9222 11613 9274
rect 11625 9222 11677 9274
rect 18315 9222 18367 9274
rect 18379 9222 18431 9274
rect 18443 9222 18495 9274
rect 18507 9222 18559 9274
rect 18571 9222 18623 9274
rect 25261 9222 25313 9274
rect 25325 9222 25377 9274
rect 25389 9222 25441 9274
rect 25453 9222 25505 9274
rect 25517 9222 25569 9274
rect 4068 9163 4120 9172
rect 4068 9129 4077 9163
rect 4077 9129 4111 9163
rect 4111 9129 4120 9163
rect 4068 9120 4120 9129
rect 1584 9027 1636 9036
rect 1584 8993 1593 9027
rect 1593 8993 1627 9027
rect 1627 8993 1636 9027
rect 1584 8984 1636 8993
rect 1768 9027 1820 9036
rect 1768 8993 1777 9027
rect 1777 8993 1811 9027
rect 1811 8993 1820 9027
rect 1768 8984 1820 8993
rect 2780 9027 2832 9036
rect 2780 8993 2789 9027
rect 2789 8993 2823 9027
rect 2823 8993 2832 9027
rect 2780 8984 2832 8993
rect 25596 9027 25648 9036
rect 25596 8993 25605 9027
rect 25605 8993 25639 9027
rect 25639 8993 25648 9027
rect 25596 8984 25648 8993
rect 25780 9027 25832 9036
rect 25780 8993 25789 9027
rect 25789 8993 25823 9027
rect 25823 8993 25832 9027
rect 25780 8984 25832 8993
rect 4344 8916 4396 8968
rect 28356 8916 28408 8968
rect 29920 8848 29972 8900
rect 7896 8678 7948 8730
rect 7960 8678 8012 8730
rect 8024 8678 8076 8730
rect 8088 8678 8140 8730
rect 8152 8678 8204 8730
rect 14842 8678 14894 8730
rect 14906 8678 14958 8730
rect 14970 8678 15022 8730
rect 15034 8678 15086 8730
rect 15098 8678 15150 8730
rect 21788 8678 21840 8730
rect 21852 8678 21904 8730
rect 21916 8678 21968 8730
rect 21980 8678 22032 8730
rect 22044 8678 22096 8730
rect 28734 8678 28786 8730
rect 28798 8678 28850 8730
rect 28862 8678 28914 8730
rect 28926 8678 28978 8730
rect 28990 8678 29042 8730
rect 1676 8483 1728 8492
rect 1676 8449 1685 8483
rect 1685 8449 1719 8483
rect 1719 8449 1728 8483
rect 1676 8440 1728 8449
rect 12716 8508 12768 8560
rect 1860 8415 1912 8424
rect 1860 8381 1869 8415
rect 1869 8381 1903 8415
rect 1903 8381 1912 8415
rect 1860 8372 1912 8381
rect 2780 8415 2832 8424
rect 2780 8381 2789 8415
rect 2789 8381 2823 8415
rect 2823 8381 2832 8415
rect 2780 8372 2832 8381
rect 4344 8372 4396 8424
rect 27712 8483 27764 8492
rect 27712 8449 27721 8483
rect 27721 8449 27755 8483
rect 27755 8449 27764 8483
rect 27712 8440 27764 8449
rect 28540 8440 28592 8492
rect 9404 8347 9456 8356
rect 9404 8313 9413 8347
rect 9413 8313 9447 8347
rect 9447 8313 9456 8347
rect 9404 8304 9456 8313
rect 3976 8279 4028 8288
rect 3976 8245 3985 8279
rect 3985 8245 4019 8279
rect 4019 8245 4028 8279
rect 3976 8236 4028 8245
rect 4160 8236 4212 8288
rect 26608 8279 26660 8288
rect 26608 8245 26617 8279
rect 26617 8245 26651 8279
rect 26651 8245 26660 8279
rect 26608 8236 26660 8245
rect 28172 8236 28224 8288
rect 4423 8134 4475 8186
rect 4487 8134 4539 8186
rect 4551 8134 4603 8186
rect 4615 8134 4667 8186
rect 4679 8134 4731 8186
rect 11369 8134 11421 8186
rect 11433 8134 11485 8186
rect 11497 8134 11549 8186
rect 11561 8134 11613 8186
rect 11625 8134 11677 8186
rect 18315 8134 18367 8186
rect 18379 8134 18431 8186
rect 18443 8134 18495 8186
rect 18507 8134 18559 8186
rect 18571 8134 18623 8186
rect 25261 8134 25313 8186
rect 25325 8134 25377 8186
rect 25389 8134 25441 8186
rect 25453 8134 25505 8186
rect 25517 8134 25569 8186
rect 1860 8032 1912 8084
rect 3976 7939 4028 7948
rect 3976 7905 3985 7939
rect 3985 7905 4019 7939
rect 4019 7905 4028 7939
rect 3976 7896 4028 7905
rect 4160 7939 4212 7948
rect 4160 7905 4169 7939
rect 4169 7905 4203 7939
rect 4203 7905 4212 7939
rect 4160 7896 4212 7905
rect 5540 7939 5592 7948
rect 5540 7905 5549 7939
rect 5549 7905 5583 7939
rect 5583 7905 5592 7939
rect 5540 7896 5592 7905
rect 27528 7939 27580 7948
rect 27528 7905 27537 7939
rect 27537 7905 27571 7939
rect 27571 7905 27580 7939
rect 27528 7896 27580 7905
rect 28172 7939 28224 7948
rect 28172 7905 28181 7939
rect 28181 7905 28215 7939
rect 28215 7905 28224 7939
rect 28172 7896 28224 7905
rect 28356 7939 28408 7948
rect 28356 7905 28365 7939
rect 28365 7905 28399 7939
rect 28399 7905 28408 7939
rect 28356 7896 28408 7905
rect 2412 7828 2464 7880
rect 7896 7590 7948 7642
rect 7960 7590 8012 7642
rect 8024 7590 8076 7642
rect 8088 7590 8140 7642
rect 8152 7590 8204 7642
rect 14842 7590 14894 7642
rect 14906 7590 14958 7642
rect 14970 7590 15022 7642
rect 15034 7590 15086 7642
rect 15098 7590 15150 7642
rect 21788 7590 21840 7642
rect 21852 7590 21904 7642
rect 21916 7590 21968 7642
rect 21980 7590 22032 7642
rect 22044 7590 22096 7642
rect 28734 7590 28786 7642
rect 28798 7590 28850 7642
rect 28862 7590 28914 7642
rect 28926 7590 28978 7642
rect 28990 7590 29042 7642
rect 2228 7395 2280 7404
rect 2228 7361 2237 7395
rect 2237 7361 2271 7395
rect 2271 7361 2280 7395
rect 2228 7352 2280 7361
rect 26608 7395 26660 7404
rect 26608 7361 26617 7395
rect 26617 7361 26651 7395
rect 26651 7361 26660 7395
rect 26608 7352 26660 7361
rect 28264 7352 28316 7404
rect 26148 7327 26200 7336
rect 26148 7293 26157 7327
rect 26157 7293 26191 7327
rect 26191 7293 26200 7327
rect 26148 7284 26200 7293
rect 1768 7148 1820 7200
rect 2964 7148 3016 7200
rect 4423 7046 4475 7098
rect 4487 7046 4539 7098
rect 4551 7046 4603 7098
rect 4615 7046 4667 7098
rect 4679 7046 4731 7098
rect 11369 7046 11421 7098
rect 11433 7046 11485 7098
rect 11497 7046 11549 7098
rect 11561 7046 11613 7098
rect 11625 7046 11677 7098
rect 18315 7046 18367 7098
rect 18379 7046 18431 7098
rect 18443 7046 18495 7098
rect 18507 7046 18559 7098
rect 18571 7046 18623 7098
rect 25261 7046 25313 7098
rect 25325 7046 25377 7098
rect 25389 7046 25441 7098
rect 25453 7046 25505 7098
rect 25517 7046 25569 7098
rect 1768 6851 1820 6860
rect 1768 6817 1777 6851
rect 1777 6817 1811 6851
rect 1811 6817 1820 6851
rect 1768 6808 1820 6817
rect 2780 6851 2832 6860
rect 2780 6817 2789 6851
rect 2789 6817 2823 6851
rect 2823 6817 2832 6851
rect 2780 6808 2832 6817
rect 19616 6808 19668 6860
rect 25136 6851 25188 6860
rect 25136 6817 25145 6851
rect 25145 6817 25179 6851
rect 25179 6817 25188 6851
rect 25136 6808 25188 6817
rect 1584 6783 1636 6792
rect 1584 6749 1593 6783
rect 1593 6749 1627 6783
rect 1627 6749 1636 6783
rect 1584 6740 1636 6749
rect 26608 6740 26660 6792
rect 23848 6604 23900 6656
rect 27344 6604 27396 6656
rect 7896 6502 7948 6554
rect 7960 6502 8012 6554
rect 8024 6502 8076 6554
rect 8088 6502 8140 6554
rect 8152 6502 8204 6554
rect 14842 6502 14894 6554
rect 14906 6502 14958 6554
rect 14970 6502 15022 6554
rect 15034 6502 15086 6554
rect 15098 6502 15150 6554
rect 21788 6502 21840 6554
rect 21852 6502 21904 6554
rect 21916 6502 21968 6554
rect 21980 6502 22032 6554
rect 22044 6502 22096 6554
rect 28734 6502 28786 6554
rect 28798 6502 28850 6554
rect 28862 6502 28914 6554
rect 28926 6502 28978 6554
rect 28990 6502 29042 6554
rect 1584 6264 1636 6316
rect 2320 6307 2372 6316
rect 2320 6273 2329 6307
rect 2329 6273 2363 6307
rect 2363 6273 2372 6307
rect 2320 6264 2372 6273
rect 2964 6307 3016 6316
rect 2964 6273 2973 6307
rect 2973 6273 3007 6307
rect 3007 6273 3016 6307
rect 2964 6264 3016 6273
rect 26608 6307 26660 6316
rect 26608 6273 26617 6307
rect 26617 6273 26651 6307
rect 26651 6273 26660 6307
rect 26608 6264 26660 6273
rect 27344 6264 27396 6316
rect 4160 6239 4212 6248
rect 4160 6205 4169 6239
rect 4169 6205 4203 6239
rect 4203 6205 4212 6239
rect 4160 6196 4212 6205
rect 26148 6239 26200 6248
rect 26148 6205 26157 6239
rect 26157 6205 26191 6239
rect 26191 6205 26200 6239
rect 26148 6196 26200 6205
rect 5356 6128 5408 6180
rect 4423 5958 4475 6010
rect 4487 5958 4539 6010
rect 4551 5958 4603 6010
rect 4615 5958 4667 6010
rect 4679 5958 4731 6010
rect 11369 5958 11421 6010
rect 11433 5958 11485 6010
rect 11497 5958 11549 6010
rect 11561 5958 11613 6010
rect 11625 5958 11677 6010
rect 18315 5958 18367 6010
rect 18379 5958 18431 6010
rect 18443 5958 18495 6010
rect 18507 5958 18559 6010
rect 18571 5958 18623 6010
rect 25261 5958 25313 6010
rect 25325 5958 25377 6010
rect 25389 5958 25441 6010
rect 25453 5958 25505 6010
rect 25517 5958 25569 6010
rect 25688 5788 25740 5840
rect 3056 5763 3108 5772
rect 3056 5729 3065 5763
rect 3065 5729 3099 5763
rect 3099 5729 3108 5763
rect 3056 5720 3108 5729
rect 27712 5788 27764 5840
rect 1584 5695 1636 5704
rect 1584 5661 1593 5695
rect 1593 5661 1627 5695
rect 1627 5661 1636 5695
rect 1584 5652 1636 5661
rect 4160 5652 4212 5704
rect 24952 5652 25004 5704
rect 26240 5652 26292 5704
rect 26424 5695 26476 5704
rect 26424 5661 26433 5695
rect 26433 5661 26467 5695
rect 26467 5661 26476 5695
rect 26424 5652 26476 5661
rect 1768 5627 1820 5636
rect 1768 5593 1777 5627
rect 1777 5593 1811 5627
rect 1811 5593 1820 5627
rect 1768 5584 1820 5593
rect 26608 5627 26660 5636
rect 26608 5593 26617 5627
rect 26617 5593 26651 5627
rect 26651 5593 26660 5627
rect 26608 5584 26660 5593
rect 29920 5584 29972 5636
rect 7896 5414 7948 5466
rect 7960 5414 8012 5466
rect 8024 5414 8076 5466
rect 8088 5414 8140 5466
rect 8152 5414 8204 5466
rect 14842 5414 14894 5466
rect 14906 5414 14958 5466
rect 14970 5414 15022 5466
rect 15034 5414 15086 5466
rect 15098 5414 15150 5466
rect 21788 5414 21840 5466
rect 21852 5414 21904 5466
rect 21916 5414 21968 5466
rect 21980 5414 22032 5466
rect 22044 5414 22096 5466
rect 28734 5414 28786 5466
rect 28798 5414 28850 5466
rect 28862 5414 28914 5466
rect 28926 5414 28978 5466
rect 28990 5414 29042 5466
rect 1768 5312 1820 5364
rect 26608 5312 26660 5364
rect 2044 5244 2096 5296
rect 1584 5176 1636 5228
rect 10508 5244 10560 5296
rect 26240 5244 26292 5296
rect 5356 5219 5408 5228
rect 5356 5185 5365 5219
rect 5365 5185 5399 5219
rect 5399 5185 5408 5219
rect 5356 5176 5408 5185
rect 27068 5244 27120 5296
rect 26424 5176 26476 5228
rect 2964 5151 3016 5160
rect 2964 5117 2973 5151
rect 2973 5117 3007 5151
rect 3007 5117 3016 5151
rect 2964 5108 3016 5117
rect 3148 5151 3200 5160
rect 3148 5117 3157 5151
rect 3157 5117 3191 5151
rect 3191 5117 3200 5151
rect 3148 5108 3200 5117
rect 4804 5151 4856 5160
rect 4804 5117 4813 5151
rect 4813 5117 4847 5151
rect 4847 5117 4856 5151
rect 4804 5108 4856 5117
rect 5448 5015 5500 5024
rect 5448 4981 5457 5015
rect 5457 4981 5491 5015
rect 5491 4981 5500 5015
rect 5448 4972 5500 4981
rect 26608 4972 26660 5024
rect 4423 4870 4475 4922
rect 4487 4870 4539 4922
rect 4551 4870 4603 4922
rect 4615 4870 4667 4922
rect 4679 4870 4731 4922
rect 11369 4870 11421 4922
rect 11433 4870 11485 4922
rect 11497 4870 11549 4922
rect 11561 4870 11613 4922
rect 11625 4870 11677 4922
rect 18315 4870 18367 4922
rect 18379 4870 18431 4922
rect 18443 4870 18495 4922
rect 18507 4870 18559 4922
rect 18571 4870 18623 4922
rect 25261 4870 25313 4922
rect 25325 4870 25377 4922
rect 25389 4870 25441 4922
rect 25453 4870 25505 4922
rect 25517 4870 25569 4922
rect 2964 4811 3016 4820
rect 2964 4777 2973 4811
rect 2973 4777 3007 4811
rect 3007 4777 3016 4811
rect 2964 4768 3016 4777
rect 5448 4675 5500 4684
rect 5448 4641 5457 4675
rect 5457 4641 5491 4675
rect 5491 4641 5500 4675
rect 5448 4632 5500 4641
rect 5816 4675 5868 4684
rect 5816 4641 5825 4675
rect 5825 4641 5859 4675
rect 5859 4641 5868 4675
rect 5816 4632 5868 4641
rect 25044 4632 25096 4684
rect 27436 4675 27488 4684
rect 27436 4641 27445 4675
rect 27445 4641 27479 4675
rect 27479 4641 27488 4675
rect 27436 4632 27488 4641
rect 1584 4607 1636 4616
rect 1584 4573 1593 4607
rect 1593 4573 1627 4607
rect 1627 4573 1636 4607
rect 1584 4564 1636 4573
rect 2504 4564 2556 4616
rect 3700 4564 3752 4616
rect 28356 4607 28408 4616
rect 28356 4573 28365 4607
rect 28365 4573 28399 4607
rect 28399 4573 28408 4607
rect 28356 4564 28408 4573
rect 22192 4496 22244 4548
rect 23756 4539 23808 4548
rect 23756 4505 23765 4539
rect 23765 4505 23799 4539
rect 23799 4505 23808 4539
rect 23756 4496 23808 4505
rect 28172 4539 28224 4548
rect 28172 4505 28181 4539
rect 28181 4505 28215 4539
rect 28215 4505 28224 4539
rect 28172 4496 28224 4505
rect 1952 4428 2004 4480
rect 7896 4326 7948 4378
rect 7960 4326 8012 4378
rect 8024 4326 8076 4378
rect 8088 4326 8140 4378
rect 8152 4326 8204 4378
rect 14842 4326 14894 4378
rect 14906 4326 14958 4378
rect 14970 4326 15022 4378
rect 15034 4326 15086 4378
rect 15098 4326 15150 4378
rect 21788 4326 21840 4378
rect 21852 4326 21904 4378
rect 21916 4326 21968 4378
rect 21980 4326 22032 4378
rect 22044 4326 22096 4378
rect 28734 4326 28786 4378
rect 28798 4326 28850 4378
rect 28862 4326 28914 4378
rect 28926 4326 28978 4378
rect 28990 4326 29042 4378
rect 2504 4224 2556 4276
rect 4436 4224 4488 4276
rect 28172 4224 28224 4276
rect 2412 4131 2464 4140
rect 2412 4097 2421 4131
rect 2421 4097 2455 4131
rect 2455 4097 2464 4131
rect 2412 4088 2464 4097
rect 3148 4088 3200 4140
rect 3240 4131 3292 4140
rect 3240 4097 3249 4131
rect 3249 4097 3283 4131
rect 3283 4097 3292 4131
rect 3240 4088 3292 4097
rect 3700 4131 3752 4140
rect 3700 4097 3709 4131
rect 3709 4097 3743 4131
rect 3743 4097 3752 4131
rect 3700 4088 3752 4097
rect 10508 4131 10560 4140
rect 4252 4020 4304 4072
rect 10508 4097 10517 4131
rect 10517 4097 10551 4131
rect 10551 4097 10560 4131
rect 10508 4088 10560 4097
rect 2872 3952 2924 4004
rect 11796 4020 11848 4072
rect 12808 4063 12860 4072
rect 12808 4029 12817 4063
rect 12817 4029 12851 4063
rect 12851 4029 12860 4063
rect 12808 4020 12860 4029
rect 12992 4063 13044 4072
rect 12992 4029 13001 4063
rect 13001 4029 13035 4063
rect 13035 4029 13044 4063
rect 12992 4020 13044 4029
rect 13636 4063 13688 4072
rect 13636 4029 13645 4063
rect 13645 4029 13679 4063
rect 13679 4029 13688 4063
rect 13636 4020 13688 4029
rect 4436 3952 4488 4004
rect 18144 3952 18196 4004
rect 21180 4088 21232 4140
rect 22100 4088 22152 4140
rect 23756 4088 23808 4140
rect 27712 4131 27764 4140
rect 27712 4097 27721 4131
rect 27721 4097 27755 4131
rect 27755 4097 27764 4131
rect 27712 4088 27764 4097
rect 24952 4020 25004 4072
rect 1768 3884 1820 3936
rect 4344 3884 4396 3936
rect 5908 3884 5960 3936
rect 6920 3884 6972 3936
rect 10600 3927 10652 3936
rect 10600 3893 10609 3927
rect 10609 3893 10643 3927
rect 10643 3893 10652 3927
rect 10600 3884 10652 3893
rect 19616 3884 19668 3936
rect 20352 3884 20404 3936
rect 20536 3884 20588 3936
rect 27620 3884 27672 3936
rect 4423 3782 4475 3834
rect 4487 3782 4539 3834
rect 4551 3782 4603 3834
rect 4615 3782 4667 3834
rect 4679 3782 4731 3834
rect 11369 3782 11421 3834
rect 11433 3782 11485 3834
rect 11497 3782 11549 3834
rect 11561 3782 11613 3834
rect 11625 3782 11677 3834
rect 18315 3782 18367 3834
rect 18379 3782 18431 3834
rect 18443 3782 18495 3834
rect 18507 3782 18559 3834
rect 18571 3782 18623 3834
rect 25261 3782 25313 3834
rect 25325 3782 25377 3834
rect 25389 3782 25441 3834
rect 25453 3782 25505 3834
rect 25517 3782 25569 3834
rect 4252 3723 4304 3732
rect 4252 3689 4261 3723
rect 4261 3689 4295 3723
rect 4295 3689 4304 3723
rect 4252 3680 4304 3689
rect 12808 3680 12860 3732
rect 664 3612 716 3664
rect 1584 3587 1636 3596
rect 1584 3553 1593 3587
rect 1593 3553 1627 3587
rect 1627 3553 1636 3587
rect 1584 3544 1636 3553
rect 1768 3587 1820 3596
rect 1768 3553 1777 3587
rect 1777 3553 1811 3587
rect 1811 3553 1820 3587
rect 1768 3544 1820 3553
rect 3884 3612 3936 3664
rect 5540 3612 5592 3664
rect 5908 3587 5960 3596
rect 5908 3553 5917 3587
rect 5917 3553 5951 3587
rect 5951 3553 5960 3587
rect 5908 3544 5960 3553
rect 6460 3587 6512 3596
rect 6460 3553 6469 3587
rect 6469 3553 6503 3587
rect 6503 3553 6512 3587
rect 6460 3544 6512 3553
rect 3240 3476 3292 3528
rect 21180 3612 21232 3664
rect 10600 3587 10652 3596
rect 10600 3553 10609 3587
rect 10609 3553 10643 3587
rect 10643 3553 10652 3587
rect 10600 3544 10652 3553
rect 10968 3587 11020 3596
rect 10968 3553 10977 3587
rect 10977 3553 11011 3587
rect 11011 3553 11020 3587
rect 10968 3544 11020 3553
rect 11796 3544 11848 3596
rect 20352 3587 20404 3596
rect 9220 3476 9272 3528
rect 13544 3519 13596 3528
rect 13544 3485 13553 3519
rect 13553 3485 13587 3519
rect 13587 3485 13596 3519
rect 13544 3476 13596 3485
rect 14004 3476 14056 3528
rect 16212 3519 16264 3528
rect 16212 3485 16221 3519
rect 16221 3485 16255 3519
rect 16255 3485 16264 3519
rect 16212 3476 16264 3485
rect 18144 3519 18196 3528
rect 18144 3485 18153 3519
rect 18153 3485 18187 3519
rect 18187 3485 18196 3519
rect 18144 3476 18196 3485
rect 19156 3408 19208 3460
rect 20352 3553 20361 3587
rect 20361 3553 20395 3587
rect 20395 3553 20404 3587
rect 20352 3544 20404 3553
rect 20536 3587 20588 3596
rect 20536 3553 20545 3587
rect 20545 3553 20579 3587
rect 20579 3553 20588 3587
rect 20536 3544 20588 3553
rect 21272 3587 21324 3596
rect 21272 3553 21281 3587
rect 21281 3553 21315 3587
rect 21315 3553 21324 3587
rect 21272 3544 21324 3553
rect 27528 3587 27580 3596
rect 27528 3553 27537 3587
rect 27537 3553 27571 3587
rect 27571 3553 27580 3587
rect 27528 3544 27580 3553
rect 19432 3519 19484 3528
rect 19432 3485 19441 3519
rect 19441 3485 19475 3519
rect 19475 3485 19484 3519
rect 19432 3476 19484 3485
rect 22100 3408 22152 3460
rect 23848 3408 23900 3460
rect 27252 3408 27304 3460
rect 7104 3340 7156 3392
rect 14188 3340 14240 3392
rect 17040 3340 17092 3392
rect 19340 3340 19392 3392
rect 7896 3238 7948 3290
rect 7960 3238 8012 3290
rect 8024 3238 8076 3290
rect 8088 3238 8140 3290
rect 8152 3238 8204 3290
rect 14842 3238 14894 3290
rect 14906 3238 14958 3290
rect 14970 3238 15022 3290
rect 15034 3238 15086 3290
rect 15098 3238 15150 3290
rect 21788 3238 21840 3290
rect 21852 3238 21904 3290
rect 21916 3238 21968 3290
rect 21980 3238 22032 3290
rect 22044 3238 22096 3290
rect 28734 3238 28786 3290
rect 28798 3238 28850 3290
rect 28862 3238 28914 3290
rect 28926 3238 28978 3290
rect 28990 3238 29042 3290
rect 2688 3136 2740 3188
rect 4804 3136 4856 3188
rect 12992 3136 13044 3188
rect 27252 3179 27304 3188
rect 27252 3145 27261 3179
rect 27261 3145 27295 3179
rect 27295 3145 27304 3179
rect 27252 3136 27304 3145
rect 1952 3111 2004 3120
rect 1952 3077 1961 3111
rect 1961 3077 1995 3111
rect 1995 3077 2004 3111
rect 1952 3068 2004 3077
rect 4344 3111 4396 3120
rect 4344 3077 4353 3111
rect 4353 3077 4387 3111
rect 4387 3077 4396 3111
rect 4344 3068 4396 3077
rect 7104 3111 7156 3120
rect 7104 3077 7113 3111
rect 7113 3077 7147 3111
rect 7147 3077 7156 3111
rect 7104 3068 7156 3077
rect 9404 3111 9456 3120
rect 9404 3077 9413 3111
rect 9413 3077 9447 3111
rect 9447 3077 9456 3111
rect 9404 3068 9456 3077
rect 14188 3111 14240 3120
rect 14188 3077 14197 3111
rect 14197 3077 14231 3111
rect 14231 3077 14240 3111
rect 14188 3068 14240 3077
rect 17040 3111 17092 3120
rect 17040 3077 17049 3111
rect 17049 3077 17083 3111
rect 17083 3077 17092 3111
rect 17040 3068 17092 3077
rect 19340 3111 19392 3120
rect 19340 3077 19349 3111
rect 19349 3077 19383 3111
rect 19383 3077 19392 3111
rect 19340 3068 19392 3077
rect 27804 3068 27856 3120
rect 4160 3043 4212 3052
rect 4160 3009 4169 3043
rect 4169 3009 4203 3043
rect 4203 3009 4212 3043
rect 4160 3000 4212 3009
rect 9220 3043 9272 3052
rect 9220 3009 9229 3043
rect 9229 3009 9263 3043
rect 9263 3009 9272 3043
rect 9220 3000 9272 3009
rect 13544 3000 13596 3052
rect 14004 3043 14056 3052
rect 14004 3009 14013 3043
rect 14013 3009 14047 3043
rect 14047 3009 14056 3043
rect 14004 3000 14056 3009
rect 16212 3000 16264 3052
rect 19156 3043 19208 3052
rect 19156 3009 19165 3043
rect 19165 3009 19199 3043
rect 19199 3009 19208 3043
rect 19156 3000 19208 3009
rect 26608 3043 26660 3052
rect 26608 3009 26617 3043
rect 26617 3009 26651 3043
rect 26651 3009 26660 3043
rect 26608 3000 26660 3009
rect 27620 3000 27672 3052
rect 28356 3000 28408 3052
rect 1768 2975 1820 2984
rect 1768 2941 1777 2975
rect 1777 2941 1811 2975
rect 1811 2941 1820 2975
rect 1768 2932 1820 2941
rect 2780 2975 2832 2984
rect 2780 2941 2789 2975
rect 2789 2941 2823 2975
rect 2823 2941 2832 2975
rect 2780 2932 2832 2941
rect 4804 2975 4856 2984
rect 4804 2941 4813 2975
rect 4813 2941 4847 2975
rect 4847 2941 4856 2975
rect 4804 2932 4856 2941
rect 6920 2975 6972 2984
rect 6920 2941 6929 2975
rect 6929 2941 6963 2975
rect 6963 2941 6972 2975
rect 8392 2975 8444 2984
rect 6920 2932 6972 2941
rect 8392 2941 8401 2975
rect 8401 2941 8435 2975
rect 8435 2941 8444 2975
rect 8392 2932 8444 2941
rect 9680 2975 9732 2984
rect 9680 2941 9689 2975
rect 9689 2941 9723 2975
rect 9723 2941 9732 2975
rect 9680 2932 9732 2941
rect 14740 2975 14792 2984
rect 14740 2941 14749 2975
rect 14749 2941 14783 2975
rect 14783 2941 14792 2975
rect 14740 2932 14792 2941
rect 16764 2932 16816 2984
rect 26148 2975 26200 2984
rect 18052 2864 18104 2916
rect 26148 2941 26157 2975
rect 26157 2941 26191 2975
rect 26191 2941 26200 2975
rect 26148 2932 26200 2941
rect 4423 2694 4475 2746
rect 4487 2694 4539 2746
rect 4551 2694 4603 2746
rect 4615 2694 4667 2746
rect 4679 2694 4731 2746
rect 11369 2694 11421 2746
rect 11433 2694 11485 2746
rect 11497 2694 11549 2746
rect 11561 2694 11613 2746
rect 11625 2694 11677 2746
rect 18315 2694 18367 2746
rect 18379 2694 18431 2746
rect 18443 2694 18495 2746
rect 18507 2694 18559 2746
rect 18571 2694 18623 2746
rect 25261 2694 25313 2746
rect 25325 2694 25377 2746
rect 25389 2694 25441 2746
rect 25453 2694 25505 2746
rect 25517 2694 25569 2746
rect 1768 2592 1820 2644
rect 17592 2635 17644 2644
rect 17592 2601 17601 2635
rect 17601 2601 17635 2635
rect 17635 2601 17644 2635
rect 17592 2592 17644 2601
rect 25872 2592 25924 2644
rect 27804 2635 27856 2644
rect 27804 2601 27813 2635
rect 27813 2601 27847 2635
rect 27847 2601 27856 2635
rect 27804 2592 27856 2601
rect 15844 2524 15896 2576
rect 3240 2456 3292 2508
rect 9496 2456 9548 2508
rect 19432 2499 19484 2508
rect 19432 2465 19441 2499
rect 19441 2465 19475 2499
rect 19475 2465 19484 2499
rect 19432 2456 19484 2465
rect 19616 2499 19668 2508
rect 19616 2465 19625 2499
rect 19625 2465 19659 2499
rect 19659 2465 19668 2499
rect 19616 2456 19668 2465
rect 19984 2499 20036 2508
rect 19984 2465 19993 2499
rect 19993 2465 20027 2499
rect 20027 2465 20036 2499
rect 19984 2456 20036 2465
rect 2596 2431 2648 2440
rect 2596 2397 2605 2431
rect 2605 2397 2639 2431
rect 2639 2397 2648 2431
rect 2596 2388 2648 2397
rect 9036 2388 9088 2440
rect 17408 2388 17460 2440
rect 27068 2388 27120 2440
rect 27620 2388 27672 2440
rect 16120 2320 16172 2372
rect 3516 2252 3568 2304
rect 8300 2252 8352 2304
rect 7896 2150 7948 2202
rect 7960 2150 8012 2202
rect 8024 2150 8076 2202
rect 8088 2150 8140 2202
rect 8152 2150 8204 2202
rect 14842 2150 14894 2202
rect 14906 2150 14958 2202
rect 14970 2150 15022 2202
rect 15034 2150 15086 2202
rect 15098 2150 15150 2202
rect 21788 2150 21840 2202
rect 21852 2150 21904 2202
rect 21916 2150 21968 2202
rect 21980 2150 22032 2202
rect 22044 2150 22096 2202
rect 28734 2150 28786 2202
rect 28798 2150 28850 2202
rect 28862 2150 28914 2202
rect 28926 2150 28978 2202
rect 28990 2150 29042 2202
<< metal2 >>
rect -10 49200 102 49800
rect 634 49314 746 49800
rect 1278 49314 1390 49800
rect 634 49286 1072 49314
rect 634 49200 746 49286
rect 1044 46034 1072 49286
rect 1136 49286 1390 49314
rect 1032 46028 1084 46034
rect 1032 45970 1084 45976
rect 1136 45554 1164 49286
rect 1278 49200 1390 49286
rect 1922 49200 2034 49800
rect 2566 49200 2678 49800
rect 3210 49200 3322 49800
rect 3514 49736 3570 49745
rect 3514 49671 3570 49680
rect 1964 46510 1992 49200
rect 2228 47048 2280 47054
rect 2228 46990 2280 46996
rect 2240 46578 2268 46990
rect 2228 46572 2280 46578
rect 2228 46514 2280 46520
rect 1952 46504 2004 46510
rect 1952 46446 2004 46452
rect 1676 46368 1728 46374
rect 1676 46310 1728 46316
rect 32 45526 1164 45554
rect 32 45354 60 45526
rect 1688 45490 1716 46310
rect 2608 46034 2636 49200
rect 2872 47048 2924 47054
rect 2872 46990 2924 46996
rect 2780 46912 2832 46918
rect 2780 46854 2832 46860
rect 2792 46646 2820 46854
rect 2780 46640 2832 46646
rect 2780 46582 2832 46588
rect 2596 46028 2648 46034
rect 2596 45970 2648 45976
rect 1676 45484 1728 45490
rect 1676 45426 1728 45432
rect 2044 45416 2096 45422
rect 2044 45358 2096 45364
rect 2504 45416 2556 45422
rect 2504 45358 2556 45364
rect 20 45348 72 45354
rect 20 45290 72 45296
rect 2056 45082 2084 45358
rect 2044 45076 2096 45082
rect 2044 45018 2096 45024
rect 2516 44878 2544 45358
rect 2778 44976 2834 44985
rect 2778 44911 2834 44920
rect 2504 44872 2556 44878
rect 2504 44814 2556 44820
rect 1584 43784 1636 43790
rect 1584 43726 1636 43732
rect 1596 42770 1624 43726
rect 1768 43104 1820 43110
rect 1768 43046 1820 43052
rect 1780 42770 1808 43046
rect 1584 42764 1636 42770
rect 1584 42706 1636 42712
rect 1768 42764 1820 42770
rect 1768 42706 1820 42712
rect 1676 42016 1728 42022
rect 1676 41958 1728 41964
rect 1584 41608 1636 41614
rect 1582 41576 1584 41585
rect 1636 41576 1638 41585
rect 1582 41511 1638 41520
rect 1688 41138 1716 41958
rect 1676 41132 1728 41138
rect 1676 41074 1728 41080
rect 2320 41064 2372 41070
rect 2320 41006 2372 41012
rect 1952 40520 2004 40526
rect 1952 40462 2004 40468
rect 1860 40384 1912 40390
rect 1860 40326 1912 40332
rect 1872 40118 1900 40326
rect 1860 40112 1912 40118
rect 1860 40054 1912 40060
rect 1964 39506 1992 40462
rect 2332 39642 2360 41006
rect 2412 40520 2464 40526
rect 2412 40462 2464 40468
rect 2424 39982 2452 40462
rect 2412 39976 2464 39982
rect 2412 39918 2464 39924
rect 2320 39636 2372 39642
rect 2320 39578 2372 39584
rect 1952 39500 2004 39506
rect 1952 39442 2004 39448
rect 1676 38344 1728 38350
rect 1676 38286 1728 38292
rect 1582 37496 1638 37505
rect 1582 37431 1638 37440
rect 1596 37262 1624 37431
rect 1584 37256 1636 37262
rect 1584 37198 1636 37204
rect 1688 36310 1716 38286
rect 1768 36576 1820 36582
rect 1768 36518 1820 36524
rect 1676 36304 1728 36310
rect 1676 36246 1728 36252
rect 1780 36242 1808 36518
rect 1768 36236 1820 36242
rect 1768 36178 1820 36184
rect 1676 35080 1728 35086
rect 1676 35022 1728 35028
rect 1688 34610 1716 35022
rect 1676 34604 1728 34610
rect 1676 34546 1728 34552
rect 1860 34536 1912 34542
rect 1860 34478 1912 34484
rect 1872 34202 1900 34478
rect 1860 34196 1912 34202
rect 1860 34138 1912 34144
rect 1584 30184 1636 30190
rect 1584 30126 1636 30132
rect 1860 30184 1912 30190
rect 1860 30126 1912 30132
rect 1596 30025 1624 30126
rect 1582 30016 1638 30025
rect 1582 29951 1638 29960
rect 1584 28076 1636 28082
rect 1584 28018 1636 28024
rect 1596 27985 1624 28018
rect 1582 27976 1638 27985
rect 1582 27911 1638 27920
rect 1768 27872 1820 27878
rect 1768 27814 1820 27820
rect 1780 27402 1808 27814
rect 1768 27396 1820 27402
rect 1768 27338 1820 27344
rect 1872 27282 1900 30126
rect 1780 27254 1900 27282
rect 1676 25832 1728 25838
rect 1676 25774 1728 25780
rect 1688 25498 1716 25774
rect 1676 25492 1728 25498
rect 1676 25434 1728 25440
rect 1582 25256 1638 25265
rect 1582 25191 1638 25200
rect 1596 24818 1624 25191
rect 1584 24812 1636 24818
rect 1584 24754 1636 24760
rect 1780 22094 1808 27254
rect 1860 26240 1912 26246
rect 1860 26182 1912 26188
rect 1872 25974 1900 26182
rect 1860 25968 1912 25974
rect 1860 25910 1912 25916
rect 1964 22094 1992 39442
rect 2516 35894 2544 44814
rect 2792 42770 2820 44911
rect 2780 42764 2832 42770
rect 2780 42706 2832 42712
rect 2778 42256 2834 42265
rect 2884 42226 2912 46990
rect 3424 45960 3476 45966
rect 3424 45902 3476 45908
rect 3240 45892 3292 45898
rect 3240 45834 3292 45840
rect 3252 44538 3280 45834
rect 3240 44532 3292 44538
rect 3240 44474 3292 44480
rect 2964 44192 3016 44198
rect 2964 44134 3016 44140
rect 2976 43314 3004 44134
rect 3436 43994 3464 45902
rect 3424 43988 3476 43994
rect 3424 43930 3476 43936
rect 3148 43648 3200 43654
rect 3148 43590 3200 43596
rect 3056 43444 3108 43450
rect 3056 43386 3108 43392
rect 2964 43308 3016 43314
rect 2964 43250 3016 43256
rect 3068 43178 3096 43386
rect 3160 43382 3188 43590
rect 3148 43376 3200 43382
rect 3148 43318 3200 43324
rect 3056 43172 3108 43178
rect 3056 43114 3108 43120
rect 2778 42191 2834 42200
rect 2872 42220 2924 42226
rect 2792 41070 2820 42191
rect 2872 42162 2924 42168
rect 2780 41064 2832 41070
rect 2780 41006 2832 41012
rect 2872 39364 2924 39370
rect 2872 39306 2924 39312
rect 2778 38856 2834 38865
rect 2778 38791 2834 38800
rect 2792 37806 2820 38791
rect 2780 37800 2832 37806
rect 2780 37742 2832 37748
rect 2884 36825 2912 39306
rect 2870 36816 2926 36825
rect 2870 36751 2926 36760
rect 2596 36712 2648 36718
rect 2596 36654 2648 36660
rect 2148 35866 2544 35894
rect 1780 22066 1900 22094
rect 1964 22066 2084 22094
rect 1768 20256 1820 20262
rect 1768 20198 1820 20204
rect 1780 19922 1808 20198
rect 1768 19916 1820 19922
rect 1768 19858 1820 19864
rect 1584 19848 1636 19854
rect 1584 19790 1636 19796
rect 1596 19378 1624 19790
rect 1584 19372 1636 19378
rect 1584 19314 1636 19320
rect 1584 18760 1636 18766
rect 1584 18702 1636 18708
rect 1596 18465 1624 18702
rect 1582 18456 1638 18465
rect 1582 18391 1638 18400
rect 1584 18080 1636 18086
rect 1584 18022 1636 18028
rect 1596 17746 1624 18022
rect 1872 17814 1900 22066
rect 2056 20466 2084 22066
rect 2044 20460 2096 20466
rect 2044 20402 2096 20408
rect 1860 17808 1912 17814
rect 1860 17750 1912 17756
rect 1584 17740 1636 17746
rect 1584 17682 1636 17688
rect 1952 17604 2004 17610
rect 1952 17546 2004 17552
rect 1964 17338 1992 17546
rect 1952 17332 2004 17338
rect 1952 17274 2004 17280
rect 2056 17202 2084 20402
rect 2044 17196 2096 17202
rect 2044 17138 2096 17144
rect 1860 16448 1912 16454
rect 1860 16390 1912 16396
rect 1872 16182 1900 16390
rect 1860 16176 1912 16182
rect 1860 16118 1912 16124
rect 1676 16040 1728 16046
rect 1676 15982 1728 15988
rect 1688 15706 1716 15982
rect 1676 15700 1728 15706
rect 1676 15642 1728 15648
rect 2056 15026 2084 17138
rect 2044 15020 2096 15026
rect 2044 14962 2096 14968
rect 1768 14816 1820 14822
rect 1768 14758 1820 14764
rect 1780 14482 1808 14758
rect 1768 14476 1820 14482
rect 1768 14418 1820 14424
rect 1584 14408 1636 14414
rect 1584 14350 1636 14356
rect 1596 13938 1624 14350
rect 1584 13932 1636 13938
rect 1584 13874 1636 13880
rect 1582 13696 1638 13705
rect 1582 13631 1638 13640
rect 1596 13394 1624 13631
rect 1584 13388 1636 13394
rect 1584 13330 1636 13336
rect 2044 13252 2096 13258
rect 2044 13194 2096 13200
rect 2056 12986 2084 13194
rect 2044 12980 2096 12986
rect 2044 12922 2096 12928
rect 2148 12850 2176 35866
rect 2332 35766 2360 35866
rect 2320 35760 2372 35766
rect 2320 35702 2372 35708
rect 2608 35698 2636 36654
rect 2780 36236 2832 36242
rect 2780 36178 2832 36184
rect 2792 36145 2820 36178
rect 2778 36136 2834 36145
rect 2778 36071 2834 36080
rect 3068 35894 3096 43114
rect 3240 42016 3292 42022
rect 3240 41958 3292 41964
rect 3424 42016 3476 42022
rect 3424 41958 3476 41964
rect 3252 41682 3280 41958
rect 3436 41682 3464 41958
rect 3240 41676 3292 41682
rect 3240 41618 3292 41624
rect 3424 41676 3476 41682
rect 3424 41618 3476 41624
rect 3528 40118 3556 49671
rect 4498 49200 4610 49800
rect 5142 49200 5254 49800
rect 5786 49200 5898 49800
rect 6430 49200 6542 49800
rect 7074 49200 7186 49800
rect 7718 49200 7830 49800
rect 8362 49200 8474 49800
rect 9650 49200 9762 49800
rect 10294 49200 10406 49800
rect 10938 49200 11050 49800
rect 11582 49200 11694 49800
rect 12226 49200 12338 49800
rect 12870 49200 12982 49800
rect 13514 49200 13626 49800
rect 14802 49314 14914 49800
rect 14802 49286 15148 49314
rect 14802 49200 14914 49286
rect 4423 47356 4731 47365
rect 4423 47354 4429 47356
rect 4485 47354 4509 47356
rect 4565 47354 4589 47356
rect 4645 47354 4669 47356
rect 4725 47354 4731 47356
rect 4485 47302 4487 47354
rect 4667 47302 4669 47354
rect 4423 47300 4429 47302
rect 4485 47300 4509 47302
rect 4565 47300 4589 47302
rect 4645 47300 4669 47302
rect 4725 47300 4731 47302
rect 4423 47291 4731 47300
rect 5828 47054 5856 49200
rect 6472 47054 6500 49200
rect 5816 47048 5868 47054
rect 5816 46990 5868 46996
rect 6460 47048 6512 47054
rect 6460 46990 6512 46996
rect 7012 47048 7064 47054
rect 7012 46990 7064 46996
rect 6000 46912 6052 46918
rect 6000 46854 6052 46860
rect 6736 46912 6788 46918
rect 6736 46854 6788 46860
rect 4423 46268 4731 46277
rect 4423 46266 4429 46268
rect 4485 46266 4509 46268
rect 4565 46266 4589 46268
rect 4645 46266 4669 46268
rect 4725 46266 4731 46268
rect 4485 46214 4487 46266
rect 4667 46214 4669 46266
rect 4423 46212 4429 46214
rect 4485 46212 4509 46214
rect 4565 46212 4589 46214
rect 4645 46212 4669 46214
rect 4725 46212 4731 46214
rect 4423 46203 4731 46212
rect 3976 45960 4028 45966
rect 3976 45902 4028 45908
rect 3988 45082 4016 45902
rect 4160 45892 4212 45898
rect 4160 45834 4212 45840
rect 4172 45558 4200 45834
rect 4160 45552 4212 45558
rect 4160 45494 4212 45500
rect 4423 45180 4731 45189
rect 4423 45178 4429 45180
rect 4485 45178 4509 45180
rect 4565 45178 4589 45180
rect 4645 45178 4669 45180
rect 4725 45178 4731 45180
rect 4485 45126 4487 45178
rect 4667 45126 4669 45178
rect 4423 45124 4429 45126
rect 4485 45124 4509 45126
rect 4565 45124 4589 45126
rect 4645 45124 4669 45126
rect 4725 45124 4731 45126
rect 4423 45115 4731 45124
rect 3976 45076 4028 45082
rect 3976 45018 4028 45024
rect 5172 44872 5224 44878
rect 5172 44814 5224 44820
rect 5184 44402 5212 44814
rect 4344 44396 4396 44402
rect 4344 44338 4396 44344
rect 5172 44396 5224 44402
rect 5172 44338 5224 44344
rect 4158 44296 4214 44305
rect 4158 44231 4214 44240
rect 4172 43246 4200 44231
rect 4160 43240 4212 43246
rect 4160 43182 4212 43188
rect 3516 40112 3568 40118
rect 3516 40054 3568 40060
rect 3148 39296 3200 39302
rect 3148 39238 3200 39244
rect 3160 37194 3188 39238
rect 3424 38820 3476 38826
rect 3424 38762 3476 38768
rect 3240 38208 3292 38214
rect 3240 38150 3292 38156
rect 3252 37330 3280 38150
rect 3240 37324 3292 37330
rect 3240 37266 3292 37272
rect 3436 37262 3464 38762
rect 3976 38752 4028 38758
rect 3976 38694 4028 38700
rect 3988 37874 4016 38694
rect 3976 37868 4028 37874
rect 3976 37810 4028 37816
rect 3424 37256 3476 37262
rect 3424 37198 3476 37204
rect 3148 37188 3200 37194
rect 3148 37130 3200 37136
rect 4160 37188 4212 37194
rect 4160 37130 4212 37136
rect 3160 36854 3188 37130
rect 4172 36922 4200 37130
rect 4160 36916 4212 36922
rect 4160 36858 4212 36864
rect 4356 36854 4384 44338
rect 4423 44092 4731 44101
rect 4423 44090 4429 44092
rect 4485 44090 4509 44092
rect 4565 44090 4589 44092
rect 4645 44090 4669 44092
rect 4725 44090 4731 44092
rect 4485 44038 4487 44090
rect 4667 44038 4669 44090
rect 4423 44036 4429 44038
rect 4485 44036 4509 44038
rect 4565 44036 4589 44038
rect 4645 44036 4669 44038
rect 4725 44036 4731 44038
rect 4423 44027 4731 44036
rect 5080 43784 5132 43790
rect 5080 43726 5132 43732
rect 4423 43004 4731 43013
rect 4423 43002 4429 43004
rect 4485 43002 4509 43004
rect 4565 43002 4589 43004
rect 4645 43002 4669 43004
rect 4725 43002 4731 43004
rect 4485 42950 4487 43002
rect 4667 42950 4669 43002
rect 4423 42948 4429 42950
rect 4485 42948 4509 42950
rect 4565 42948 4589 42950
rect 4645 42948 4669 42950
rect 4725 42948 4731 42950
rect 4423 42939 4731 42948
rect 4423 41916 4731 41925
rect 4423 41914 4429 41916
rect 4485 41914 4509 41916
rect 4565 41914 4589 41916
rect 4645 41914 4669 41916
rect 4725 41914 4731 41916
rect 4485 41862 4487 41914
rect 4667 41862 4669 41914
rect 4423 41860 4429 41862
rect 4485 41860 4509 41862
rect 4565 41860 4589 41862
rect 4645 41860 4669 41862
rect 4725 41860 4731 41862
rect 4423 41851 4731 41860
rect 4423 40828 4731 40837
rect 4423 40826 4429 40828
rect 4485 40826 4509 40828
rect 4565 40826 4589 40828
rect 4645 40826 4669 40828
rect 4725 40826 4731 40828
rect 4485 40774 4487 40826
rect 4667 40774 4669 40826
rect 4423 40772 4429 40774
rect 4485 40772 4509 40774
rect 4565 40772 4589 40774
rect 4645 40772 4669 40774
rect 4725 40772 4731 40774
rect 4423 40763 4731 40772
rect 4423 39740 4731 39749
rect 4423 39738 4429 39740
rect 4485 39738 4509 39740
rect 4565 39738 4589 39740
rect 4645 39738 4669 39740
rect 4725 39738 4731 39740
rect 4485 39686 4487 39738
rect 4667 39686 4669 39738
rect 4423 39684 4429 39686
rect 4485 39684 4509 39686
rect 4565 39684 4589 39686
rect 4645 39684 4669 39686
rect 4725 39684 4731 39686
rect 4423 39675 4731 39684
rect 4423 38652 4731 38661
rect 4423 38650 4429 38652
rect 4485 38650 4509 38652
rect 4565 38650 4589 38652
rect 4645 38650 4669 38652
rect 4725 38650 4731 38652
rect 4485 38598 4487 38650
rect 4667 38598 4669 38650
rect 4423 38596 4429 38598
rect 4485 38596 4509 38598
rect 4565 38596 4589 38598
rect 4645 38596 4669 38598
rect 4725 38596 4731 38598
rect 4423 38587 4731 38596
rect 4896 37868 4948 37874
rect 4896 37810 4948 37816
rect 4423 37564 4731 37573
rect 4423 37562 4429 37564
rect 4485 37562 4509 37564
rect 4565 37562 4589 37564
rect 4645 37562 4669 37564
rect 4725 37562 4731 37564
rect 4485 37510 4487 37562
rect 4667 37510 4669 37562
rect 4423 37508 4429 37510
rect 4485 37508 4509 37510
rect 4565 37508 4589 37510
rect 4645 37508 4669 37510
rect 4725 37508 4731 37510
rect 4423 37499 4731 37508
rect 3148 36848 3200 36854
rect 3148 36790 3200 36796
rect 4344 36848 4396 36854
rect 4344 36790 4396 36796
rect 4252 36780 4304 36786
rect 4252 36722 4304 36728
rect 4160 36644 4212 36650
rect 4160 36586 4212 36592
rect 2884 35866 3096 35894
rect 2596 35692 2648 35698
rect 2596 35634 2648 35640
rect 2884 35154 2912 35866
rect 4172 35630 4200 36586
rect 4264 36174 4292 36722
rect 4344 36712 4396 36718
rect 4344 36654 4396 36660
rect 4252 36168 4304 36174
rect 4252 36110 4304 36116
rect 4264 35698 4292 36110
rect 4252 35692 4304 35698
rect 4252 35634 4304 35640
rect 4160 35624 4212 35630
rect 4160 35566 4212 35572
rect 2872 35148 2924 35154
rect 2872 35090 2924 35096
rect 2778 34776 2834 34785
rect 2778 34711 2834 34720
rect 2792 34542 2820 34711
rect 2780 34536 2832 34542
rect 2780 34478 2832 34484
rect 2884 33998 2912 35090
rect 4264 35086 4292 35634
rect 4356 35154 4384 36654
rect 4423 36476 4731 36485
rect 4423 36474 4429 36476
rect 4485 36474 4509 36476
rect 4565 36474 4589 36476
rect 4645 36474 4669 36476
rect 4725 36474 4731 36476
rect 4485 36422 4487 36474
rect 4667 36422 4669 36474
rect 4423 36420 4429 36422
rect 4485 36420 4509 36422
rect 4565 36420 4589 36422
rect 4645 36420 4669 36422
rect 4725 36420 4731 36422
rect 4423 36411 4731 36420
rect 4908 36106 4936 37810
rect 4988 36848 5040 36854
rect 4988 36790 5040 36796
rect 5000 36378 5028 36790
rect 4988 36372 5040 36378
rect 4988 36314 5040 36320
rect 4896 36100 4948 36106
rect 4896 36042 4948 36048
rect 4804 35624 4856 35630
rect 4804 35566 4856 35572
rect 4423 35388 4731 35397
rect 4423 35386 4429 35388
rect 4485 35386 4509 35388
rect 4565 35386 4589 35388
rect 4645 35386 4669 35388
rect 4725 35386 4731 35388
rect 4485 35334 4487 35386
rect 4667 35334 4669 35386
rect 4423 35332 4429 35334
rect 4485 35332 4509 35334
rect 4565 35332 4589 35334
rect 4645 35332 4669 35334
rect 4725 35332 4731 35334
rect 4423 35323 4731 35332
rect 4344 35148 4396 35154
rect 4344 35090 4396 35096
rect 4252 35080 4304 35086
rect 4252 35022 4304 35028
rect 4264 34610 4292 35022
rect 4356 35018 4384 35090
rect 4344 35012 4396 35018
rect 4344 34954 4396 34960
rect 4252 34604 4304 34610
rect 4252 34546 4304 34552
rect 4264 33998 4292 34546
rect 2320 33992 2372 33998
rect 2320 33934 2372 33940
rect 2872 33992 2924 33998
rect 2872 33934 2924 33940
rect 4252 33992 4304 33998
rect 4252 33934 4304 33940
rect 2228 17876 2280 17882
rect 2228 17818 2280 17824
rect 2240 16658 2268 17818
rect 2228 16652 2280 16658
rect 2228 16594 2280 16600
rect 2136 12844 2188 12850
rect 2136 12786 2188 12792
rect 2148 12434 2176 12786
rect 2056 12406 2176 12434
rect 1676 11688 1728 11694
rect 1676 11630 1728 11636
rect 1688 11354 1716 11630
rect 1676 11348 1728 11354
rect 1676 11290 1728 11296
rect 1676 10056 1728 10062
rect 1676 9998 1728 10004
rect 1584 9376 1636 9382
rect 1584 9318 1636 9324
rect 1596 9042 1624 9318
rect 1584 9036 1636 9042
rect 1584 8978 1636 8984
rect 1688 8498 1716 9998
rect 1768 9376 1820 9382
rect 1768 9318 1820 9324
rect 1780 9042 1808 9318
rect 1768 9036 1820 9042
rect 1768 8978 1820 8984
rect 1676 8492 1728 8498
rect 1676 8434 1728 8440
rect 1860 8424 1912 8430
rect 1860 8366 1912 8372
rect 1872 8090 1900 8366
rect 1860 8084 1912 8090
rect 1860 8026 1912 8032
rect 1768 7200 1820 7206
rect 1768 7142 1820 7148
rect 1780 6866 1808 7142
rect 1768 6860 1820 6866
rect 1768 6802 1820 6808
rect 1584 6792 1636 6798
rect 1584 6734 1636 6740
rect 1596 6322 1624 6734
rect 1584 6316 1636 6322
rect 1584 6258 1636 6264
rect 1584 5704 1636 5710
rect 1584 5646 1636 5652
rect 1596 5234 1624 5646
rect 1768 5636 1820 5642
rect 1768 5578 1820 5584
rect 1780 5370 1808 5578
rect 1768 5364 1820 5370
rect 1768 5306 1820 5312
rect 2056 5302 2084 12406
rect 2240 11150 2268 16594
rect 2228 11144 2280 11150
rect 2228 11086 2280 11092
rect 2240 7410 2268 11086
rect 2228 7404 2280 7410
rect 2228 7346 2280 7352
rect 2332 6322 2360 33934
rect 4160 33924 4212 33930
rect 4160 33866 4212 33872
rect 3514 33416 3570 33425
rect 3514 33351 3570 33360
rect 3528 33318 3556 33351
rect 3516 33312 3568 33318
rect 3516 33254 3568 33260
rect 2962 32056 3018 32065
rect 2962 31991 3018 32000
rect 2976 28014 3004 31991
rect 2964 28008 3016 28014
rect 2964 27950 3016 27956
rect 2596 27600 2648 27606
rect 2596 27542 2648 27548
rect 2608 26382 2636 27542
rect 2596 26376 2648 26382
rect 2596 26318 2648 26324
rect 2504 15020 2556 15026
rect 2504 14962 2556 14968
rect 2412 11688 2464 11694
rect 2412 11630 2464 11636
rect 2424 11354 2452 11630
rect 2412 11348 2464 11354
rect 2412 11290 2464 11296
rect 2516 9586 2544 14962
rect 2504 9580 2556 9586
rect 2504 9522 2556 9528
rect 2412 7880 2464 7886
rect 2412 7822 2464 7828
rect 2320 6316 2372 6322
rect 2320 6258 2372 6264
rect 2044 5296 2096 5302
rect 2044 5238 2096 5244
rect 1584 5228 1636 5234
rect 1584 5170 1636 5176
rect 1584 4616 1636 4622
rect 1584 4558 1636 4564
rect 664 3664 716 3670
rect 664 3606 716 3612
rect 676 800 704 3606
rect 1596 3602 1624 4558
rect 1952 4480 2004 4486
rect 1952 4422 2004 4428
rect 1768 3936 1820 3942
rect 1768 3878 1820 3884
rect 1780 3602 1808 3878
rect 1584 3596 1636 3602
rect 1584 3538 1636 3544
rect 1768 3596 1820 3602
rect 1768 3538 1820 3544
rect 1964 3126 1992 4422
rect 2424 4146 2452 7822
rect 2504 4616 2556 4622
rect 2504 4558 2556 4564
rect 2516 4282 2544 4558
rect 2504 4276 2556 4282
rect 2504 4218 2556 4224
rect 2412 4140 2464 4146
rect 2412 4082 2464 4088
rect 1952 3120 2004 3126
rect 1952 3062 2004 3068
rect 1768 2984 1820 2990
rect 1768 2926 1820 2932
rect 1780 2650 1808 2926
rect 1768 2644 1820 2650
rect 1768 2586 1820 2592
rect 2608 2446 2636 26318
rect 2778 25936 2834 25945
rect 2778 25871 2834 25880
rect 2792 25838 2820 25871
rect 2780 25832 2832 25838
rect 2780 25774 2832 25780
rect 2780 19916 2832 19922
rect 2780 19858 2832 19864
rect 2792 19825 2820 19858
rect 2778 19816 2834 19825
rect 2778 19751 2834 19760
rect 3330 19136 3386 19145
rect 3330 19071 3386 19080
rect 3344 18698 3372 19071
rect 3332 18692 3384 18698
rect 3332 18634 3384 18640
rect 2778 17776 2834 17785
rect 2778 17711 2780 17720
rect 2832 17711 2834 17720
rect 2780 17682 2832 17688
rect 2780 16040 2832 16046
rect 2780 15982 2832 15988
rect 2792 15745 2820 15982
rect 2778 15736 2834 15745
rect 2778 15671 2834 15680
rect 2780 14476 2832 14482
rect 2780 14418 2832 14424
rect 2792 14385 2820 14418
rect 2778 14376 2834 14385
rect 2778 14311 2834 14320
rect 3700 13932 3752 13938
rect 3700 13874 3752 13880
rect 3424 13864 3476 13870
rect 3424 13806 3476 13812
rect 3436 13394 3464 13806
rect 3424 13388 3476 13394
rect 3424 13330 3476 13336
rect 3608 12436 3660 12442
rect 3608 12378 3660 12384
rect 3620 12345 3648 12378
rect 3606 12336 3662 12345
rect 3606 12271 3662 12280
rect 2780 11688 2832 11694
rect 2778 11656 2780 11665
rect 2832 11656 2834 11665
rect 2778 11591 2834 11600
rect 3056 10056 3108 10062
rect 3056 9998 3108 10004
rect 3068 9586 3096 9998
rect 3056 9580 3108 9586
rect 3056 9522 3108 9528
rect 2780 9036 2832 9042
rect 2780 8978 2832 8984
rect 2792 8945 2820 8978
rect 2778 8936 2834 8945
rect 2778 8871 2834 8880
rect 2780 8424 2832 8430
rect 2780 8366 2832 8372
rect 2792 7585 2820 8366
rect 2778 7576 2834 7585
rect 2778 7511 2834 7520
rect 2964 7200 3016 7206
rect 2964 7142 3016 7148
rect 2780 6860 2832 6866
rect 2780 6802 2832 6808
rect 2792 4865 2820 6802
rect 2976 6322 3004 7142
rect 3712 6914 3740 13874
rect 4172 11778 4200 33866
rect 4356 26234 4384 34954
rect 4423 34300 4731 34309
rect 4423 34298 4429 34300
rect 4485 34298 4509 34300
rect 4565 34298 4589 34300
rect 4645 34298 4669 34300
rect 4725 34298 4731 34300
rect 4485 34246 4487 34298
rect 4667 34246 4669 34298
rect 4423 34244 4429 34246
rect 4485 34244 4509 34246
rect 4565 34244 4589 34246
rect 4645 34244 4669 34246
rect 4725 34244 4731 34246
rect 4423 34235 4731 34244
rect 4423 33212 4731 33221
rect 4423 33210 4429 33212
rect 4485 33210 4509 33212
rect 4565 33210 4589 33212
rect 4645 33210 4669 33212
rect 4725 33210 4731 33212
rect 4485 33158 4487 33210
rect 4667 33158 4669 33210
rect 4423 33156 4429 33158
rect 4485 33156 4509 33158
rect 4565 33156 4589 33158
rect 4645 33156 4669 33158
rect 4725 33156 4731 33158
rect 4423 33147 4731 33156
rect 4423 32124 4731 32133
rect 4423 32122 4429 32124
rect 4485 32122 4509 32124
rect 4565 32122 4589 32124
rect 4645 32122 4669 32124
rect 4725 32122 4731 32124
rect 4485 32070 4487 32122
rect 4667 32070 4669 32122
rect 4423 32068 4429 32070
rect 4485 32068 4509 32070
rect 4565 32068 4589 32070
rect 4645 32068 4669 32070
rect 4725 32068 4731 32070
rect 4423 32059 4731 32068
rect 4423 31036 4731 31045
rect 4423 31034 4429 31036
rect 4485 31034 4509 31036
rect 4565 31034 4589 31036
rect 4645 31034 4669 31036
rect 4725 31034 4731 31036
rect 4485 30982 4487 31034
rect 4667 30982 4669 31034
rect 4423 30980 4429 30982
rect 4485 30980 4509 30982
rect 4565 30980 4589 30982
rect 4645 30980 4669 30982
rect 4725 30980 4731 30982
rect 4423 30971 4731 30980
rect 4423 29948 4731 29957
rect 4423 29946 4429 29948
rect 4485 29946 4509 29948
rect 4565 29946 4589 29948
rect 4645 29946 4669 29948
rect 4725 29946 4731 29948
rect 4485 29894 4487 29946
rect 4667 29894 4669 29946
rect 4423 29892 4429 29894
rect 4485 29892 4509 29894
rect 4565 29892 4589 29894
rect 4645 29892 4669 29894
rect 4725 29892 4731 29894
rect 4423 29883 4731 29892
rect 4816 29238 4844 35566
rect 4804 29232 4856 29238
rect 4804 29174 4856 29180
rect 4423 28860 4731 28869
rect 4423 28858 4429 28860
rect 4485 28858 4509 28860
rect 4565 28858 4589 28860
rect 4645 28858 4669 28860
rect 4725 28858 4731 28860
rect 4485 28806 4487 28858
rect 4667 28806 4669 28858
rect 4423 28804 4429 28806
rect 4485 28804 4509 28806
rect 4565 28804 4589 28806
rect 4645 28804 4669 28806
rect 4725 28804 4731 28806
rect 4423 28795 4731 28804
rect 4423 27772 4731 27781
rect 4423 27770 4429 27772
rect 4485 27770 4509 27772
rect 4565 27770 4589 27772
rect 4645 27770 4669 27772
rect 4725 27770 4731 27772
rect 4485 27718 4487 27770
rect 4667 27718 4669 27770
rect 4423 27716 4429 27718
rect 4485 27716 4509 27718
rect 4565 27716 4589 27718
rect 4645 27716 4669 27718
rect 4725 27716 4731 27718
rect 4423 27707 4731 27716
rect 5000 27606 5028 36314
rect 5092 33930 5120 43726
rect 5540 38344 5592 38350
rect 5540 38286 5592 38292
rect 5552 35894 5580 38286
rect 6012 36786 6040 46854
rect 6748 37126 6776 46854
rect 7024 46578 7052 46990
rect 7896 46812 8204 46821
rect 7896 46810 7902 46812
rect 7958 46810 7982 46812
rect 8038 46810 8062 46812
rect 8118 46810 8142 46812
rect 8198 46810 8204 46812
rect 7958 46758 7960 46810
rect 8140 46758 8142 46810
rect 7896 46756 7902 46758
rect 7958 46756 7982 46758
rect 8038 46756 8062 46758
rect 8118 46756 8142 46758
rect 8198 46756 8204 46758
rect 7896 46747 8204 46756
rect 7012 46572 7064 46578
rect 7012 46514 7064 46520
rect 8404 46510 8432 49200
rect 10336 47122 10364 49200
rect 10324 47116 10376 47122
rect 10324 47058 10376 47064
rect 9312 47048 9364 47054
rect 9312 46990 9364 46996
rect 9220 46980 9272 46986
rect 9220 46922 9272 46928
rect 7932 46504 7984 46510
rect 7932 46446 7984 46452
rect 8392 46504 8444 46510
rect 8392 46446 8444 46452
rect 7944 46170 7972 46446
rect 7932 46164 7984 46170
rect 7932 46106 7984 46112
rect 9232 45966 9260 46922
rect 7748 45960 7800 45966
rect 7748 45902 7800 45908
rect 9220 45960 9272 45966
rect 9220 45902 9272 45908
rect 6736 37120 6788 37126
rect 6736 37062 6788 37068
rect 6000 36780 6052 36786
rect 6000 36722 6052 36728
rect 5552 35866 5764 35894
rect 5736 35630 5764 35866
rect 5724 35624 5776 35630
rect 5724 35566 5776 35572
rect 5736 34542 5764 35566
rect 7760 34678 7788 45902
rect 7896 45724 8204 45733
rect 7896 45722 7902 45724
rect 7958 45722 7982 45724
rect 8038 45722 8062 45724
rect 8118 45722 8142 45724
rect 8198 45722 8204 45724
rect 7958 45670 7960 45722
rect 8140 45670 8142 45722
rect 7896 45668 7902 45670
rect 7958 45668 7982 45670
rect 8038 45668 8062 45670
rect 8118 45668 8142 45670
rect 8198 45668 8204 45670
rect 7896 45659 8204 45668
rect 9324 45490 9352 46990
rect 9496 46980 9548 46986
rect 9496 46922 9548 46928
rect 9508 46170 9536 46922
rect 10980 46510 11008 49200
rect 11624 47546 11652 49200
rect 11624 47518 11836 47546
rect 11369 47356 11677 47365
rect 11369 47354 11375 47356
rect 11431 47354 11455 47356
rect 11511 47354 11535 47356
rect 11591 47354 11615 47356
rect 11671 47354 11677 47356
rect 11431 47302 11433 47354
rect 11613 47302 11615 47354
rect 11369 47300 11375 47302
rect 11431 47300 11455 47302
rect 11511 47300 11535 47302
rect 11591 47300 11615 47302
rect 11671 47300 11677 47302
rect 11369 47291 11677 47300
rect 10140 46504 10192 46510
rect 10140 46446 10192 46452
rect 10968 46504 11020 46510
rect 10968 46446 11020 46452
rect 10152 46170 10180 46446
rect 10416 46436 10468 46442
rect 10416 46378 10468 46384
rect 9496 46164 9548 46170
rect 9496 46106 9548 46112
rect 10140 46164 10192 46170
rect 10140 46106 10192 46112
rect 10428 45490 10456 46378
rect 11704 46368 11756 46374
rect 11704 46310 11756 46316
rect 11369 46268 11677 46277
rect 11369 46266 11375 46268
rect 11431 46266 11455 46268
rect 11511 46266 11535 46268
rect 11591 46266 11615 46268
rect 11671 46266 11677 46268
rect 11431 46214 11433 46266
rect 11613 46214 11615 46266
rect 11369 46212 11375 46214
rect 11431 46212 11455 46214
rect 11511 46212 11535 46214
rect 11591 46212 11615 46214
rect 11671 46212 11677 46214
rect 11369 46203 11677 46212
rect 11716 46034 11744 46310
rect 11808 46034 11836 47518
rect 12900 47048 12952 47054
rect 12900 46990 12952 46996
rect 12912 46578 12940 46990
rect 12900 46572 12952 46578
rect 12900 46514 12952 46520
rect 13556 46510 13584 49200
rect 15120 47002 15148 49286
rect 15446 49200 15558 49800
rect 16090 49200 16202 49800
rect 16734 49200 16846 49800
rect 17378 49200 17490 49800
rect 18022 49200 18134 49800
rect 18666 49200 18778 49800
rect 19954 49200 20066 49800
rect 20598 49200 20710 49800
rect 21242 49200 21354 49800
rect 21886 49200 21998 49800
rect 22530 49200 22642 49800
rect 23174 49200 23286 49800
rect 23818 49314 23930 49800
rect 23818 49286 24072 49314
rect 23818 49200 23930 49286
rect 15120 46974 15240 47002
rect 14842 46812 15150 46821
rect 14842 46810 14848 46812
rect 14904 46810 14928 46812
rect 14984 46810 15008 46812
rect 15064 46810 15088 46812
rect 15144 46810 15150 46812
rect 14904 46758 14906 46810
rect 15086 46758 15088 46810
rect 14842 46756 14848 46758
rect 14904 46756 14928 46758
rect 14984 46756 15008 46758
rect 15064 46756 15088 46758
rect 15144 46756 15150 46758
rect 14842 46747 15150 46756
rect 13084 46504 13136 46510
rect 13084 46446 13136 46452
rect 13544 46504 13596 46510
rect 13544 46446 13596 46452
rect 11704 46028 11756 46034
rect 11704 45970 11756 45976
rect 11796 46028 11848 46034
rect 11796 45970 11848 45976
rect 10692 45960 10744 45966
rect 10692 45902 10744 45908
rect 9312 45484 9364 45490
rect 9312 45426 9364 45432
rect 10416 45484 10468 45490
rect 10416 45426 10468 45432
rect 7896 44636 8204 44645
rect 7896 44634 7902 44636
rect 7958 44634 7982 44636
rect 8038 44634 8062 44636
rect 8118 44634 8142 44636
rect 8198 44634 8204 44636
rect 7958 44582 7960 44634
rect 8140 44582 8142 44634
rect 7896 44580 7902 44582
rect 7958 44580 7982 44582
rect 8038 44580 8062 44582
rect 8118 44580 8142 44582
rect 8198 44580 8204 44582
rect 7896 44571 8204 44580
rect 10704 43790 10732 45902
rect 12716 45824 12768 45830
rect 12716 45766 12768 45772
rect 11369 45180 11677 45189
rect 11369 45178 11375 45180
rect 11431 45178 11455 45180
rect 11511 45178 11535 45180
rect 11591 45178 11615 45180
rect 11671 45178 11677 45180
rect 11431 45126 11433 45178
rect 11613 45126 11615 45178
rect 11369 45124 11375 45126
rect 11431 45124 11455 45126
rect 11511 45124 11535 45126
rect 11591 45124 11615 45126
rect 11671 45124 11677 45126
rect 11369 45115 11677 45124
rect 11369 44092 11677 44101
rect 11369 44090 11375 44092
rect 11431 44090 11455 44092
rect 11511 44090 11535 44092
rect 11591 44090 11615 44092
rect 11671 44090 11677 44092
rect 11431 44038 11433 44090
rect 11613 44038 11615 44090
rect 11369 44036 11375 44038
rect 11431 44036 11455 44038
rect 11511 44036 11535 44038
rect 11591 44036 11615 44038
rect 11671 44036 11677 44038
rect 11369 44027 11677 44036
rect 10692 43784 10744 43790
rect 10692 43726 10744 43732
rect 7896 43548 8204 43557
rect 7896 43546 7902 43548
rect 7958 43546 7982 43548
rect 8038 43546 8062 43548
rect 8118 43546 8142 43548
rect 8198 43546 8204 43548
rect 7958 43494 7960 43546
rect 8140 43494 8142 43546
rect 7896 43492 7902 43494
rect 7958 43492 7982 43494
rect 8038 43492 8062 43494
rect 8118 43492 8142 43494
rect 8198 43492 8204 43494
rect 7896 43483 8204 43492
rect 11369 43004 11677 43013
rect 11369 43002 11375 43004
rect 11431 43002 11455 43004
rect 11511 43002 11535 43004
rect 11591 43002 11615 43004
rect 11671 43002 11677 43004
rect 11431 42950 11433 43002
rect 11613 42950 11615 43002
rect 11369 42948 11375 42950
rect 11431 42948 11455 42950
rect 11511 42948 11535 42950
rect 11591 42948 11615 42950
rect 11671 42948 11677 42950
rect 11369 42939 11677 42948
rect 7896 42460 8204 42469
rect 7896 42458 7902 42460
rect 7958 42458 7982 42460
rect 8038 42458 8062 42460
rect 8118 42458 8142 42460
rect 8198 42458 8204 42460
rect 7958 42406 7960 42458
rect 8140 42406 8142 42458
rect 7896 42404 7902 42406
rect 7958 42404 7982 42406
rect 8038 42404 8062 42406
rect 8118 42404 8142 42406
rect 8198 42404 8204 42406
rect 7896 42395 8204 42404
rect 11369 41916 11677 41925
rect 11369 41914 11375 41916
rect 11431 41914 11455 41916
rect 11511 41914 11535 41916
rect 11591 41914 11615 41916
rect 11671 41914 11677 41916
rect 11431 41862 11433 41914
rect 11613 41862 11615 41914
rect 11369 41860 11375 41862
rect 11431 41860 11455 41862
rect 11511 41860 11535 41862
rect 11591 41860 11615 41862
rect 11671 41860 11677 41862
rect 11369 41851 11677 41860
rect 7896 41372 8204 41381
rect 7896 41370 7902 41372
rect 7958 41370 7982 41372
rect 8038 41370 8062 41372
rect 8118 41370 8142 41372
rect 8198 41370 8204 41372
rect 7958 41318 7960 41370
rect 8140 41318 8142 41370
rect 7896 41316 7902 41318
rect 7958 41316 7982 41318
rect 8038 41316 8062 41318
rect 8118 41316 8142 41318
rect 8198 41316 8204 41318
rect 7896 41307 8204 41316
rect 11369 40828 11677 40837
rect 11369 40826 11375 40828
rect 11431 40826 11455 40828
rect 11511 40826 11535 40828
rect 11591 40826 11615 40828
rect 11671 40826 11677 40828
rect 11431 40774 11433 40826
rect 11613 40774 11615 40826
rect 11369 40772 11375 40774
rect 11431 40772 11455 40774
rect 11511 40772 11535 40774
rect 11591 40772 11615 40774
rect 11671 40772 11677 40774
rect 11369 40763 11677 40772
rect 7896 40284 8204 40293
rect 7896 40282 7902 40284
rect 7958 40282 7982 40284
rect 8038 40282 8062 40284
rect 8118 40282 8142 40284
rect 8198 40282 8204 40284
rect 7958 40230 7960 40282
rect 8140 40230 8142 40282
rect 7896 40228 7902 40230
rect 7958 40228 7982 40230
rect 8038 40228 8062 40230
rect 8118 40228 8142 40230
rect 8198 40228 8204 40230
rect 7896 40219 8204 40228
rect 11369 39740 11677 39749
rect 11369 39738 11375 39740
rect 11431 39738 11455 39740
rect 11511 39738 11535 39740
rect 11591 39738 11615 39740
rect 11671 39738 11677 39740
rect 11431 39686 11433 39738
rect 11613 39686 11615 39738
rect 11369 39684 11375 39686
rect 11431 39684 11455 39686
rect 11511 39684 11535 39686
rect 11591 39684 11615 39686
rect 11671 39684 11677 39686
rect 11369 39675 11677 39684
rect 7896 39196 8204 39205
rect 7896 39194 7902 39196
rect 7958 39194 7982 39196
rect 8038 39194 8062 39196
rect 8118 39194 8142 39196
rect 8198 39194 8204 39196
rect 7958 39142 7960 39194
rect 8140 39142 8142 39194
rect 7896 39140 7902 39142
rect 7958 39140 7982 39142
rect 8038 39140 8062 39142
rect 8118 39140 8142 39142
rect 8198 39140 8204 39142
rect 7896 39131 8204 39140
rect 11369 38652 11677 38661
rect 11369 38650 11375 38652
rect 11431 38650 11455 38652
rect 11511 38650 11535 38652
rect 11591 38650 11615 38652
rect 11671 38650 11677 38652
rect 11431 38598 11433 38650
rect 11613 38598 11615 38650
rect 11369 38596 11375 38598
rect 11431 38596 11455 38598
rect 11511 38596 11535 38598
rect 11591 38596 11615 38598
rect 11671 38596 11677 38598
rect 11369 38587 11677 38596
rect 7896 38108 8204 38117
rect 7896 38106 7902 38108
rect 7958 38106 7982 38108
rect 8038 38106 8062 38108
rect 8118 38106 8142 38108
rect 8198 38106 8204 38108
rect 7958 38054 7960 38106
rect 8140 38054 8142 38106
rect 7896 38052 7902 38054
rect 7958 38052 7982 38054
rect 8038 38052 8062 38054
rect 8118 38052 8142 38054
rect 8198 38052 8204 38054
rect 7896 38043 8204 38052
rect 11369 37564 11677 37573
rect 11369 37562 11375 37564
rect 11431 37562 11455 37564
rect 11511 37562 11535 37564
rect 11591 37562 11615 37564
rect 11671 37562 11677 37564
rect 11431 37510 11433 37562
rect 11613 37510 11615 37562
rect 11369 37508 11375 37510
rect 11431 37508 11455 37510
rect 11511 37508 11535 37510
rect 11591 37508 11615 37510
rect 11671 37508 11677 37510
rect 11369 37499 11677 37508
rect 7896 37020 8204 37029
rect 7896 37018 7902 37020
rect 7958 37018 7982 37020
rect 8038 37018 8062 37020
rect 8118 37018 8142 37020
rect 8198 37018 8204 37020
rect 7958 36966 7960 37018
rect 8140 36966 8142 37018
rect 7896 36964 7902 36966
rect 7958 36964 7982 36966
rect 8038 36964 8062 36966
rect 8118 36964 8142 36966
rect 8198 36964 8204 36966
rect 7896 36955 8204 36964
rect 11369 36476 11677 36485
rect 11369 36474 11375 36476
rect 11431 36474 11455 36476
rect 11511 36474 11535 36476
rect 11591 36474 11615 36476
rect 11671 36474 11677 36476
rect 11431 36422 11433 36474
rect 11613 36422 11615 36474
rect 11369 36420 11375 36422
rect 11431 36420 11455 36422
rect 11511 36420 11535 36422
rect 11591 36420 11615 36422
rect 11671 36420 11677 36422
rect 11369 36411 11677 36420
rect 12072 36100 12124 36106
rect 12072 36042 12124 36048
rect 7896 35932 8204 35941
rect 7896 35930 7902 35932
rect 7958 35930 7982 35932
rect 8038 35930 8062 35932
rect 8118 35930 8142 35932
rect 8198 35930 8204 35932
rect 7958 35878 7960 35930
rect 8140 35878 8142 35930
rect 7896 35876 7902 35878
rect 7958 35876 7982 35878
rect 8038 35876 8062 35878
rect 8118 35876 8142 35878
rect 8198 35876 8204 35878
rect 7896 35867 8204 35876
rect 12084 35834 12112 36042
rect 12072 35828 12124 35834
rect 12072 35770 12124 35776
rect 12728 35766 12756 45766
rect 13096 45626 13124 46446
rect 14188 45960 14240 45966
rect 14188 45902 14240 45908
rect 13268 45824 13320 45830
rect 13268 45766 13320 45772
rect 13084 45620 13136 45626
rect 13084 45562 13136 45568
rect 13280 45490 13308 45766
rect 14200 45490 14228 45902
rect 14842 45724 15150 45733
rect 14842 45722 14848 45724
rect 14904 45722 14928 45724
rect 14984 45722 15008 45724
rect 15064 45722 15088 45724
rect 15144 45722 15150 45724
rect 14904 45670 14906 45722
rect 15086 45670 15088 45722
rect 14842 45668 14848 45670
rect 14904 45668 14928 45670
rect 14984 45668 15008 45670
rect 15064 45668 15088 45670
rect 15144 45668 15150 45670
rect 14842 45659 15150 45668
rect 13268 45484 13320 45490
rect 13268 45426 13320 45432
rect 14188 45484 14240 45490
rect 14188 45426 14240 45432
rect 15212 45422 15240 46974
rect 15844 46572 15896 46578
rect 15844 46514 15896 46520
rect 15856 45830 15884 46514
rect 15936 46504 15988 46510
rect 15936 46446 15988 46452
rect 15948 46034 15976 46446
rect 16120 46368 16172 46374
rect 16120 46310 16172 46316
rect 16132 46034 16160 46310
rect 16776 46034 16804 49200
rect 18315 47356 18623 47365
rect 18315 47354 18321 47356
rect 18377 47354 18401 47356
rect 18457 47354 18481 47356
rect 18537 47354 18561 47356
rect 18617 47354 18623 47356
rect 18377 47302 18379 47354
rect 18559 47302 18561 47354
rect 18315 47300 18321 47302
rect 18377 47300 18401 47302
rect 18457 47300 18481 47302
rect 18537 47300 18561 47302
rect 18617 47300 18623 47302
rect 18315 47291 18623 47300
rect 18236 47048 18288 47054
rect 18236 46990 18288 46996
rect 18248 46578 18276 46990
rect 18236 46572 18288 46578
rect 18236 46514 18288 46520
rect 18708 46510 18736 49200
rect 19996 46918 20024 49200
rect 19984 46912 20036 46918
rect 19984 46854 20036 46860
rect 18144 46504 18196 46510
rect 18144 46446 18196 46452
rect 18696 46504 18748 46510
rect 18696 46446 18748 46452
rect 17224 46436 17276 46442
rect 17224 46378 17276 46384
rect 17236 46170 17264 46378
rect 18156 46170 18184 46446
rect 20260 46368 20312 46374
rect 20260 46310 20312 46316
rect 18315 46268 18623 46277
rect 18315 46266 18321 46268
rect 18377 46266 18401 46268
rect 18457 46266 18481 46268
rect 18537 46266 18561 46268
rect 18617 46266 18623 46268
rect 18377 46214 18379 46266
rect 18559 46214 18561 46266
rect 18315 46212 18321 46214
rect 18377 46212 18401 46214
rect 18457 46212 18481 46214
rect 18537 46212 18561 46214
rect 18617 46212 18623 46214
rect 18315 46203 18623 46212
rect 17224 46164 17276 46170
rect 17224 46106 17276 46112
rect 18144 46164 18196 46170
rect 18144 46106 18196 46112
rect 20272 46034 20300 46310
rect 21284 46034 21312 49200
rect 21788 46812 22096 46821
rect 21788 46810 21794 46812
rect 21850 46810 21874 46812
rect 21930 46810 21954 46812
rect 22010 46810 22034 46812
rect 22090 46810 22096 46812
rect 21850 46758 21852 46810
rect 22032 46758 22034 46810
rect 21788 46756 21794 46758
rect 21850 46756 21874 46758
rect 21930 46756 21954 46758
rect 22010 46756 22034 46758
rect 22090 46756 22096 46758
rect 21788 46747 22096 46756
rect 15936 46028 15988 46034
rect 15936 45970 15988 45976
rect 16120 46028 16172 46034
rect 16120 45970 16172 45976
rect 16764 46028 16816 46034
rect 16764 45970 16816 45976
rect 20260 46028 20312 46034
rect 20260 45970 20312 45976
rect 21272 46028 21324 46034
rect 21272 45970 21324 45976
rect 18328 45960 18380 45966
rect 18328 45902 18380 45908
rect 15844 45824 15896 45830
rect 15844 45766 15896 45772
rect 14372 45416 14424 45422
rect 14372 45358 14424 45364
rect 15200 45416 15252 45422
rect 15200 45358 15252 45364
rect 14384 44538 14412 45358
rect 14842 44636 15150 44645
rect 14842 44634 14848 44636
rect 14904 44634 14928 44636
rect 14984 44634 15008 44636
rect 15064 44634 15088 44636
rect 15144 44634 15150 44636
rect 14904 44582 14906 44634
rect 15086 44582 15088 44634
rect 14842 44580 14848 44582
rect 14904 44580 14928 44582
rect 14984 44580 15008 44582
rect 15064 44580 15088 44582
rect 15144 44580 15150 44582
rect 14842 44571 15150 44580
rect 14372 44532 14424 44538
rect 14372 44474 14424 44480
rect 14372 44396 14424 44402
rect 14372 44338 14424 44344
rect 12716 35760 12768 35766
rect 12716 35702 12768 35708
rect 11369 35388 11677 35397
rect 11369 35386 11375 35388
rect 11431 35386 11455 35388
rect 11511 35386 11535 35388
rect 11591 35386 11615 35388
rect 11671 35386 11677 35388
rect 11431 35334 11433 35386
rect 11613 35334 11615 35386
rect 11369 35332 11375 35334
rect 11431 35332 11455 35334
rect 11511 35332 11535 35334
rect 11591 35332 11615 35334
rect 11671 35332 11677 35334
rect 11369 35323 11677 35332
rect 12728 35290 12756 35702
rect 12716 35284 12768 35290
rect 12716 35226 12768 35232
rect 7896 34844 8204 34853
rect 7896 34842 7902 34844
rect 7958 34842 7982 34844
rect 8038 34842 8062 34844
rect 8118 34842 8142 34844
rect 8198 34842 8204 34844
rect 7958 34790 7960 34842
rect 8140 34790 8142 34842
rect 7896 34788 7902 34790
rect 7958 34788 7982 34790
rect 8038 34788 8062 34790
rect 8118 34788 8142 34790
rect 8198 34788 8204 34790
rect 7896 34779 8204 34788
rect 7748 34672 7800 34678
rect 7748 34614 7800 34620
rect 5172 34536 5224 34542
rect 5172 34478 5224 34484
rect 5724 34536 5776 34542
rect 5724 34478 5776 34484
rect 8392 34536 8444 34542
rect 8392 34478 8444 34484
rect 5080 33924 5132 33930
rect 5080 33866 5132 33872
rect 4988 27600 5040 27606
rect 4988 27542 5040 27548
rect 4423 26684 4731 26693
rect 4423 26682 4429 26684
rect 4485 26682 4509 26684
rect 4565 26682 4589 26684
rect 4645 26682 4669 26684
rect 4725 26682 4731 26684
rect 4485 26630 4487 26682
rect 4667 26630 4669 26682
rect 4423 26628 4429 26630
rect 4485 26628 4509 26630
rect 4565 26628 4589 26630
rect 4645 26628 4669 26630
rect 4725 26628 4731 26630
rect 4423 26619 4731 26628
rect 4264 26206 4384 26234
rect 4264 16574 4292 26206
rect 4423 25596 4731 25605
rect 4423 25594 4429 25596
rect 4485 25594 4509 25596
rect 4565 25594 4589 25596
rect 4645 25594 4669 25596
rect 4725 25594 4731 25596
rect 4485 25542 4487 25594
rect 4667 25542 4669 25594
rect 4423 25540 4429 25542
rect 4485 25540 4509 25542
rect 4565 25540 4589 25542
rect 4645 25540 4669 25542
rect 4725 25540 4731 25542
rect 4423 25531 4731 25540
rect 4423 24508 4731 24517
rect 4423 24506 4429 24508
rect 4485 24506 4509 24508
rect 4565 24506 4589 24508
rect 4645 24506 4669 24508
rect 4725 24506 4731 24508
rect 4485 24454 4487 24506
rect 4667 24454 4669 24506
rect 4423 24452 4429 24454
rect 4485 24452 4509 24454
rect 4565 24452 4589 24454
rect 4645 24452 4669 24454
rect 4725 24452 4731 24454
rect 4423 24443 4731 24452
rect 4423 23420 4731 23429
rect 4423 23418 4429 23420
rect 4485 23418 4509 23420
rect 4565 23418 4589 23420
rect 4645 23418 4669 23420
rect 4725 23418 4731 23420
rect 4485 23366 4487 23418
rect 4667 23366 4669 23418
rect 4423 23364 4429 23366
rect 4485 23364 4509 23366
rect 4565 23364 4589 23366
rect 4645 23364 4669 23366
rect 4725 23364 4731 23366
rect 4423 23355 4731 23364
rect 4423 22332 4731 22341
rect 4423 22330 4429 22332
rect 4485 22330 4509 22332
rect 4565 22330 4589 22332
rect 4645 22330 4669 22332
rect 4725 22330 4731 22332
rect 4485 22278 4487 22330
rect 4667 22278 4669 22330
rect 4423 22276 4429 22278
rect 4485 22276 4509 22278
rect 4565 22276 4589 22278
rect 4645 22276 4669 22278
rect 4725 22276 4731 22278
rect 4423 22267 4731 22276
rect 4423 21244 4731 21253
rect 4423 21242 4429 21244
rect 4485 21242 4509 21244
rect 4565 21242 4589 21244
rect 4645 21242 4669 21244
rect 4725 21242 4731 21244
rect 4485 21190 4487 21242
rect 4667 21190 4669 21242
rect 4423 21188 4429 21190
rect 4485 21188 4509 21190
rect 4565 21188 4589 21190
rect 4645 21188 4669 21190
rect 4725 21188 4731 21190
rect 4423 21179 4731 21188
rect 4423 20156 4731 20165
rect 4423 20154 4429 20156
rect 4485 20154 4509 20156
rect 4565 20154 4589 20156
rect 4645 20154 4669 20156
rect 4725 20154 4731 20156
rect 4485 20102 4487 20154
rect 4667 20102 4669 20154
rect 4423 20100 4429 20102
rect 4485 20100 4509 20102
rect 4565 20100 4589 20102
rect 4645 20100 4669 20102
rect 4725 20100 4731 20102
rect 4423 20091 4731 20100
rect 4423 19068 4731 19077
rect 4423 19066 4429 19068
rect 4485 19066 4509 19068
rect 4565 19066 4589 19068
rect 4645 19066 4669 19068
rect 4725 19066 4731 19068
rect 4485 19014 4487 19066
rect 4667 19014 4669 19066
rect 4423 19012 4429 19014
rect 4485 19012 4509 19014
rect 4565 19012 4589 19014
rect 4645 19012 4669 19014
rect 4725 19012 4731 19014
rect 4423 19003 4731 19012
rect 4423 17980 4731 17989
rect 4423 17978 4429 17980
rect 4485 17978 4509 17980
rect 4565 17978 4589 17980
rect 4645 17978 4669 17980
rect 4725 17978 4731 17980
rect 4485 17926 4487 17978
rect 4667 17926 4669 17978
rect 4423 17924 4429 17926
rect 4485 17924 4509 17926
rect 4565 17924 4589 17926
rect 4645 17924 4669 17926
rect 4725 17924 4731 17926
rect 4423 17915 4731 17924
rect 5184 17882 5212 34478
rect 7896 33756 8204 33765
rect 7896 33754 7902 33756
rect 7958 33754 7982 33756
rect 8038 33754 8062 33756
rect 8118 33754 8142 33756
rect 8198 33754 8204 33756
rect 7958 33702 7960 33754
rect 8140 33702 8142 33754
rect 7896 33700 7902 33702
rect 7958 33700 7982 33702
rect 8038 33700 8062 33702
rect 8118 33700 8142 33702
rect 8198 33700 8204 33702
rect 7896 33691 8204 33700
rect 7896 32668 8204 32677
rect 7896 32666 7902 32668
rect 7958 32666 7982 32668
rect 8038 32666 8062 32668
rect 8118 32666 8142 32668
rect 8198 32666 8204 32668
rect 7958 32614 7960 32666
rect 8140 32614 8142 32666
rect 7896 32612 7902 32614
rect 7958 32612 7982 32614
rect 8038 32612 8062 32614
rect 8118 32612 8142 32614
rect 8198 32612 8204 32614
rect 7896 32603 8204 32612
rect 7896 31580 8204 31589
rect 7896 31578 7902 31580
rect 7958 31578 7982 31580
rect 8038 31578 8062 31580
rect 8118 31578 8142 31580
rect 8198 31578 8204 31580
rect 7958 31526 7960 31578
rect 8140 31526 8142 31578
rect 7896 31524 7902 31526
rect 7958 31524 7982 31526
rect 8038 31524 8062 31526
rect 8118 31524 8142 31526
rect 8198 31524 8204 31526
rect 7896 31515 8204 31524
rect 7896 30492 8204 30501
rect 7896 30490 7902 30492
rect 7958 30490 7982 30492
rect 8038 30490 8062 30492
rect 8118 30490 8142 30492
rect 8198 30490 8204 30492
rect 7958 30438 7960 30490
rect 8140 30438 8142 30490
rect 7896 30436 7902 30438
rect 7958 30436 7982 30438
rect 8038 30436 8062 30438
rect 8118 30436 8142 30438
rect 8198 30436 8204 30438
rect 7896 30427 8204 30436
rect 7896 29404 8204 29413
rect 7896 29402 7902 29404
rect 7958 29402 7982 29404
rect 8038 29402 8062 29404
rect 8118 29402 8142 29404
rect 8198 29402 8204 29404
rect 7958 29350 7960 29402
rect 8140 29350 8142 29402
rect 7896 29348 7902 29350
rect 7958 29348 7982 29350
rect 8038 29348 8062 29350
rect 8118 29348 8142 29350
rect 8198 29348 8204 29350
rect 7896 29339 8204 29348
rect 7896 28316 8204 28325
rect 7896 28314 7902 28316
rect 7958 28314 7982 28316
rect 8038 28314 8062 28316
rect 8118 28314 8142 28316
rect 8198 28314 8204 28316
rect 7958 28262 7960 28314
rect 8140 28262 8142 28314
rect 7896 28260 7902 28262
rect 7958 28260 7982 28262
rect 8038 28260 8062 28262
rect 8118 28260 8142 28262
rect 8198 28260 8204 28262
rect 7896 28251 8204 28260
rect 7896 27228 8204 27237
rect 7896 27226 7902 27228
rect 7958 27226 7982 27228
rect 8038 27226 8062 27228
rect 8118 27226 8142 27228
rect 8198 27226 8204 27228
rect 7958 27174 7960 27226
rect 8140 27174 8142 27226
rect 7896 27172 7902 27174
rect 7958 27172 7982 27174
rect 8038 27172 8062 27174
rect 8118 27172 8142 27174
rect 8198 27172 8204 27174
rect 7896 27163 8204 27172
rect 7896 26140 8204 26149
rect 7896 26138 7902 26140
rect 7958 26138 7982 26140
rect 8038 26138 8062 26140
rect 8118 26138 8142 26140
rect 8198 26138 8204 26140
rect 7958 26086 7960 26138
rect 8140 26086 8142 26138
rect 7896 26084 7902 26086
rect 7958 26084 7982 26086
rect 8038 26084 8062 26086
rect 8118 26084 8142 26086
rect 8198 26084 8204 26086
rect 7896 26075 8204 26084
rect 7896 25052 8204 25061
rect 7896 25050 7902 25052
rect 7958 25050 7982 25052
rect 8038 25050 8062 25052
rect 8118 25050 8142 25052
rect 8198 25050 8204 25052
rect 7958 24998 7960 25050
rect 8140 24998 8142 25050
rect 7896 24996 7902 24998
rect 7958 24996 7982 24998
rect 8038 24996 8062 24998
rect 8118 24996 8142 24998
rect 8198 24996 8204 24998
rect 7896 24987 8204 24996
rect 7896 23964 8204 23973
rect 7896 23962 7902 23964
rect 7958 23962 7982 23964
rect 8038 23962 8062 23964
rect 8118 23962 8142 23964
rect 8198 23962 8204 23964
rect 7958 23910 7960 23962
rect 8140 23910 8142 23962
rect 7896 23908 7902 23910
rect 7958 23908 7982 23910
rect 8038 23908 8062 23910
rect 8118 23908 8142 23910
rect 8198 23908 8204 23910
rect 7896 23899 8204 23908
rect 7896 22876 8204 22885
rect 7896 22874 7902 22876
rect 7958 22874 7982 22876
rect 8038 22874 8062 22876
rect 8118 22874 8142 22876
rect 8198 22874 8204 22876
rect 7958 22822 7960 22874
rect 8140 22822 8142 22874
rect 7896 22820 7902 22822
rect 7958 22820 7982 22822
rect 8038 22820 8062 22822
rect 8118 22820 8142 22822
rect 8198 22820 8204 22822
rect 7896 22811 8204 22820
rect 7896 21788 8204 21797
rect 7896 21786 7902 21788
rect 7958 21786 7982 21788
rect 8038 21786 8062 21788
rect 8118 21786 8142 21788
rect 8198 21786 8204 21788
rect 7958 21734 7960 21786
rect 8140 21734 8142 21786
rect 7896 21732 7902 21734
rect 7958 21732 7982 21734
rect 8038 21732 8062 21734
rect 8118 21732 8142 21734
rect 8198 21732 8204 21734
rect 7896 21723 8204 21732
rect 7896 20700 8204 20709
rect 7896 20698 7902 20700
rect 7958 20698 7982 20700
rect 8038 20698 8062 20700
rect 8118 20698 8142 20700
rect 8198 20698 8204 20700
rect 7958 20646 7960 20698
rect 8140 20646 8142 20698
rect 7896 20644 7902 20646
rect 7958 20644 7982 20646
rect 8038 20644 8062 20646
rect 8118 20644 8142 20646
rect 8198 20644 8204 20646
rect 7896 20635 8204 20644
rect 7896 19612 8204 19621
rect 7896 19610 7902 19612
rect 7958 19610 7982 19612
rect 8038 19610 8062 19612
rect 8118 19610 8142 19612
rect 8198 19610 8204 19612
rect 7958 19558 7960 19610
rect 8140 19558 8142 19610
rect 7896 19556 7902 19558
rect 7958 19556 7982 19558
rect 8038 19556 8062 19558
rect 8118 19556 8142 19558
rect 8198 19556 8204 19558
rect 7896 19547 8204 19556
rect 7896 18524 8204 18533
rect 7896 18522 7902 18524
rect 7958 18522 7982 18524
rect 8038 18522 8062 18524
rect 8118 18522 8142 18524
rect 8198 18522 8204 18524
rect 7958 18470 7960 18522
rect 8140 18470 8142 18522
rect 7896 18468 7902 18470
rect 7958 18468 7982 18470
rect 8038 18468 8062 18470
rect 8118 18468 8142 18470
rect 8198 18468 8204 18470
rect 7896 18459 8204 18468
rect 5172 17876 5224 17882
rect 5172 17818 5224 17824
rect 7896 17436 8204 17445
rect 7896 17434 7902 17436
rect 7958 17434 7982 17436
rect 8038 17434 8062 17436
rect 8118 17434 8142 17436
rect 8198 17434 8204 17436
rect 7958 17382 7960 17434
rect 8140 17382 8142 17434
rect 7896 17380 7902 17382
rect 7958 17380 7982 17382
rect 8038 17380 8062 17382
rect 8118 17380 8142 17382
rect 8198 17380 8204 17382
rect 7896 17371 8204 17380
rect 4423 16892 4731 16901
rect 4423 16890 4429 16892
rect 4485 16890 4509 16892
rect 4565 16890 4589 16892
rect 4645 16890 4669 16892
rect 4725 16890 4731 16892
rect 4485 16838 4487 16890
rect 4667 16838 4669 16890
rect 4423 16836 4429 16838
rect 4485 16836 4509 16838
rect 4565 16836 4589 16838
rect 4645 16836 4669 16838
rect 4725 16836 4731 16838
rect 4423 16827 4731 16836
rect 4264 16546 4384 16574
rect 4172 11750 4292 11778
rect 4068 9512 4120 9518
rect 4068 9454 4120 9460
rect 4160 9512 4212 9518
rect 4160 9454 4212 9460
rect 4080 9178 4108 9454
rect 4068 9172 4120 9178
rect 4068 9114 4120 9120
rect 4172 8378 4200 9454
rect 4080 8350 4200 8378
rect 3976 8288 4028 8294
rect 4080 8265 4108 8350
rect 4160 8288 4212 8294
rect 3976 8230 4028 8236
rect 4066 8256 4122 8265
rect 3988 7954 4016 8230
rect 4160 8230 4212 8236
rect 4066 8191 4122 8200
rect 4172 7954 4200 8230
rect 3976 7948 4028 7954
rect 3976 7890 4028 7896
rect 4160 7948 4212 7954
rect 4160 7890 4212 7896
rect 3620 6886 3740 6914
rect 4264 6914 4292 11750
rect 4356 8974 4384 16546
rect 7896 16348 8204 16357
rect 7896 16346 7902 16348
rect 7958 16346 7982 16348
rect 8038 16346 8062 16348
rect 8118 16346 8142 16348
rect 8198 16346 8204 16348
rect 7958 16294 7960 16346
rect 8140 16294 8142 16346
rect 7896 16292 7902 16294
rect 7958 16292 7982 16294
rect 8038 16292 8062 16294
rect 8118 16292 8142 16294
rect 8198 16292 8204 16294
rect 7896 16283 8204 16292
rect 4423 15804 4731 15813
rect 4423 15802 4429 15804
rect 4485 15802 4509 15804
rect 4565 15802 4589 15804
rect 4645 15802 4669 15804
rect 4725 15802 4731 15804
rect 4485 15750 4487 15802
rect 4667 15750 4669 15802
rect 4423 15748 4429 15750
rect 4485 15748 4509 15750
rect 4565 15748 4589 15750
rect 4645 15748 4669 15750
rect 4725 15748 4731 15750
rect 4423 15739 4731 15748
rect 7896 15260 8204 15269
rect 7896 15258 7902 15260
rect 7958 15258 7982 15260
rect 8038 15258 8062 15260
rect 8118 15258 8142 15260
rect 8198 15258 8204 15260
rect 7958 15206 7960 15258
rect 8140 15206 8142 15258
rect 7896 15204 7902 15206
rect 7958 15204 7982 15206
rect 8038 15204 8062 15206
rect 8118 15204 8142 15206
rect 8198 15204 8204 15206
rect 7896 15195 8204 15204
rect 4423 14716 4731 14725
rect 4423 14714 4429 14716
rect 4485 14714 4509 14716
rect 4565 14714 4589 14716
rect 4645 14714 4669 14716
rect 4725 14714 4731 14716
rect 4485 14662 4487 14714
rect 4667 14662 4669 14714
rect 4423 14660 4429 14662
rect 4485 14660 4509 14662
rect 4565 14660 4589 14662
rect 4645 14660 4669 14662
rect 4725 14660 4731 14662
rect 4423 14651 4731 14660
rect 8404 14414 8432 34478
rect 11369 34300 11677 34309
rect 11369 34298 11375 34300
rect 11431 34298 11455 34300
rect 11511 34298 11535 34300
rect 11591 34298 11615 34300
rect 11671 34298 11677 34300
rect 11431 34246 11433 34298
rect 11613 34246 11615 34298
rect 11369 34244 11375 34246
rect 11431 34244 11455 34246
rect 11511 34244 11535 34246
rect 11591 34244 11615 34246
rect 11671 34244 11677 34246
rect 11369 34235 11677 34244
rect 11369 33212 11677 33221
rect 11369 33210 11375 33212
rect 11431 33210 11455 33212
rect 11511 33210 11535 33212
rect 11591 33210 11615 33212
rect 11671 33210 11677 33212
rect 11431 33158 11433 33210
rect 11613 33158 11615 33210
rect 11369 33156 11375 33158
rect 11431 33156 11455 33158
rect 11511 33156 11535 33158
rect 11591 33156 11615 33158
rect 11671 33156 11677 33158
rect 11369 33147 11677 33156
rect 11369 32124 11677 32133
rect 11369 32122 11375 32124
rect 11431 32122 11455 32124
rect 11511 32122 11535 32124
rect 11591 32122 11615 32124
rect 11671 32122 11677 32124
rect 11431 32070 11433 32122
rect 11613 32070 11615 32122
rect 11369 32068 11375 32070
rect 11431 32068 11455 32070
rect 11511 32068 11535 32070
rect 11591 32068 11615 32070
rect 11671 32068 11677 32070
rect 11369 32059 11677 32068
rect 11369 31036 11677 31045
rect 11369 31034 11375 31036
rect 11431 31034 11455 31036
rect 11511 31034 11535 31036
rect 11591 31034 11615 31036
rect 11671 31034 11677 31036
rect 11431 30982 11433 31034
rect 11613 30982 11615 31034
rect 11369 30980 11375 30982
rect 11431 30980 11455 30982
rect 11511 30980 11535 30982
rect 11591 30980 11615 30982
rect 11671 30980 11677 30982
rect 11369 30971 11677 30980
rect 11369 29948 11677 29957
rect 11369 29946 11375 29948
rect 11431 29946 11455 29948
rect 11511 29946 11535 29948
rect 11591 29946 11615 29948
rect 11671 29946 11677 29948
rect 11431 29894 11433 29946
rect 11613 29894 11615 29946
rect 11369 29892 11375 29894
rect 11431 29892 11455 29894
rect 11511 29892 11535 29894
rect 11591 29892 11615 29894
rect 11671 29892 11677 29894
rect 11369 29883 11677 29892
rect 11369 28860 11677 28869
rect 11369 28858 11375 28860
rect 11431 28858 11455 28860
rect 11511 28858 11535 28860
rect 11591 28858 11615 28860
rect 11671 28858 11677 28860
rect 11431 28806 11433 28858
rect 11613 28806 11615 28858
rect 11369 28804 11375 28806
rect 11431 28804 11455 28806
rect 11511 28804 11535 28806
rect 11591 28804 11615 28806
rect 11671 28804 11677 28806
rect 11369 28795 11677 28804
rect 11369 27772 11677 27781
rect 11369 27770 11375 27772
rect 11431 27770 11455 27772
rect 11511 27770 11535 27772
rect 11591 27770 11615 27772
rect 11671 27770 11677 27772
rect 11431 27718 11433 27770
rect 11613 27718 11615 27770
rect 11369 27716 11375 27718
rect 11431 27716 11455 27718
rect 11511 27716 11535 27718
rect 11591 27716 11615 27718
rect 11671 27716 11677 27718
rect 11369 27707 11677 27716
rect 11369 26684 11677 26693
rect 11369 26682 11375 26684
rect 11431 26682 11455 26684
rect 11511 26682 11535 26684
rect 11591 26682 11615 26684
rect 11671 26682 11677 26684
rect 11431 26630 11433 26682
rect 11613 26630 11615 26682
rect 11369 26628 11375 26630
rect 11431 26628 11455 26630
rect 11511 26628 11535 26630
rect 11591 26628 11615 26630
rect 11671 26628 11677 26630
rect 11369 26619 11677 26628
rect 11369 25596 11677 25605
rect 11369 25594 11375 25596
rect 11431 25594 11455 25596
rect 11511 25594 11535 25596
rect 11591 25594 11615 25596
rect 11671 25594 11677 25596
rect 11431 25542 11433 25594
rect 11613 25542 11615 25594
rect 11369 25540 11375 25542
rect 11431 25540 11455 25542
rect 11511 25540 11535 25542
rect 11591 25540 11615 25542
rect 11671 25540 11677 25542
rect 11369 25531 11677 25540
rect 9496 25152 9548 25158
rect 9496 25094 9548 25100
rect 8392 14408 8444 14414
rect 8392 14350 8444 14356
rect 7896 14172 8204 14181
rect 7896 14170 7902 14172
rect 7958 14170 7982 14172
rect 8038 14170 8062 14172
rect 8118 14170 8142 14172
rect 8198 14170 8204 14172
rect 7958 14118 7960 14170
rect 8140 14118 8142 14170
rect 7896 14116 7902 14118
rect 7958 14116 7982 14118
rect 8038 14116 8062 14118
rect 8118 14116 8142 14118
rect 8198 14116 8204 14118
rect 7896 14107 8204 14116
rect 8300 13864 8352 13870
rect 8300 13806 8352 13812
rect 4423 13628 4731 13637
rect 4423 13626 4429 13628
rect 4485 13626 4509 13628
rect 4565 13626 4589 13628
rect 4645 13626 4669 13628
rect 4725 13626 4731 13628
rect 4485 13574 4487 13626
rect 4667 13574 4669 13626
rect 4423 13572 4429 13574
rect 4485 13572 4509 13574
rect 4565 13572 4589 13574
rect 4645 13572 4669 13574
rect 4725 13572 4731 13574
rect 4423 13563 4731 13572
rect 7896 13084 8204 13093
rect 7896 13082 7902 13084
rect 7958 13082 7982 13084
rect 8038 13082 8062 13084
rect 8118 13082 8142 13084
rect 8198 13082 8204 13084
rect 7958 13030 7960 13082
rect 8140 13030 8142 13082
rect 7896 13028 7902 13030
rect 7958 13028 7982 13030
rect 8038 13028 8062 13030
rect 8118 13028 8142 13030
rect 8198 13028 8204 13030
rect 7896 13019 8204 13028
rect 4423 12540 4731 12549
rect 4423 12538 4429 12540
rect 4485 12538 4509 12540
rect 4565 12538 4589 12540
rect 4645 12538 4669 12540
rect 4725 12538 4731 12540
rect 4485 12486 4487 12538
rect 4667 12486 4669 12538
rect 4423 12484 4429 12486
rect 4485 12484 4509 12486
rect 4565 12484 4589 12486
rect 4645 12484 4669 12486
rect 4725 12484 4731 12486
rect 4423 12475 4731 12484
rect 7896 11996 8204 12005
rect 7896 11994 7902 11996
rect 7958 11994 7982 11996
rect 8038 11994 8062 11996
rect 8118 11994 8142 11996
rect 8198 11994 8204 11996
rect 7958 11942 7960 11994
rect 8140 11942 8142 11994
rect 7896 11940 7902 11942
rect 7958 11940 7982 11942
rect 8038 11940 8062 11942
rect 8118 11940 8142 11942
rect 8198 11940 8204 11942
rect 7896 11931 8204 11940
rect 4423 11452 4731 11461
rect 4423 11450 4429 11452
rect 4485 11450 4509 11452
rect 4565 11450 4589 11452
rect 4645 11450 4669 11452
rect 4725 11450 4731 11452
rect 4485 11398 4487 11450
rect 4667 11398 4669 11450
rect 4423 11396 4429 11398
rect 4485 11396 4509 11398
rect 4565 11396 4589 11398
rect 4645 11396 4669 11398
rect 4725 11396 4731 11398
rect 4423 11387 4731 11396
rect 7896 10908 8204 10917
rect 7896 10906 7902 10908
rect 7958 10906 7982 10908
rect 8038 10906 8062 10908
rect 8118 10906 8142 10908
rect 8198 10906 8204 10908
rect 7958 10854 7960 10906
rect 8140 10854 8142 10906
rect 7896 10852 7902 10854
rect 7958 10852 7982 10854
rect 8038 10852 8062 10854
rect 8118 10852 8142 10854
rect 8198 10852 8204 10854
rect 7896 10843 8204 10852
rect 4423 10364 4731 10373
rect 4423 10362 4429 10364
rect 4485 10362 4509 10364
rect 4565 10362 4589 10364
rect 4645 10362 4669 10364
rect 4725 10362 4731 10364
rect 4485 10310 4487 10362
rect 4667 10310 4669 10362
rect 4423 10308 4429 10310
rect 4485 10308 4509 10310
rect 4565 10308 4589 10310
rect 4645 10308 4669 10310
rect 4725 10308 4731 10310
rect 4423 10299 4731 10308
rect 7896 9820 8204 9829
rect 7896 9818 7902 9820
rect 7958 9818 7982 9820
rect 8038 9818 8062 9820
rect 8118 9818 8142 9820
rect 8198 9818 8204 9820
rect 7958 9766 7960 9818
rect 8140 9766 8142 9818
rect 7896 9764 7902 9766
rect 7958 9764 7982 9766
rect 8038 9764 8062 9766
rect 8118 9764 8142 9766
rect 8198 9764 8204 9766
rect 7896 9755 8204 9764
rect 4423 9276 4731 9285
rect 4423 9274 4429 9276
rect 4485 9274 4509 9276
rect 4565 9274 4589 9276
rect 4645 9274 4669 9276
rect 4725 9274 4731 9276
rect 4485 9222 4487 9274
rect 4667 9222 4669 9274
rect 4423 9220 4429 9222
rect 4485 9220 4509 9222
rect 4565 9220 4589 9222
rect 4645 9220 4669 9222
rect 4725 9220 4731 9222
rect 4423 9211 4731 9220
rect 4344 8968 4396 8974
rect 4344 8910 4396 8916
rect 4356 8430 4384 8910
rect 7896 8732 8204 8741
rect 7896 8730 7902 8732
rect 7958 8730 7982 8732
rect 8038 8730 8062 8732
rect 8118 8730 8142 8732
rect 8198 8730 8204 8732
rect 7958 8678 7960 8730
rect 8140 8678 8142 8730
rect 7896 8676 7902 8678
rect 7958 8676 7982 8678
rect 8038 8676 8062 8678
rect 8118 8676 8142 8678
rect 8198 8676 8204 8678
rect 7896 8667 8204 8676
rect 4344 8424 4396 8430
rect 4344 8366 4396 8372
rect 4423 8188 4731 8197
rect 4423 8186 4429 8188
rect 4485 8186 4509 8188
rect 4565 8186 4589 8188
rect 4645 8186 4669 8188
rect 4725 8186 4731 8188
rect 4485 8134 4487 8186
rect 4667 8134 4669 8186
rect 4423 8132 4429 8134
rect 4485 8132 4509 8134
rect 4565 8132 4589 8134
rect 4645 8132 4669 8134
rect 4725 8132 4731 8134
rect 4423 8123 4731 8132
rect 5540 7948 5592 7954
rect 5540 7890 5592 7896
rect 4423 7100 4731 7109
rect 4423 7098 4429 7100
rect 4485 7098 4509 7100
rect 4565 7098 4589 7100
rect 4645 7098 4669 7100
rect 4725 7098 4731 7100
rect 4485 7046 4487 7098
rect 4667 7046 4669 7098
rect 4423 7044 4429 7046
rect 4485 7044 4509 7046
rect 4565 7044 4589 7046
rect 4645 7044 4669 7046
rect 4725 7044 4731 7046
rect 4423 7035 4731 7044
rect 4264 6886 4384 6914
rect 2964 6316 3016 6322
rect 2964 6258 3016 6264
rect 3620 6225 3648 6886
rect 4160 6248 4212 6254
rect 3606 6216 3662 6225
rect 4160 6190 4212 6196
rect 3606 6151 3662 6160
rect 4172 5794 4200 6190
rect 3056 5772 3108 5778
rect 3056 5714 3108 5720
rect 4080 5766 4200 5794
rect 2964 5160 3016 5166
rect 2964 5102 3016 5108
rect 2778 4856 2834 4865
rect 2976 4826 3004 5102
rect 2778 4791 2834 4800
rect 2964 4820 3016 4826
rect 2964 4762 3016 4768
rect 2872 4004 2924 4010
rect 2872 3946 2924 3952
rect 2688 3188 2740 3194
rect 2688 3130 2740 3136
rect 2596 2440 2648 2446
rect 2596 2382 2648 2388
rect 2700 2258 2728 3130
rect 2780 2984 2832 2990
rect 2780 2926 2832 2932
rect 2608 2230 2728 2258
rect 2608 800 2636 2230
rect 2792 1465 2820 2926
rect 2884 2825 2912 3946
rect 3068 3505 3096 5714
rect 3148 5160 3200 5166
rect 3148 5102 3200 5108
rect 3160 4146 3188 5102
rect 3700 4616 3752 4622
rect 3700 4558 3752 4564
rect 3712 4146 3740 4558
rect 4080 4185 4108 5766
rect 4160 5704 4212 5710
rect 4160 5646 4212 5652
rect 4066 4176 4122 4185
rect 3148 4140 3200 4146
rect 3148 4082 3200 4088
rect 3240 4140 3292 4146
rect 3240 4082 3292 4088
rect 3700 4140 3752 4146
rect 4066 4111 4122 4120
rect 3700 4082 3752 4088
rect 3252 3534 3280 4082
rect 3884 3664 3936 3670
rect 3884 3606 3936 3612
rect 3240 3528 3292 3534
rect 3054 3496 3110 3505
rect 3240 3470 3292 3476
rect 3054 3431 3110 3440
rect 2870 2816 2926 2825
rect 2870 2751 2926 2760
rect 3240 2508 3292 2514
rect 3240 2450 3292 2456
rect 2778 1456 2834 1465
rect 2778 1391 2834 1400
rect 3252 800 3280 2450
rect 3516 2304 3568 2310
rect 3516 2246 3568 2252
rect 3528 2145 3556 2246
rect 3514 2136 3570 2145
rect 3514 2071 3570 2080
rect 3896 800 3924 3606
rect 4172 3058 4200 5646
rect 4356 4706 4384 6886
rect 5356 6180 5408 6186
rect 5356 6122 5408 6128
rect 4423 6012 4731 6021
rect 4423 6010 4429 6012
rect 4485 6010 4509 6012
rect 4565 6010 4589 6012
rect 4645 6010 4669 6012
rect 4725 6010 4731 6012
rect 4485 5958 4487 6010
rect 4667 5958 4669 6010
rect 4423 5956 4429 5958
rect 4485 5956 4509 5958
rect 4565 5956 4589 5958
rect 4645 5956 4669 5958
rect 4725 5956 4731 5958
rect 4423 5947 4731 5956
rect 5368 5234 5396 6122
rect 5356 5228 5408 5234
rect 5356 5170 5408 5176
rect 4804 5160 4856 5166
rect 4804 5102 4856 5108
rect 4423 4924 4731 4933
rect 4423 4922 4429 4924
rect 4485 4922 4509 4924
rect 4565 4922 4589 4924
rect 4645 4922 4669 4924
rect 4725 4922 4731 4924
rect 4485 4870 4487 4922
rect 4667 4870 4669 4922
rect 4423 4868 4429 4870
rect 4485 4868 4509 4870
rect 4565 4868 4589 4870
rect 4645 4868 4669 4870
rect 4725 4868 4731 4870
rect 4423 4859 4731 4868
rect 4356 4678 4476 4706
rect 4448 4282 4476 4678
rect 4436 4276 4488 4282
rect 4436 4218 4488 4224
rect 4252 4072 4304 4078
rect 4252 4014 4304 4020
rect 4264 3738 4292 4014
rect 4448 4010 4476 4218
rect 4436 4004 4488 4010
rect 4436 3946 4488 3952
rect 4344 3936 4396 3942
rect 4344 3878 4396 3884
rect 4252 3732 4304 3738
rect 4252 3674 4304 3680
rect 4356 3126 4384 3878
rect 4423 3836 4731 3845
rect 4423 3834 4429 3836
rect 4485 3834 4509 3836
rect 4565 3834 4589 3836
rect 4645 3834 4669 3836
rect 4725 3834 4731 3836
rect 4485 3782 4487 3834
rect 4667 3782 4669 3834
rect 4423 3780 4429 3782
rect 4485 3780 4509 3782
rect 4565 3780 4589 3782
rect 4645 3780 4669 3782
rect 4725 3780 4731 3782
rect 4423 3771 4731 3780
rect 4816 3194 4844 5102
rect 5448 5024 5500 5030
rect 5448 4966 5500 4972
rect 5460 4690 5488 4966
rect 5448 4684 5500 4690
rect 5448 4626 5500 4632
rect 5552 3670 5580 7890
rect 7896 7644 8204 7653
rect 7896 7642 7902 7644
rect 7958 7642 7982 7644
rect 8038 7642 8062 7644
rect 8118 7642 8142 7644
rect 8198 7642 8204 7644
rect 7958 7590 7960 7642
rect 8140 7590 8142 7642
rect 7896 7588 7902 7590
rect 7958 7588 7982 7590
rect 8038 7588 8062 7590
rect 8118 7588 8142 7590
rect 8198 7588 8204 7590
rect 7896 7579 8204 7588
rect 7896 6556 8204 6565
rect 7896 6554 7902 6556
rect 7958 6554 7982 6556
rect 8038 6554 8062 6556
rect 8118 6554 8142 6556
rect 8198 6554 8204 6556
rect 7958 6502 7960 6554
rect 8140 6502 8142 6554
rect 7896 6500 7902 6502
rect 7958 6500 7982 6502
rect 8038 6500 8062 6502
rect 8118 6500 8142 6502
rect 8198 6500 8204 6502
rect 7896 6491 8204 6500
rect 7896 5468 8204 5477
rect 7896 5466 7902 5468
rect 7958 5466 7982 5468
rect 8038 5466 8062 5468
rect 8118 5466 8142 5468
rect 8198 5466 8204 5468
rect 7958 5414 7960 5466
rect 8140 5414 8142 5466
rect 7896 5412 7902 5414
rect 7958 5412 7982 5414
rect 8038 5412 8062 5414
rect 8118 5412 8142 5414
rect 8198 5412 8204 5414
rect 7896 5403 8204 5412
rect 5816 4684 5868 4690
rect 5816 4626 5868 4632
rect 5540 3664 5592 3670
rect 5540 3606 5592 3612
rect 4804 3188 4856 3194
rect 4804 3130 4856 3136
rect 4344 3120 4396 3126
rect 4344 3062 4396 3068
rect 4160 3052 4212 3058
rect 4160 2994 4212 3000
rect 4804 2984 4856 2990
rect 4804 2926 4856 2932
rect 4423 2748 4731 2757
rect 4423 2746 4429 2748
rect 4485 2746 4509 2748
rect 4565 2746 4589 2748
rect 4645 2746 4669 2748
rect 4725 2746 4731 2748
rect 4485 2694 4487 2746
rect 4667 2694 4669 2746
rect 4423 2692 4429 2694
rect 4485 2692 4509 2694
rect 4565 2692 4589 2694
rect 4645 2692 4669 2694
rect 4725 2692 4731 2694
rect 4423 2683 4731 2692
rect 4816 1714 4844 2926
rect 4540 1686 4844 1714
rect 4540 800 4568 1686
rect 5828 800 5856 4626
rect 7896 4380 8204 4389
rect 7896 4378 7902 4380
rect 7958 4378 7982 4380
rect 8038 4378 8062 4380
rect 8118 4378 8142 4380
rect 8198 4378 8204 4380
rect 7958 4326 7960 4378
rect 8140 4326 8142 4378
rect 7896 4324 7902 4326
rect 7958 4324 7982 4326
rect 8038 4324 8062 4326
rect 8118 4324 8142 4326
rect 8198 4324 8204 4326
rect 7896 4315 8204 4324
rect 5908 3936 5960 3942
rect 5908 3878 5960 3884
rect 6920 3936 6972 3942
rect 6920 3878 6972 3884
rect 5920 3602 5948 3878
rect 5908 3596 5960 3602
rect 5908 3538 5960 3544
rect 6460 3596 6512 3602
rect 6460 3538 6512 3544
rect 6472 800 6500 3538
rect 6932 2990 6960 3878
rect 7104 3392 7156 3398
rect 7104 3334 7156 3340
rect 7116 3126 7144 3334
rect 7896 3292 8204 3301
rect 7896 3290 7902 3292
rect 7958 3290 7982 3292
rect 8038 3290 8062 3292
rect 8118 3290 8142 3292
rect 8198 3290 8204 3292
rect 7958 3238 7960 3290
rect 8140 3238 8142 3290
rect 7896 3236 7902 3238
rect 7958 3236 7982 3238
rect 8038 3236 8062 3238
rect 8118 3236 8142 3238
rect 8198 3236 8204 3238
rect 7896 3227 8204 3236
rect 7104 3120 7156 3126
rect 7104 3062 7156 3068
rect 6920 2984 6972 2990
rect 6920 2926 6972 2932
rect 8312 2310 8340 13806
rect 9404 8356 9456 8362
rect 9404 8298 9456 8304
rect 9220 3528 9272 3534
rect 9220 3470 9272 3476
rect 9232 3058 9260 3470
rect 9416 3126 9444 8298
rect 9404 3120 9456 3126
rect 9404 3062 9456 3068
rect 9220 3052 9272 3058
rect 9220 2994 9272 3000
rect 8392 2984 8444 2990
rect 8392 2926 8444 2932
rect 8300 2304 8352 2310
rect 8300 2246 8352 2252
rect 7896 2204 8204 2213
rect 7896 2202 7902 2204
rect 7958 2202 7982 2204
rect 8038 2202 8062 2204
rect 8118 2202 8142 2204
rect 8198 2202 8204 2204
rect 7958 2150 7960 2202
rect 8140 2150 8142 2202
rect 7896 2148 7902 2150
rect 7958 2148 7982 2150
rect 8038 2148 8062 2150
rect 8118 2148 8142 2150
rect 8198 2148 8204 2150
rect 7896 2139 8204 2148
rect 8404 800 8432 2926
rect 9508 2514 9536 25094
rect 11369 24508 11677 24517
rect 11369 24506 11375 24508
rect 11431 24506 11455 24508
rect 11511 24506 11535 24508
rect 11591 24506 11615 24508
rect 11671 24506 11677 24508
rect 11431 24454 11433 24506
rect 11613 24454 11615 24506
rect 11369 24452 11375 24454
rect 11431 24452 11455 24454
rect 11511 24452 11535 24454
rect 11591 24452 11615 24454
rect 11671 24452 11677 24454
rect 11369 24443 11677 24452
rect 11369 23420 11677 23429
rect 11369 23418 11375 23420
rect 11431 23418 11455 23420
rect 11511 23418 11535 23420
rect 11591 23418 11615 23420
rect 11671 23418 11677 23420
rect 11431 23366 11433 23418
rect 11613 23366 11615 23418
rect 11369 23364 11375 23366
rect 11431 23364 11455 23366
rect 11511 23364 11535 23366
rect 11591 23364 11615 23366
rect 11671 23364 11677 23366
rect 11369 23355 11677 23364
rect 11369 22332 11677 22341
rect 11369 22330 11375 22332
rect 11431 22330 11455 22332
rect 11511 22330 11535 22332
rect 11591 22330 11615 22332
rect 11671 22330 11677 22332
rect 11431 22278 11433 22330
rect 11613 22278 11615 22330
rect 11369 22276 11375 22278
rect 11431 22276 11455 22278
rect 11511 22276 11535 22278
rect 11591 22276 11615 22278
rect 11671 22276 11677 22278
rect 11369 22267 11677 22276
rect 11369 21244 11677 21253
rect 11369 21242 11375 21244
rect 11431 21242 11455 21244
rect 11511 21242 11535 21244
rect 11591 21242 11615 21244
rect 11671 21242 11677 21244
rect 11431 21190 11433 21242
rect 11613 21190 11615 21242
rect 11369 21188 11375 21190
rect 11431 21188 11455 21190
rect 11511 21188 11535 21190
rect 11591 21188 11615 21190
rect 11671 21188 11677 21190
rect 11369 21179 11677 21188
rect 11369 20156 11677 20165
rect 11369 20154 11375 20156
rect 11431 20154 11455 20156
rect 11511 20154 11535 20156
rect 11591 20154 11615 20156
rect 11671 20154 11677 20156
rect 11431 20102 11433 20154
rect 11613 20102 11615 20154
rect 11369 20100 11375 20102
rect 11431 20100 11455 20102
rect 11511 20100 11535 20102
rect 11591 20100 11615 20102
rect 11671 20100 11677 20102
rect 11369 20091 11677 20100
rect 11369 19068 11677 19077
rect 11369 19066 11375 19068
rect 11431 19066 11455 19068
rect 11511 19066 11535 19068
rect 11591 19066 11615 19068
rect 11671 19066 11677 19068
rect 11431 19014 11433 19066
rect 11613 19014 11615 19066
rect 11369 19012 11375 19014
rect 11431 19012 11455 19014
rect 11511 19012 11535 19014
rect 11591 19012 11615 19014
rect 11671 19012 11677 19014
rect 11369 19003 11677 19012
rect 11369 17980 11677 17989
rect 11369 17978 11375 17980
rect 11431 17978 11455 17980
rect 11511 17978 11535 17980
rect 11591 17978 11615 17980
rect 11671 17978 11677 17980
rect 11431 17926 11433 17978
rect 11613 17926 11615 17978
rect 11369 17924 11375 17926
rect 11431 17924 11455 17926
rect 11511 17924 11535 17926
rect 11591 17924 11615 17926
rect 11671 17924 11677 17926
rect 11369 17915 11677 17924
rect 11369 16892 11677 16901
rect 11369 16890 11375 16892
rect 11431 16890 11455 16892
rect 11511 16890 11535 16892
rect 11591 16890 11615 16892
rect 11671 16890 11677 16892
rect 11431 16838 11433 16890
rect 11613 16838 11615 16890
rect 11369 16836 11375 16838
rect 11431 16836 11455 16838
rect 11511 16836 11535 16838
rect 11591 16836 11615 16838
rect 11671 16836 11677 16838
rect 11369 16827 11677 16836
rect 11369 15804 11677 15813
rect 11369 15802 11375 15804
rect 11431 15802 11455 15804
rect 11511 15802 11535 15804
rect 11591 15802 11615 15804
rect 11671 15802 11677 15804
rect 11431 15750 11433 15802
rect 11613 15750 11615 15802
rect 11369 15748 11375 15750
rect 11431 15748 11455 15750
rect 11511 15748 11535 15750
rect 11591 15748 11615 15750
rect 11671 15748 11677 15750
rect 11369 15739 11677 15748
rect 12624 14884 12676 14890
rect 12624 14826 12676 14832
rect 11369 14716 11677 14725
rect 11369 14714 11375 14716
rect 11431 14714 11455 14716
rect 11511 14714 11535 14716
rect 11591 14714 11615 14716
rect 11671 14714 11677 14716
rect 11431 14662 11433 14714
rect 11613 14662 11615 14714
rect 11369 14660 11375 14662
rect 11431 14660 11455 14662
rect 11511 14660 11535 14662
rect 11591 14660 11615 14662
rect 11671 14660 11677 14662
rect 11369 14651 11677 14660
rect 12636 14482 12664 14826
rect 9680 14476 9732 14482
rect 9680 14418 9732 14424
rect 12624 14476 12676 14482
rect 12624 14418 12676 14424
rect 9692 12442 9720 14418
rect 10968 14340 11020 14346
rect 10968 14282 11020 14288
rect 11244 14340 11296 14346
rect 11244 14282 11296 14288
rect 9956 14272 10008 14278
rect 9956 14214 10008 14220
rect 9968 14006 9996 14214
rect 9956 14000 10008 14006
rect 9956 13942 10008 13948
rect 10980 13938 11008 14282
rect 10968 13932 11020 13938
rect 10968 13874 11020 13880
rect 11256 13530 11284 14282
rect 11369 13628 11677 13637
rect 11369 13626 11375 13628
rect 11431 13626 11455 13628
rect 11511 13626 11535 13628
rect 11591 13626 11615 13628
rect 11671 13626 11677 13628
rect 11431 13574 11433 13626
rect 11613 13574 11615 13626
rect 11369 13572 11375 13574
rect 11431 13572 11455 13574
rect 11511 13572 11535 13574
rect 11591 13572 11615 13574
rect 11671 13572 11677 13574
rect 11369 13563 11677 13572
rect 11244 13524 11296 13530
rect 11244 13466 11296 13472
rect 9772 13320 9824 13326
rect 9772 13262 9824 13268
rect 9680 12436 9732 12442
rect 9680 12378 9732 12384
rect 9784 11150 9812 13262
rect 11369 12540 11677 12549
rect 11369 12538 11375 12540
rect 11431 12538 11455 12540
rect 11511 12538 11535 12540
rect 11591 12538 11615 12540
rect 11671 12538 11677 12540
rect 11431 12486 11433 12538
rect 11613 12486 11615 12538
rect 11369 12484 11375 12486
rect 11431 12484 11455 12486
rect 11511 12484 11535 12486
rect 11591 12484 11615 12486
rect 11671 12484 11677 12486
rect 11369 12475 11677 12484
rect 11369 11452 11677 11461
rect 11369 11450 11375 11452
rect 11431 11450 11455 11452
rect 11511 11450 11535 11452
rect 11591 11450 11615 11452
rect 11671 11450 11677 11452
rect 11431 11398 11433 11450
rect 11613 11398 11615 11450
rect 11369 11396 11375 11398
rect 11431 11396 11455 11398
rect 11511 11396 11535 11398
rect 11591 11396 11615 11398
rect 11671 11396 11677 11398
rect 11369 11387 11677 11396
rect 9772 11144 9824 11150
rect 9772 11086 9824 11092
rect 11369 10364 11677 10373
rect 11369 10362 11375 10364
rect 11431 10362 11455 10364
rect 11511 10362 11535 10364
rect 11591 10362 11615 10364
rect 11671 10362 11677 10364
rect 11431 10310 11433 10362
rect 11613 10310 11615 10362
rect 11369 10308 11375 10310
rect 11431 10308 11455 10310
rect 11511 10308 11535 10310
rect 11591 10308 11615 10310
rect 11671 10308 11677 10310
rect 11369 10299 11677 10308
rect 11369 9276 11677 9285
rect 11369 9274 11375 9276
rect 11431 9274 11455 9276
rect 11511 9274 11535 9276
rect 11591 9274 11615 9276
rect 11671 9274 11677 9276
rect 11431 9222 11433 9274
rect 11613 9222 11615 9274
rect 11369 9220 11375 9222
rect 11431 9220 11455 9222
rect 11511 9220 11535 9222
rect 11591 9220 11615 9222
rect 11671 9220 11677 9222
rect 11369 9211 11677 9220
rect 12728 8566 12756 35226
rect 14384 35018 14412 44338
rect 14842 43548 15150 43557
rect 14842 43546 14848 43548
rect 14904 43546 14928 43548
rect 14984 43546 15008 43548
rect 15064 43546 15088 43548
rect 15144 43546 15150 43548
rect 14904 43494 14906 43546
rect 15086 43494 15088 43546
rect 14842 43492 14848 43494
rect 14904 43492 14928 43494
rect 14984 43492 15008 43494
rect 15064 43492 15088 43494
rect 15144 43492 15150 43494
rect 14842 43483 15150 43492
rect 15856 43450 15884 45766
rect 18340 45626 18368 45902
rect 22572 45898 22600 49200
rect 22836 47048 22888 47054
rect 22836 46990 22888 46996
rect 22848 46578 22876 46990
rect 22836 46572 22888 46578
rect 22836 46514 22888 46520
rect 23216 46510 23244 49200
rect 23756 47184 23808 47190
rect 23756 47126 23808 47132
rect 23480 46912 23532 46918
rect 23480 46854 23532 46860
rect 23112 46504 23164 46510
rect 23112 46446 23164 46452
rect 23204 46504 23256 46510
rect 23204 46446 23256 46452
rect 23124 46170 23152 46446
rect 23112 46164 23164 46170
rect 23112 46106 23164 46112
rect 23204 45960 23256 45966
rect 23204 45902 23256 45908
rect 20444 45892 20496 45898
rect 20444 45834 20496 45840
rect 21272 45892 21324 45898
rect 21272 45834 21324 45840
rect 22560 45892 22612 45898
rect 22560 45834 22612 45840
rect 20352 45824 20404 45830
rect 20352 45766 20404 45772
rect 18328 45620 18380 45626
rect 18328 45562 18380 45568
rect 20364 45490 20392 45766
rect 20456 45626 20484 45834
rect 20444 45620 20496 45626
rect 20444 45562 20496 45568
rect 20352 45484 20404 45490
rect 20352 45426 20404 45432
rect 20364 45286 20392 45426
rect 20352 45280 20404 45286
rect 20352 45222 20404 45228
rect 18315 45180 18623 45189
rect 18315 45178 18321 45180
rect 18377 45178 18401 45180
rect 18457 45178 18481 45180
rect 18537 45178 18561 45180
rect 18617 45178 18623 45180
rect 18377 45126 18379 45178
rect 18559 45126 18561 45178
rect 18315 45124 18321 45126
rect 18377 45124 18401 45126
rect 18457 45124 18481 45126
rect 18537 45124 18561 45126
rect 18617 45124 18623 45126
rect 18315 45115 18623 45124
rect 19340 44396 19392 44402
rect 19340 44338 19392 44344
rect 18315 44092 18623 44101
rect 18315 44090 18321 44092
rect 18377 44090 18401 44092
rect 18457 44090 18481 44092
rect 18537 44090 18561 44092
rect 18617 44090 18623 44092
rect 18377 44038 18379 44090
rect 18559 44038 18561 44090
rect 18315 44036 18321 44038
rect 18377 44036 18401 44038
rect 18457 44036 18481 44038
rect 18537 44036 18561 44038
rect 18617 44036 18623 44038
rect 18315 44027 18623 44036
rect 15844 43444 15896 43450
rect 15844 43386 15896 43392
rect 19352 43314 19380 44338
rect 21284 43858 21312 45834
rect 21788 45724 22096 45733
rect 21788 45722 21794 45724
rect 21850 45722 21874 45724
rect 21930 45722 21954 45724
rect 22010 45722 22034 45724
rect 22090 45722 22096 45724
rect 21850 45670 21852 45722
rect 22032 45670 22034 45722
rect 21788 45668 21794 45670
rect 21850 45668 21874 45670
rect 21930 45668 21954 45670
rect 22010 45668 22034 45670
rect 22090 45668 22096 45670
rect 21788 45659 22096 45668
rect 21640 45280 21692 45286
rect 21640 45222 21692 45228
rect 21272 43852 21324 43858
rect 21272 43794 21324 43800
rect 19432 43784 19484 43790
rect 19432 43726 19484 43732
rect 19340 43308 19392 43314
rect 19340 43250 19392 43256
rect 18315 43004 18623 43013
rect 18315 43002 18321 43004
rect 18377 43002 18401 43004
rect 18457 43002 18481 43004
rect 18537 43002 18561 43004
rect 18617 43002 18623 43004
rect 18377 42950 18379 43002
rect 18559 42950 18561 43002
rect 18315 42948 18321 42950
rect 18377 42948 18401 42950
rect 18457 42948 18481 42950
rect 18537 42948 18561 42950
rect 18617 42948 18623 42950
rect 18315 42939 18623 42948
rect 19444 42945 19472 43726
rect 19616 43716 19668 43722
rect 19616 43658 19668 43664
rect 19628 43450 19656 43658
rect 19616 43444 19668 43450
rect 19616 43386 19668 43392
rect 19430 42936 19486 42945
rect 19430 42871 19486 42880
rect 14842 42460 15150 42469
rect 14842 42458 14848 42460
rect 14904 42458 14928 42460
rect 14984 42458 15008 42460
rect 15064 42458 15088 42460
rect 15144 42458 15150 42460
rect 14904 42406 14906 42458
rect 15086 42406 15088 42458
rect 14842 42404 14848 42406
rect 14904 42404 14928 42406
rect 14984 42404 15008 42406
rect 15064 42404 15088 42406
rect 15144 42404 15150 42406
rect 14842 42395 15150 42404
rect 18315 41916 18623 41925
rect 18315 41914 18321 41916
rect 18377 41914 18401 41916
rect 18457 41914 18481 41916
rect 18537 41914 18561 41916
rect 18617 41914 18623 41916
rect 18377 41862 18379 41914
rect 18559 41862 18561 41914
rect 18315 41860 18321 41862
rect 18377 41860 18401 41862
rect 18457 41860 18481 41862
rect 18537 41860 18561 41862
rect 18617 41860 18623 41862
rect 18315 41851 18623 41860
rect 14842 41372 15150 41381
rect 14842 41370 14848 41372
rect 14904 41370 14928 41372
rect 14984 41370 15008 41372
rect 15064 41370 15088 41372
rect 15144 41370 15150 41372
rect 14904 41318 14906 41370
rect 15086 41318 15088 41370
rect 14842 41316 14848 41318
rect 14904 41316 14928 41318
rect 14984 41316 15008 41318
rect 15064 41316 15088 41318
rect 15144 41316 15150 41318
rect 14842 41307 15150 41316
rect 18315 40828 18623 40837
rect 18315 40826 18321 40828
rect 18377 40826 18401 40828
rect 18457 40826 18481 40828
rect 18537 40826 18561 40828
rect 18617 40826 18623 40828
rect 18377 40774 18379 40826
rect 18559 40774 18561 40826
rect 18315 40772 18321 40774
rect 18377 40772 18401 40774
rect 18457 40772 18481 40774
rect 18537 40772 18561 40774
rect 18617 40772 18623 40774
rect 18315 40763 18623 40772
rect 17868 40520 17920 40526
rect 17868 40462 17920 40468
rect 18604 40520 18656 40526
rect 18604 40462 18656 40468
rect 17500 40384 17552 40390
rect 17500 40326 17552 40332
rect 14842 40284 15150 40293
rect 14842 40282 14848 40284
rect 14904 40282 14928 40284
rect 14984 40282 15008 40284
rect 15064 40282 15088 40284
rect 15144 40282 15150 40284
rect 14904 40230 14906 40282
rect 15086 40230 15088 40282
rect 14842 40228 14848 40230
rect 14904 40228 14928 40230
rect 14984 40228 15008 40230
rect 15064 40228 15088 40230
rect 15144 40228 15150 40230
rect 14842 40219 15150 40228
rect 17512 40050 17540 40326
rect 17880 40118 17908 40462
rect 18236 40452 18288 40458
rect 18236 40394 18288 40400
rect 17868 40112 17920 40118
rect 17868 40054 17920 40060
rect 17224 40044 17276 40050
rect 17224 39986 17276 39992
rect 17500 40044 17552 40050
rect 17500 39986 17552 39992
rect 16304 39976 16356 39982
rect 16304 39918 16356 39924
rect 14842 39196 15150 39205
rect 14842 39194 14848 39196
rect 14904 39194 14928 39196
rect 14984 39194 15008 39196
rect 15064 39194 15088 39196
rect 15144 39194 15150 39196
rect 14904 39142 14906 39194
rect 15086 39142 15088 39194
rect 14842 39140 14848 39142
rect 14904 39140 14928 39142
rect 14984 39140 15008 39142
rect 15064 39140 15088 39142
rect 15144 39140 15150 39142
rect 14842 39131 15150 39140
rect 15292 38548 15344 38554
rect 15292 38490 15344 38496
rect 15304 38282 15332 38490
rect 16120 38480 16172 38486
rect 16120 38422 16172 38428
rect 15476 38412 15528 38418
rect 15476 38354 15528 38360
rect 15844 38412 15896 38418
rect 15844 38354 15896 38360
rect 15292 38276 15344 38282
rect 15292 38218 15344 38224
rect 14842 38108 15150 38117
rect 14842 38106 14848 38108
rect 14904 38106 14928 38108
rect 14984 38106 15008 38108
rect 15064 38106 15088 38108
rect 15144 38106 15150 38108
rect 14904 38054 14906 38106
rect 15086 38054 15088 38106
rect 14842 38052 14848 38054
rect 14904 38052 14928 38054
rect 14984 38052 15008 38054
rect 15064 38052 15088 38054
rect 15144 38052 15150 38054
rect 14842 38043 15150 38052
rect 14842 37020 15150 37029
rect 14842 37018 14848 37020
rect 14904 37018 14928 37020
rect 14984 37018 15008 37020
rect 15064 37018 15088 37020
rect 15144 37018 15150 37020
rect 14904 36966 14906 37018
rect 15086 36966 15088 37018
rect 14842 36964 14848 36966
rect 14904 36964 14928 36966
rect 14984 36964 15008 36966
rect 15064 36964 15088 36966
rect 15144 36964 15150 36966
rect 14842 36955 15150 36964
rect 14842 35932 15150 35941
rect 14842 35930 14848 35932
rect 14904 35930 14928 35932
rect 14984 35930 15008 35932
rect 15064 35930 15088 35932
rect 15144 35930 15150 35932
rect 14904 35878 14906 35930
rect 15086 35878 15088 35930
rect 14842 35876 14848 35878
rect 14904 35876 14928 35878
rect 14984 35876 15008 35878
rect 15064 35876 15088 35878
rect 15144 35876 15150 35878
rect 14842 35867 15150 35876
rect 14372 35012 14424 35018
rect 14372 34954 14424 34960
rect 12808 34536 12860 34542
rect 12808 34478 12860 34484
rect 12820 31958 12848 34478
rect 13820 33312 13872 33318
rect 13820 33254 13872 33260
rect 13832 32366 13860 33254
rect 12900 32360 12952 32366
rect 12900 32302 12952 32308
rect 13820 32360 13872 32366
rect 13820 32302 13872 32308
rect 12912 32026 12940 32302
rect 13268 32292 13320 32298
rect 13268 32234 13320 32240
rect 12900 32020 12952 32026
rect 12900 31962 12952 31968
rect 12808 31952 12860 31958
rect 12808 31894 12860 31900
rect 13280 16794 13308 32234
rect 14384 27470 14412 34954
rect 14842 34844 15150 34853
rect 14842 34842 14848 34844
rect 14904 34842 14928 34844
rect 14984 34842 15008 34844
rect 15064 34842 15088 34844
rect 15144 34842 15150 34844
rect 14904 34790 14906 34842
rect 15086 34790 15088 34842
rect 14842 34788 14848 34790
rect 14904 34788 14928 34790
rect 14984 34788 15008 34790
rect 15064 34788 15088 34790
rect 15144 34788 15150 34790
rect 14842 34779 15150 34788
rect 14842 33756 15150 33765
rect 14842 33754 14848 33756
rect 14904 33754 14928 33756
rect 14984 33754 15008 33756
rect 15064 33754 15088 33756
rect 15144 33754 15150 33756
rect 14904 33702 14906 33754
rect 15086 33702 15088 33754
rect 14842 33700 14848 33702
rect 14904 33700 14928 33702
rect 14984 33700 15008 33702
rect 15064 33700 15088 33702
rect 15144 33700 15150 33702
rect 14842 33691 15150 33700
rect 14842 32668 15150 32677
rect 14842 32666 14848 32668
rect 14904 32666 14928 32668
rect 14984 32666 15008 32668
rect 15064 32666 15088 32668
rect 15144 32666 15150 32668
rect 14904 32614 14906 32666
rect 15086 32614 15088 32666
rect 14842 32612 14848 32614
rect 14904 32612 14928 32614
rect 14984 32612 15008 32614
rect 15064 32612 15088 32614
rect 15144 32612 15150 32614
rect 14842 32603 15150 32612
rect 14842 31580 15150 31589
rect 14842 31578 14848 31580
rect 14904 31578 14928 31580
rect 14984 31578 15008 31580
rect 15064 31578 15088 31580
rect 15144 31578 15150 31580
rect 14904 31526 14906 31578
rect 15086 31526 15088 31578
rect 14842 31524 14848 31526
rect 14904 31524 14928 31526
rect 14984 31524 15008 31526
rect 15064 31524 15088 31526
rect 15144 31524 15150 31526
rect 14842 31515 15150 31524
rect 14842 30492 15150 30501
rect 14842 30490 14848 30492
rect 14904 30490 14928 30492
rect 14984 30490 15008 30492
rect 15064 30490 15088 30492
rect 15144 30490 15150 30492
rect 14904 30438 14906 30490
rect 15086 30438 15088 30490
rect 14842 30436 14848 30438
rect 14904 30436 14928 30438
rect 14984 30436 15008 30438
rect 15064 30436 15088 30438
rect 15144 30436 15150 30438
rect 14842 30427 15150 30436
rect 14842 29404 15150 29413
rect 14842 29402 14848 29404
rect 14904 29402 14928 29404
rect 14984 29402 15008 29404
rect 15064 29402 15088 29404
rect 15144 29402 15150 29404
rect 14904 29350 14906 29402
rect 15086 29350 15088 29402
rect 14842 29348 14848 29350
rect 14904 29348 14928 29350
rect 14984 29348 15008 29350
rect 15064 29348 15088 29350
rect 15144 29348 15150 29350
rect 14842 29339 15150 29348
rect 14842 28316 15150 28325
rect 14842 28314 14848 28316
rect 14904 28314 14928 28316
rect 14984 28314 15008 28316
rect 15064 28314 15088 28316
rect 15144 28314 15150 28316
rect 14904 28262 14906 28314
rect 15086 28262 15088 28314
rect 14842 28260 14848 28262
rect 14904 28260 14928 28262
rect 14984 28260 15008 28262
rect 15064 28260 15088 28262
rect 15144 28260 15150 28262
rect 14842 28251 15150 28260
rect 15200 28008 15252 28014
rect 15200 27950 15252 27956
rect 15212 27606 15240 27950
rect 15200 27600 15252 27606
rect 15200 27542 15252 27548
rect 14372 27464 14424 27470
rect 14372 27406 14424 27412
rect 14384 19786 14412 27406
rect 14842 27228 15150 27237
rect 14842 27226 14848 27228
rect 14904 27226 14928 27228
rect 14984 27226 15008 27228
rect 15064 27226 15088 27228
rect 15144 27226 15150 27228
rect 14904 27174 14906 27226
rect 15086 27174 15088 27226
rect 14842 27172 14848 27174
rect 14904 27172 14928 27174
rect 14984 27172 15008 27174
rect 15064 27172 15088 27174
rect 15144 27172 15150 27174
rect 14842 27163 15150 27172
rect 14842 26140 15150 26149
rect 14842 26138 14848 26140
rect 14904 26138 14928 26140
rect 14984 26138 15008 26140
rect 15064 26138 15088 26140
rect 15144 26138 15150 26140
rect 14904 26086 14906 26138
rect 15086 26086 15088 26138
rect 14842 26084 14848 26086
rect 14904 26084 14928 26086
rect 14984 26084 15008 26086
rect 15064 26084 15088 26086
rect 15144 26084 15150 26086
rect 14842 26075 15150 26084
rect 14842 25052 15150 25061
rect 14842 25050 14848 25052
rect 14904 25050 14928 25052
rect 14984 25050 15008 25052
rect 15064 25050 15088 25052
rect 15144 25050 15150 25052
rect 14904 24998 14906 25050
rect 15086 24998 15088 25050
rect 14842 24996 14848 24998
rect 14904 24996 14928 24998
rect 14984 24996 15008 24998
rect 15064 24996 15088 24998
rect 15144 24996 15150 24998
rect 14842 24987 15150 24996
rect 14842 23964 15150 23973
rect 14842 23962 14848 23964
rect 14904 23962 14928 23964
rect 14984 23962 15008 23964
rect 15064 23962 15088 23964
rect 15144 23962 15150 23964
rect 14904 23910 14906 23962
rect 15086 23910 15088 23962
rect 14842 23908 14848 23910
rect 14904 23908 14928 23910
rect 14984 23908 15008 23910
rect 15064 23908 15088 23910
rect 15144 23908 15150 23910
rect 14842 23899 15150 23908
rect 14842 22876 15150 22885
rect 14842 22874 14848 22876
rect 14904 22874 14928 22876
rect 14984 22874 15008 22876
rect 15064 22874 15088 22876
rect 15144 22874 15150 22876
rect 14904 22822 14906 22874
rect 15086 22822 15088 22874
rect 14842 22820 14848 22822
rect 14904 22820 14928 22822
rect 14984 22820 15008 22822
rect 15064 22820 15088 22822
rect 15144 22820 15150 22822
rect 14842 22811 15150 22820
rect 14842 21788 15150 21797
rect 14842 21786 14848 21788
rect 14904 21786 14928 21788
rect 14984 21786 15008 21788
rect 15064 21786 15088 21788
rect 15144 21786 15150 21788
rect 14904 21734 14906 21786
rect 15086 21734 15088 21786
rect 14842 21732 14848 21734
rect 14904 21732 14928 21734
rect 14984 21732 15008 21734
rect 15064 21732 15088 21734
rect 15144 21732 15150 21734
rect 14842 21723 15150 21732
rect 14842 20700 15150 20709
rect 14842 20698 14848 20700
rect 14904 20698 14928 20700
rect 14984 20698 15008 20700
rect 15064 20698 15088 20700
rect 15144 20698 15150 20700
rect 14904 20646 14906 20698
rect 15086 20646 15088 20698
rect 14842 20644 14848 20646
rect 14904 20644 14928 20646
rect 14984 20644 15008 20646
rect 15064 20644 15088 20646
rect 15144 20644 15150 20646
rect 14842 20635 15150 20644
rect 15200 20460 15252 20466
rect 15200 20402 15252 20408
rect 15212 20058 15240 20402
rect 15304 20262 15332 38218
rect 15488 38010 15516 38354
rect 15476 38004 15528 38010
rect 15476 37946 15528 37952
rect 15476 37324 15528 37330
rect 15476 37266 15528 37272
rect 15488 26450 15516 37266
rect 15752 36576 15804 36582
rect 15752 36518 15804 36524
rect 15764 35698 15792 36518
rect 15752 35692 15804 35698
rect 15752 35634 15804 35640
rect 15568 35624 15620 35630
rect 15568 35566 15620 35572
rect 15580 34746 15608 35566
rect 15568 34740 15620 34746
rect 15568 34682 15620 34688
rect 15856 33522 15884 38354
rect 16132 38350 16160 38422
rect 16120 38344 16172 38350
rect 16120 38286 16172 38292
rect 16028 38208 16080 38214
rect 16028 38150 16080 38156
rect 16040 37874 16068 38150
rect 16028 37868 16080 37874
rect 16028 37810 16080 37816
rect 16132 37194 16160 38286
rect 16212 37392 16264 37398
rect 16212 37334 16264 37340
rect 16120 37188 16172 37194
rect 16120 37130 16172 37136
rect 16028 37120 16080 37126
rect 16028 37062 16080 37068
rect 16040 34610 16068 37062
rect 16028 34604 16080 34610
rect 16028 34546 16080 34552
rect 16028 34400 16080 34406
rect 16028 34342 16080 34348
rect 16040 33998 16068 34342
rect 16028 33992 16080 33998
rect 16028 33934 16080 33940
rect 16132 33522 16160 37130
rect 16224 36718 16252 37334
rect 16212 36712 16264 36718
rect 16212 36654 16264 36660
rect 16212 33856 16264 33862
rect 16212 33798 16264 33804
rect 16224 33590 16252 33798
rect 16212 33584 16264 33590
rect 16212 33526 16264 33532
rect 15752 33516 15804 33522
rect 15752 33458 15804 33464
rect 15844 33516 15896 33522
rect 15844 33458 15896 33464
rect 16120 33516 16172 33522
rect 16120 33458 16172 33464
rect 15764 33046 15792 33458
rect 15752 33040 15804 33046
rect 15752 32982 15804 32988
rect 15856 30938 15884 33458
rect 16028 33312 16080 33318
rect 16028 33254 16080 33260
rect 16040 32910 16068 33254
rect 16028 32904 16080 32910
rect 16028 32846 16080 32852
rect 15844 30932 15896 30938
rect 15844 30874 15896 30880
rect 15856 30190 15884 30874
rect 15844 30184 15896 30190
rect 15844 30126 15896 30132
rect 16040 28762 16068 32846
rect 16212 31476 16264 31482
rect 16316 31464 16344 39918
rect 17040 39840 17092 39846
rect 17040 39782 17092 39788
rect 16396 37868 16448 37874
rect 16396 37810 16448 37816
rect 16408 32774 16436 37810
rect 16580 37800 16632 37806
rect 16580 37742 16632 37748
rect 16592 37194 16620 37742
rect 16948 37664 17000 37670
rect 16948 37606 17000 37612
rect 16580 37188 16632 37194
rect 16580 37130 16632 37136
rect 16592 33658 16620 37130
rect 16580 33652 16632 33658
rect 16580 33594 16632 33600
rect 16764 33108 16816 33114
rect 16764 33050 16816 33056
rect 16488 33040 16540 33046
rect 16488 32982 16540 32988
rect 16396 32768 16448 32774
rect 16396 32710 16448 32716
rect 16500 31890 16528 32982
rect 16776 32910 16804 33050
rect 16764 32904 16816 32910
rect 16764 32846 16816 32852
rect 16580 32020 16632 32026
rect 16580 31962 16632 31968
rect 16592 31906 16620 31962
rect 16488 31884 16540 31890
rect 16592 31878 16712 31906
rect 16488 31826 16540 31832
rect 16580 31816 16632 31822
rect 16580 31758 16632 31764
rect 16264 31436 16344 31464
rect 16212 31418 16264 31424
rect 16316 30802 16344 31436
rect 16592 31210 16620 31758
rect 16684 31482 16712 31878
rect 16672 31476 16724 31482
rect 16672 31418 16724 31424
rect 16776 31346 16804 32846
rect 16856 31748 16908 31754
rect 16856 31690 16908 31696
rect 16764 31340 16816 31346
rect 16764 31282 16816 31288
rect 16580 31204 16632 31210
rect 16580 31146 16632 31152
rect 16304 30796 16356 30802
rect 16304 30738 16356 30744
rect 16316 30258 16344 30738
rect 16304 30252 16356 30258
rect 16304 30194 16356 30200
rect 16028 28756 16080 28762
rect 16028 28698 16080 28704
rect 15660 28484 15712 28490
rect 15660 28426 15712 28432
rect 15752 28484 15804 28490
rect 15752 28426 15804 28432
rect 15672 27674 15700 28426
rect 15660 27668 15712 27674
rect 15660 27610 15712 27616
rect 15764 27554 15792 28426
rect 15672 27526 15792 27554
rect 15844 27532 15896 27538
rect 15476 26444 15528 26450
rect 15476 26386 15528 26392
rect 15488 25362 15516 26386
rect 15476 25356 15528 25362
rect 15476 25298 15528 25304
rect 15292 20256 15344 20262
rect 15292 20198 15344 20204
rect 15200 20052 15252 20058
rect 15200 19994 15252 20000
rect 15304 19854 15332 20198
rect 15488 19922 15516 25298
rect 15672 20466 15700 27526
rect 15844 27474 15896 27480
rect 15752 26308 15804 26314
rect 15752 26250 15804 26256
rect 15764 24614 15792 26250
rect 15752 24608 15804 24614
rect 15752 24550 15804 24556
rect 15752 22976 15804 22982
rect 15752 22918 15804 22924
rect 15764 22710 15792 22918
rect 15752 22704 15804 22710
rect 15752 22646 15804 22652
rect 15856 22094 15884 27474
rect 16040 27470 16068 28698
rect 16028 27464 16080 27470
rect 16028 27406 16080 27412
rect 16304 27464 16356 27470
rect 16304 27406 16356 27412
rect 16316 27130 16344 27406
rect 16304 27124 16356 27130
rect 16304 27066 16356 27072
rect 15936 26988 15988 26994
rect 15936 26930 15988 26936
rect 15948 26586 15976 26930
rect 15936 26580 15988 26586
rect 15936 26522 15988 26528
rect 16488 26036 16540 26042
rect 16488 25978 16540 25984
rect 16120 25900 16172 25906
rect 16120 25842 16172 25848
rect 16132 25498 16160 25842
rect 16120 25492 16172 25498
rect 16120 25434 16172 25440
rect 16500 25294 16528 25978
rect 16488 25288 16540 25294
rect 16488 25230 16540 25236
rect 16592 23798 16620 31146
rect 16672 31136 16724 31142
rect 16672 31078 16724 31084
rect 16684 30734 16712 31078
rect 16672 30728 16724 30734
rect 16672 30670 16724 30676
rect 16684 30326 16712 30670
rect 16868 30326 16896 31690
rect 16672 30320 16724 30326
rect 16672 30262 16724 30268
rect 16856 30320 16908 30326
rect 16856 30262 16908 30268
rect 16684 29850 16712 30262
rect 16856 30048 16908 30054
rect 16856 29990 16908 29996
rect 16672 29844 16724 29850
rect 16672 29786 16724 29792
rect 16868 29646 16896 29990
rect 16856 29640 16908 29646
rect 16856 29582 16908 29588
rect 16764 28416 16816 28422
rect 16764 28358 16816 28364
rect 16776 28082 16804 28358
rect 16764 28076 16816 28082
rect 16764 28018 16816 28024
rect 16960 27010 16988 37606
rect 17052 36174 17080 39782
rect 17236 39302 17264 39986
rect 17316 39908 17368 39914
rect 17316 39850 17368 39856
rect 17328 39642 17356 39850
rect 17316 39636 17368 39642
rect 17316 39578 17368 39584
rect 17224 39296 17276 39302
rect 17224 39238 17276 39244
rect 17512 38434 17540 39986
rect 17880 39370 17908 40054
rect 18248 39846 18276 40394
rect 18616 40186 18644 40462
rect 18696 40384 18748 40390
rect 18696 40326 18748 40332
rect 18604 40180 18656 40186
rect 18604 40122 18656 40128
rect 18236 39840 18288 39846
rect 18236 39782 18288 39788
rect 18248 39574 18276 39782
rect 18315 39740 18623 39749
rect 18315 39738 18321 39740
rect 18377 39738 18401 39740
rect 18457 39738 18481 39740
rect 18537 39738 18561 39740
rect 18617 39738 18623 39740
rect 18377 39686 18379 39738
rect 18559 39686 18561 39738
rect 18315 39684 18321 39686
rect 18377 39684 18401 39686
rect 18457 39684 18481 39686
rect 18537 39684 18561 39686
rect 18617 39684 18623 39686
rect 18315 39675 18623 39684
rect 18708 39574 18736 40326
rect 19248 40180 19300 40186
rect 19248 40122 19300 40128
rect 18880 40044 18932 40050
rect 18880 39986 18932 39992
rect 18892 39574 18920 39986
rect 19260 39846 19288 40122
rect 19616 40044 19668 40050
rect 19616 39986 19668 39992
rect 19248 39840 19300 39846
rect 19248 39782 19300 39788
rect 18236 39568 18288 39574
rect 18236 39510 18288 39516
rect 18696 39568 18748 39574
rect 18696 39510 18748 39516
rect 18880 39568 18932 39574
rect 18880 39510 18932 39516
rect 17868 39364 17920 39370
rect 17868 39306 17920 39312
rect 17328 38406 17632 38434
rect 17328 38350 17356 38406
rect 17604 38350 17632 38406
rect 17316 38344 17368 38350
rect 17316 38286 17368 38292
rect 17592 38344 17644 38350
rect 17592 38286 17644 38292
rect 17132 38208 17184 38214
rect 17132 38150 17184 38156
rect 17144 37738 17172 38150
rect 17316 37868 17368 37874
rect 17316 37810 17368 37816
rect 17132 37732 17184 37738
rect 17132 37674 17184 37680
rect 17144 37466 17172 37674
rect 17328 37466 17356 37810
rect 17592 37664 17644 37670
rect 17592 37606 17644 37612
rect 17132 37460 17184 37466
rect 17132 37402 17184 37408
rect 17316 37460 17368 37466
rect 17316 37402 17368 37408
rect 17604 37194 17632 37606
rect 17592 37188 17644 37194
rect 17592 37130 17644 37136
rect 17040 36168 17092 36174
rect 17040 36110 17092 36116
rect 17316 36032 17368 36038
rect 17316 35974 17368 35980
rect 17132 35488 17184 35494
rect 17132 35430 17184 35436
rect 17144 35086 17172 35430
rect 17132 35080 17184 35086
rect 17132 35022 17184 35028
rect 17040 35012 17092 35018
rect 17040 34954 17092 34960
rect 17052 34610 17080 34954
rect 17328 34610 17356 35974
rect 17880 34746 17908 39306
rect 18144 39296 18196 39302
rect 18144 39238 18196 39244
rect 18052 39024 18104 39030
rect 18052 38966 18104 38972
rect 17960 38344 18012 38350
rect 17960 38286 18012 38292
rect 17972 38214 18000 38286
rect 18064 38282 18092 38966
rect 18052 38276 18104 38282
rect 18052 38218 18104 38224
rect 17960 38208 18012 38214
rect 17960 38150 18012 38156
rect 17972 36922 18000 38150
rect 18156 37448 18184 39238
rect 18248 38962 18276 39510
rect 18892 39438 18920 39510
rect 19260 39506 19288 39782
rect 19248 39500 19300 39506
rect 19248 39442 19300 39448
rect 18604 39432 18656 39438
rect 18604 39374 18656 39380
rect 18696 39432 18748 39438
rect 18696 39374 18748 39380
rect 18880 39432 18932 39438
rect 18880 39374 18932 39380
rect 18616 39098 18644 39374
rect 18604 39092 18656 39098
rect 18604 39034 18656 39040
rect 18708 39030 18736 39374
rect 19248 39296 19300 39302
rect 19248 39238 19300 39244
rect 18696 39024 18748 39030
rect 18696 38966 18748 38972
rect 18236 38956 18288 38962
rect 18236 38898 18288 38904
rect 18248 37874 18276 38898
rect 18788 38752 18840 38758
rect 18788 38694 18840 38700
rect 18315 38652 18623 38661
rect 18315 38650 18321 38652
rect 18377 38650 18401 38652
rect 18457 38650 18481 38652
rect 18537 38650 18561 38652
rect 18617 38650 18623 38652
rect 18377 38598 18379 38650
rect 18559 38598 18561 38650
rect 18315 38596 18321 38598
rect 18377 38596 18401 38598
rect 18457 38596 18481 38598
rect 18537 38596 18561 38598
rect 18617 38596 18623 38598
rect 18315 38587 18623 38596
rect 18800 38298 18828 38694
rect 18524 38270 18828 38298
rect 18420 38208 18472 38214
rect 18420 38150 18472 38156
rect 18432 37874 18460 38150
rect 18236 37868 18288 37874
rect 18236 37810 18288 37816
rect 18420 37868 18472 37874
rect 18420 37810 18472 37816
rect 18248 37670 18276 37810
rect 18524 37806 18552 38270
rect 18696 37868 18748 37874
rect 18696 37810 18748 37816
rect 18512 37800 18564 37806
rect 18512 37742 18564 37748
rect 18236 37664 18288 37670
rect 18236 37606 18288 37612
rect 18315 37564 18623 37573
rect 18315 37562 18321 37564
rect 18377 37562 18401 37564
rect 18457 37562 18481 37564
rect 18537 37562 18561 37564
rect 18617 37562 18623 37564
rect 18377 37510 18379 37562
rect 18559 37510 18561 37562
rect 18315 37508 18321 37510
rect 18377 37508 18401 37510
rect 18457 37508 18481 37510
rect 18537 37508 18561 37510
rect 18617 37508 18623 37510
rect 18315 37499 18623 37508
rect 18708 37466 18736 37810
rect 19156 37664 19208 37670
rect 19156 37606 19208 37612
rect 18696 37460 18748 37466
rect 18156 37420 18368 37448
rect 18340 37262 18368 37420
rect 18696 37402 18748 37408
rect 18144 37256 18196 37262
rect 18144 37198 18196 37204
rect 18328 37256 18380 37262
rect 18328 37198 18380 37204
rect 17960 36916 18012 36922
rect 17960 36858 18012 36864
rect 17972 35290 18000 36858
rect 18156 36242 18184 37198
rect 18236 37120 18288 37126
rect 18236 37062 18288 37068
rect 19064 37120 19116 37126
rect 19064 37062 19116 37068
rect 18144 36236 18196 36242
rect 18144 36178 18196 36184
rect 18248 35698 18276 37062
rect 19076 36786 19104 37062
rect 19064 36780 19116 36786
rect 19064 36722 19116 36728
rect 18315 36476 18623 36485
rect 18315 36474 18321 36476
rect 18377 36474 18401 36476
rect 18457 36474 18481 36476
rect 18537 36474 18561 36476
rect 18617 36474 18623 36476
rect 18377 36422 18379 36474
rect 18559 36422 18561 36474
rect 18315 36420 18321 36422
rect 18377 36420 18401 36422
rect 18457 36420 18481 36422
rect 18537 36420 18561 36422
rect 18617 36420 18623 36422
rect 18315 36411 18623 36420
rect 19076 36242 19104 36722
rect 19064 36236 19116 36242
rect 19064 36178 19116 36184
rect 18788 35760 18840 35766
rect 18788 35702 18840 35708
rect 18236 35692 18288 35698
rect 18236 35634 18288 35640
rect 18315 35388 18623 35397
rect 18315 35386 18321 35388
rect 18377 35386 18401 35388
rect 18457 35386 18481 35388
rect 18537 35386 18561 35388
rect 18617 35386 18623 35388
rect 18377 35334 18379 35386
rect 18559 35334 18561 35386
rect 18315 35332 18321 35334
rect 18377 35332 18401 35334
rect 18457 35332 18481 35334
rect 18537 35332 18561 35334
rect 18617 35332 18623 35334
rect 18315 35323 18623 35332
rect 17960 35284 18012 35290
rect 17960 35226 18012 35232
rect 18800 35086 18828 35702
rect 19168 35562 19196 37606
rect 19260 36786 19288 39238
rect 19628 38962 19656 39986
rect 20904 39976 20956 39982
rect 20904 39918 20956 39924
rect 20916 39438 20944 39918
rect 19800 39432 19852 39438
rect 19800 39374 19852 39380
rect 20260 39432 20312 39438
rect 20260 39374 20312 39380
rect 20904 39432 20956 39438
rect 20904 39374 20956 39380
rect 19812 39098 19840 39374
rect 19984 39296 20036 39302
rect 19984 39238 20036 39244
rect 19800 39092 19852 39098
rect 19800 39034 19852 39040
rect 19616 38956 19668 38962
rect 19616 38898 19668 38904
rect 19524 37868 19576 37874
rect 19524 37810 19576 37816
rect 19248 36780 19300 36786
rect 19248 36722 19300 36728
rect 19536 36666 19564 37810
rect 19616 37664 19668 37670
rect 19616 37606 19668 37612
rect 19444 36638 19564 36666
rect 19156 35556 19208 35562
rect 19156 35498 19208 35504
rect 18788 35080 18840 35086
rect 18788 35022 18840 35028
rect 17868 34740 17920 34746
rect 17868 34682 17920 34688
rect 17040 34604 17092 34610
rect 17040 34546 17092 34552
rect 17316 34604 17368 34610
rect 17316 34546 17368 34552
rect 18315 34300 18623 34309
rect 18315 34298 18321 34300
rect 18377 34298 18401 34300
rect 18457 34298 18481 34300
rect 18537 34298 18561 34300
rect 18617 34298 18623 34300
rect 18377 34246 18379 34298
rect 18559 34246 18561 34298
rect 18315 34244 18321 34246
rect 18377 34244 18401 34246
rect 18457 34244 18481 34246
rect 18537 34244 18561 34246
rect 18617 34244 18623 34246
rect 18315 34235 18623 34244
rect 18800 33454 18828 35022
rect 18788 33448 18840 33454
rect 18788 33390 18840 33396
rect 18315 33212 18623 33221
rect 18315 33210 18321 33212
rect 18377 33210 18401 33212
rect 18457 33210 18481 33212
rect 18537 33210 18561 33212
rect 18617 33210 18623 33212
rect 18377 33158 18379 33210
rect 18559 33158 18561 33210
rect 18315 33156 18321 33158
rect 18377 33156 18401 33158
rect 18457 33156 18481 33158
rect 18537 33156 18561 33158
rect 18617 33156 18623 33158
rect 18315 33147 18623 33156
rect 17040 32836 17092 32842
rect 17040 32778 17092 32784
rect 17052 31822 17080 32778
rect 17592 32428 17644 32434
rect 17592 32370 17644 32376
rect 17604 31822 17632 32370
rect 18800 32314 18828 33390
rect 18880 32768 18932 32774
rect 18880 32710 18932 32716
rect 18892 32434 18920 32710
rect 18880 32428 18932 32434
rect 18880 32370 18932 32376
rect 18800 32298 18920 32314
rect 18800 32292 18932 32298
rect 18800 32286 18880 32292
rect 18880 32234 18932 32240
rect 18315 32124 18623 32133
rect 18315 32122 18321 32124
rect 18377 32122 18401 32124
rect 18457 32122 18481 32124
rect 18537 32122 18561 32124
rect 18617 32122 18623 32124
rect 18377 32070 18379 32122
rect 18559 32070 18561 32122
rect 18315 32068 18321 32070
rect 18377 32068 18401 32070
rect 18457 32068 18481 32070
rect 18537 32068 18561 32070
rect 18617 32068 18623 32070
rect 18315 32059 18623 32068
rect 18604 31884 18656 31890
rect 18604 31826 18656 31832
rect 17040 31816 17092 31822
rect 17040 31758 17092 31764
rect 17592 31816 17644 31822
rect 17592 31758 17644 31764
rect 17052 30258 17080 31758
rect 17224 31340 17276 31346
rect 17224 31282 17276 31288
rect 17236 30598 17264 31282
rect 17224 30592 17276 30598
rect 17224 30534 17276 30540
rect 17236 30258 17264 30534
rect 17040 30252 17092 30258
rect 17224 30252 17276 30258
rect 17092 30212 17172 30240
rect 17040 30194 17092 30200
rect 17040 28484 17092 28490
rect 17040 28426 17092 28432
rect 17052 28218 17080 28426
rect 17040 28212 17092 28218
rect 17040 28154 17092 28160
rect 17144 27418 17172 30212
rect 17224 30194 17276 30200
rect 17500 30252 17552 30258
rect 17500 30194 17552 30200
rect 17512 29850 17540 30194
rect 17500 29844 17552 29850
rect 17500 29786 17552 29792
rect 17604 29714 17632 31758
rect 18616 31414 18644 31826
rect 18604 31408 18656 31414
rect 18604 31350 18656 31356
rect 18892 31278 18920 32234
rect 19444 32026 19472 36638
rect 19524 36576 19576 36582
rect 19524 36518 19576 36524
rect 19536 35086 19564 36518
rect 19628 36378 19656 37606
rect 19996 36922 20024 39238
rect 20076 37800 20128 37806
rect 20076 37742 20128 37748
rect 20088 37466 20116 37742
rect 20076 37460 20128 37466
rect 20076 37402 20128 37408
rect 20168 37256 20220 37262
rect 20168 37198 20220 37204
rect 19984 36916 20036 36922
rect 19984 36858 20036 36864
rect 19616 36372 19668 36378
rect 19616 36314 19668 36320
rect 19800 36100 19852 36106
rect 19800 36042 19852 36048
rect 19524 35080 19576 35086
rect 19524 35022 19576 35028
rect 19432 32020 19484 32026
rect 19432 31962 19484 31968
rect 19812 31754 19840 36042
rect 19996 32842 20024 36858
rect 20180 36242 20208 37198
rect 20272 36854 20300 39374
rect 20628 39296 20680 39302
rect 20628 39238 20680 39244
rect 20444 38888 20496 38894
rect 20444 38830 20496 38836
rect 20456 37466 20484 38830
rect 20444 37460 20496 37466
rect 20444 37402 20496 37408
rect 20536 37324 20588 37330
rect 20536 37266 20588 37272
rect 20444 37256 20496 37262
rect 20444 37198 20496 37204
rect 20456 36854 20484 37198
rect 20260 36848 20312 36854
rect 20260 36790 20312 36796
rect 20444 36848 20496 36854
rect 20444 36790 20496 36796
rect 20168 36236 20220 36242
rect 20168 36178 20220 36184
rect 20076 34604 20128 34610
rect 20076 34546 20128 34552
rect 19984 32836 20036 32842
rect 19984 32778 20036 32784
rect 20088 32450 20116 34546
rect 20168 32904 20220 32910
rect 20168 32846 20220 32852
rect 20180 32570 20208 32846
rect 20272 32842 20300 36790
rect 20352 36712 20404 36718
rect 20456 36700 20484 36790
rect 20404 36672 20484 36700
rect 20352 36654 20404 36660
rect 20352 36168 20404 36174
rect 20352 36110 20404 36116
rect 20364 34202 20392 36110
rect 20456 36106 20484 36672
rect 20444 36100 20496 36106
rect 20444 36042 20496 36048
rect 20548 35018 20576 37266
rect 20640 37262 20668 39238
rect 20916 38962 20944 39374
rect 20904 38956 20956 38962
rect 20904 38898 20956 38904
rect 20720 37460 20772 37466
rect 20720 37402 20772 37408
rect 20628 37256 20680 37262
rect 20628 37198 20680 37204
rect 20628 36916 20680 36922
rect 20628 36858 20680 36864
rect 20640 36786 20668 36858
rect 20628 36780 20680 36786
rect 20628 36722 20680 36728
rect 20732 36718 20760 37402
rect 20812 37256 20864 37262
rect 20812 37198 20864 37204
rect 20824 36922 20852 37198
rect 20812 36916 20864 36922
rect 20812 36858 20864 36864
rect 20720 36712 20772 36718
rect 20720 36654 20772 36660
rect 20536 35012 20588 35018
rect 20536 34954 20588 34960
rect 20732 34542 20760 36654
rect 20812 36644 20864 36650
rect 20812 36586 20864 36592
rect 20824 36378 20852 36586
rect 20812 36372 20864 36378
rect 20812 36314 20864 36320
rect 20812 36168 20864 36174
rect 20812 36110 20864 36116
rect 20720 34536 20772 34542
rect 20720 34478 20772 34484
rect 20720 34400 20772 34406
rect 20720 34342 20772 34348
rect 20352 34196 20404 34202
rect 20352 34138 20404 34144
rect 20364 32910 20392 34138
rect 20732 33998 20760 34342
rect 20720 33992 20772 33998
rect 20720 33934 20772 33940
rect 20352 32904 20404 32910
rect 20352 32846 20404 32852
rect 20260 32836 20312 32842
rect 20260 32778 20312 32784
rect 20168 32564 20220 32570
rect 20168 32506 20220 32512
rect 20088 32422 20208 32450
rect 19892 31816 19944 31822
rect 19892 31758 19944 31764
rect 20076 31816 20128 31822
rect 20076 31758 20128 31764
rect 19616 31748 19840 31754
rect 19668 31726 19840 31748
rect 19616 31690 19668 31696
rect 18880 31272 18932 31278
rect 18880 31214 18932 31220
rect 18315 31036 18623 31045
rect 18315 31034 18321 31036
rect 18377 31034 18401 31036
rect 18457 31034 18481 31036
rect 18537 31034 18561 31036
rect 18617 31034 18623 31036
rect 18377 30982 18379 31034
rect 18559 30982 18561 31034
rect 18315 30980 18321 30982
rect 18377 30980 18401 30982
rect 18457 30980 18481 30982
rect 18537 30980 18561 30982
rect 18617 30980 18623 30982
rect 18315 30971 18623 30980
rect 18315 29948 18623 29957
rect 18315 29946 18321 29948
rect 18377 29946 18401 29948
rect 18457 29946 18481 29948
rect 18537 29946 18561 29948
rect 18617 29946 18623 29948
rect 18377 29894 18379 29946
rect 18559 29894 18561 29946
rect 18315 29892 18321 29894
rect 18377 29892 18401 29894
rect 18457 29892 18481 29894
rect 18537 29892 18561 29894
rect 18617 29892 18623 29894
rect 18315 29883 18623 29892
rect 17776 29844 17828 29850
rect 17776 29786 17828 29792
rect 17592 29708 17644 29714
rect 17592 29650 17644 29656
rect 17144 27390 17264 27418
rect 17132 27328 17184 27334
rect 17132 27270 17184 27276
rect 16684 26982 16988 27010
rect 17144 26994 17172 27270
rect 17132 26988 17184 26994
rect 16580 23792 16632 23798
rect 16580 23734 16632 23740
rect 16396 23520 16448 23526
rect 16396 23462 16448 23468
rect 16408 23118 16436 23462
rect 16592 23118 16620 23734
rect 16396 23112 16448 23118
rect 16396 23054 16448 23060
rect 16580 23112 16632 23118
rect 16580 23054 16632 23060
rect 16212 23044 16264 23050
rect 16212 22986 16264 22992
rect 15856 22066 15976 22094
rect 15660 20460 15712 20466
rect 15660 20402 15712 20408
rect 15844 20460 15896 20466
rect 15844 20402 15896 20408
rect 15476 19916 15528 19922
rect 15476 19858 15528 19864
rect 15292 19848 15344 19854
rect 15292 19790 15344 19796
rect 14372 19780 14424 19786
rect 14372 19722 14424 19728
rect 14842 19612 15150 19621
rect 14842 19610 14848 19612
rect 14904 19610 14928 19612
rect 14984 19610 15008 19612
rect 15064 19610 15088 19612
rect 15144 19610 15150 19612
rect 14904 19558 14906 19610
rect 15086 19558 15088 19610
rect 14842 19556 14848 19558
rect 14904 19556 14928 19558
rect 14984 19556 15008 19558
rect 15064 19556 15088 19558
rect 15144 19556 15150 19558
rect 14842 19547 15150 19556
rect 14842 18524 15150 18533
rect 14842 18522 14848 18524
rect 14904 18522 14928 18524
rect 14984 18522 15008 18524
rect 15064 18522 15088 18524
rect 15144 18522 15150 18524
rect 14904 18470 14906 18522
rect 15086 18470 15088 18522
rect 14842 18468 14848 18470
rect 14904 18468 14928 18470
rect 14984 18468 15008 18470
rect 15064 18468 15088 18470
rect 15144 18468 15150 18470
rect 14842 18459 15150 18468
rect 14842 17436 15150 17445
rect 14842 17434 14848 17436
rect 14904 17434 14928 17436
rect 14984 17434 15008 17436
rect 15064 17434 15088 17436
rect 15144 17434 15150 17436
rect 14904 17382 14906 17434
rect 15086 17382 15088 17434
rect 14842 17380 14848 17382
rect 14904 17380 14928 17382
rect 14984 17380 15008 17382
rect 15064 17380 15088 17382
rect 15144 17380 15150 17382
rect 14842 17371 15150 17380
rect 15488 17270 15516 19858
rect 15660 19712 15712 19718
rect 15660 19654 15712 19660
rect 15672 18630 15700 19654
rect 15660 18624 15712 18630
rect 15660 18566 15712 18572
rect 15856 18290 15884 20402
rect 15660 18284 15712 18290
rect 15660 18226 15712 18232
rect 15844 18284 15896 18290
rect 15844 18226 15896 18232
rect 15672 17882 15700 18226
rect 15660 17876 15712 17882
rect 15660 17818 15712 17824
rect 15948 17746 15976 22066
rect 16120 21888 16172 21894
rect 16120 21830 16172 21836
rect 16132 21622 16160 21830
rect 16224 21690 16252 22986
rect 16212 21684 16264 21690
rect 16212 21626 16264 21632
rect 16120 21616 16172 21622
rect 16120 21558 16172 21564
rect 16028 20936 16080 20942
rect 16028 20878 16080 20884
rect 16040 20602 16068 20878
rect 16028 20596 16080 20602
rect 16028 20538 16080 20544
rect 16120 19372 16172 19378
rect 16224 19360 16252 21626
rect 16684 19514 16712 26982
rect 17132 26930 17184 26936
rect 16764 26920 16816 26926
rect 16764 26862 16816 26868
rect 16856 26920 16908 26926
rect 16856 26862 16908 26868
rect 16776 25226 16804 26862
rect 16868 25838 16896 26862
rect 16856 25832 16908 25838
rect 16856 25774 16908 25780
rect 16764 25220 16816 25226
rect 16764 25162 16816 25168
rect 16868 24818 16896 25774
rect 17132 25220 17184 25226
rect 17132 25162 17184 25168
rect 16856 24812 16908 24818
rect 16856 24754 16908 24760
rect 17144 24206 17172 25162
rect 17132 24200 17184 24206
rect 17132 24142 17184 24148
rect 17040 23112 17092 23118
rect 17040 23054 17092 23060
rect 17052 22778 17080 23054
rect 17040 22772 17092 22778
rect 17040 22714 17092 22720
rect 17052 22642 17080 22714
rect 17040 22636 17092 22642
rect 17040 22578 17092 22584
rect 16856 22432 16908 22438
rect 16856 22374 16908 22380
rect 16868 22030 16896 22374
rect 17144 22098 17172 24142
rect 17236 23186 17264 27390
rect 17788 27282 17816 29786
rect 18892 29646 18920 31214
rect 19340 30728 19392 30734
rect 19340 30670 19392 30676
rect 19352 30394 19380 30670
rect 19340 30388 19392 30394
rect 19340 30330 19392 30336
rect 18880 29640 18932 29646
rect 18880 29582 18932 29588
rect 18892 28966 18920 29582
rect 18880 28960 18932 28966
rect 18880 28902 18932 28908
rect 18315 28860 18623 28869
rect 18315 28858 18321 28860
rect 18377 28858 18401 28860
rect 18457 28858 18481 28860
rect 18537 28858 18561 28860
rect 18617 28858 18623 28860
rect 18377 28806 18379 28858
rect 18559 28806 18561 28858
rect 18315 28804 18321 28806
rect 18377 28804 18401 28806
rect 18457 28804 18481 28806
rect 18537 28804 18561 28806
rect 18617 28804 18623 28806
rect 18315 28795 18623 28804
rect 18892 28558 18920 28902
rect 18880 28552 18932 28558
rect 18880 28494 18932 28500
rect 18315 27772 18623 27781
rect 18315 27770 18321 27772
rect 18377 27770 18401 27772
rect 18457 27770 18481 27772
rect 18537 27770 18561 27772
rect 18617 27770 18623 27772
rect 18377 27718 18379 27770
rect 18559 27718 18561 27770
rect 18315 27716 18321 27718
rect 18377 27716 18401 27718
rect 18457 27716 18481 27718
rect 18537 27716 18561 27718
rect 18617 27716 18623 27718
rect 18315 27707 18623 27716
rect 18892 27470 18920 28494
rect 19352 28422 19380 30330
rect 19524 30048 19576 30054
rect 19524 29990 19576 29996
rect 19536 29646 19564 29990
rect 19524 29640 19576 29646
rect 19524 29582 19576 29588
rect 19340 28416 19392 28422
rect 19340 28358 19392 28364
rect 19352 28082 19380 28358
rect 19340 28076 19392 28082
rect 19340 28018 19392 28024
rect 18880 27464 18932 27470
rect 18880 27406 18932 27412
rect 17788 27254 17908 27282
rect 17500 24812 17552 24818
rect 17500 24754 17552 24760
rect 17512 24410 17540 24754
rect 17500 24404 17552 24410
rect 17500 24346 17552 24352
rect 17316 24200 17368 24206
rect 17316 24142 17368 24148
rect 17328 23322 17356 24142
rect 17592 23588 17644 23594
rect 17592 23530 17644 23536
rect 17316 23316 17368 23322
rect 17316 23258 17368 23264
rect 17224 23180 17276 23186
rect 17224 23122 17276 23128
rect 17604 23118 17632 23530
rect 17684 23520 17736 23526
rect 17684 23462 17736 23468
rect 17696 23186 17724 23462
rect 17684 23180 17736 23186
rect 17684 23122 17736 23128
rect 17592 23112 17644 23118
rect 17592 23054 17644 23060
rect 17224 23044 17276 23050
rect 17224 22986 17276 22992
rect 17236 22642 17264 22986
rect 17224 22636 17276 22642
rect 17224 22578 17276 22584
rect 17316 22568 17368 22574
rect 17316 22510 17368 22516
rect 17132 22092 17184 22098
rect 17328 22094 17356 22510
rect 17132 22034 17184 22040
rect 17236 22066 17356 22094
rect 16856 22024 16908 22030
rect 16856 21966 16908 21972
rect 16948 20800 17000 20806
rect 16948 20742 17000 20748
rect 16960 20466 16988 20742
rect 16948 20460 17000 20466
rect 16948 20402 17000 20408
rect 16672 19508 16724 19514
rect 16672 19450 16724 19456
rect 17236 19446 17264 22066
rect 17224 19440 17276 19446
rect 17224 19382 17276 19388
rect 16172 19332 16252 19360
rect 16120 19314 16172 19320
rect 16224 18222 16252 19332
rect 16856 19372 16908 19378
rect 16856 19314 16908 19320
rect 16868 18426 16896 19314
rect 17236 18766 17264 19382
rect 17408 19372 17460 19378
rect 17408 19314 17460 19320
rect 17224 18760 17276 18766
rect 17224 18702 17276 18708
rect 17224 18624 17276 18630
rect 17224 18566 17276 18572
rect 17236 18426 17264 18566
rect 16856 18420 16908 18426
rect 16856 18362 16908 18368
rect 17224 18420 17276 18426
rect 17224 18362 17276 18368
rect 17132 18284 17184 18290
rect 17132 18226 17184 18232
rect 16212 18216 16264 18222
rect 16212 18158 16264 18164
rect 16856 18080 16908 18086
rect 16856 18022 16908 18028
rect 15936 17740 15988 17746
rect 15936 17682 15988 17688
rect 15476 17264 15528 17270
rect 15476 17206 15528 17212
rect 15844 17196 15896 17202
rect 15948 17184 15976 17682
rect 16868 17202 16896 18022
rect 17144 17882 17172 18226
rect 17132 17876 17184 17882
rect 17132 17818 17184 17824
rect 17236 17746 17264 18362
rect 17316 18284 17368 18290
rect 17316 18226 17368 18232
rect 17224 17740 17276 17746
rect 17224 17682 17276 17688
rect 17328 17610 17356 18226
rect 17420 17882 17448 19314
rect 17696 18850 17724 23122
rect 17880 23118 17908 27254
rect 18892 26994 18920 27406
rect 18880 26988 18932 26994
rect 18880 26930 18932 26936
rect 18972 26988 19024 26994
rect 18972 26930 19024 26936
rect 18236 26784 18288 26790
rect 18236 26726 18288 26732
rect 18248 26382 18276 26726
rect 18315 26684 18623 26693
rect 18315 26682 18321 26684
rect 18377 26682 18401 26684
rect 18457 26682 18481 26684
rect 18537 26682 18561 26684
rect 18617 26682 18623 26684
rect 18377 26630 18379 26682
rect 18559 26630 18561 26682
rect 18315 26628 18321 26630
rect 18377 26628 18401 26630
rect 18457 26628 18481 26630
rect 18537 26628 18561 26630
rect 18617 26628 18623 26630
rect 18315 26619 18623 26628
rect 18892 26450 18920 26930
rect 18880 26444 18932 26450
rect 18880 26386 18932 26392
rect 18236 26376 18288 26382
rect 18236 26318 18288 26324
rect 18315 25596 18623 25605
rect 18315 25594 18321 25596
rect 18377 25594 18401 25596
rect 18457 25594 18481 25596
rect 18537 25594 18561 25596
rect 18617 25594 18623 25596
rect 18377 25542 18379 25594
rect 18559 25542 18561 25594
rect 18315 25540 18321 25542
rect 18377 25540 18401 25542
rect 18457 25540 18481 25542
rect 18537 25540 18561 25542
rect 18617 25540 18623 25542
rect 18315 25531 18623 25540
rect 18984 25498 19012 26930
rect 19628 26790 19656 31690
rect 19904 31226 19932 31758
rect 19720 31198 19932 31226
rect 19616 26784 19668 26790
rect 19616 26726 19668 26732
rect 19720 26042 19748 31198
rect 20088 31142 20116 31758
rect 19892 31136 19944 31142
rect 19892 31078 19944 31084
rect 20076 31136 20128 31142
rect 20076 31078 20128 31084
rect 19904 30326 19932 31078
rect 19892 30320 19944 30326
rect 19892 30262 19944 30268
rect 20076 30252 20128 30258
rect 20076 30194 20128 30200
rect 20088 29170 20116 30194
rect 20076 29164 20128 29170
rect 20076 29106 20128 29112
rect 19800 27396 19852 27402
rect 19800 27338 19852 27344
rect 19812 26586 19840 27338
rect 19800 26580 19852 26586
rect 19800 26522 19852 26528
rect 19984 26376 20036 26382
rect 19984 26318 20036 26324
rect 19996 26042 20024 26318
rect 19708 26036 19760 26042
rect 19708 25978 19760 25984
rect 19984 26036 20036 26042
rect 19984 25978 20036 25984
rect 19984 25900 20036 25906
rect 19984 25842 20036 25848
rect 18972 25492 19024 25498
rect 18972 25434 19024 25440
rect 18236 25288 18288 25294
rect 18236 25230 18288 25236
rect 17868 23112 17920 23118
rect 17868 23054 17920 23060
rect 17880 22794 17908 23054
rect 17788 22766 17908 22794
rect 18248 22778 18276 25230
rect 19996 24954 20024 25842
rect 19984 24948 20036 24954
rect 19984 24890 20036 24896
rect 18786 24712 18842 24721
rect 18786 24647 18788 24656
rect 18840 24647 18842 24656
rect 18788 24618 18840 24624
rect 18315 24508 18623 24517
rect 18315 24506 18321 24508
rect 18377 24506 18401 24508
rect 18457 24506 18481 24508
rect 18537 24506 18561 24508
rect 18617 24506 18623 24508
rect 18377 24454 18379 24506
rect 18559 24454 18561 24506
rect 18315 24452 18321 24454
rect 18377 24452 18401 24454
rect 18457 24452 18481 24454
rect 18537 24452 18561 24454
rect 18617 24452 18623 24454
rect 18315 24443 18623 24452
rect 18800 23746 18828 24618
rect 19892 24608 19944 24614
rect 19892 24550 19944 24556
rect 19432 24200 19484 24206
rect 19432 24142 19484 24148
rect 18708 23730 18828 23746
rect 18696 23724 18828 23730
rect 18748 23718 18828 23724
rect 18696 23666 18748 23672
rect 18315 23420 18623 23429
rect 18315 23418 18321 23420
rect 18377 23418 18401 23420
rect 18457 23418 18481 23420
rect 18537 23418 18561 23420
rect 18617 23418 18623 23420
rect 18377 23366 18379 23418
rect 18559 23366 18561 23418
rect 18315 23364 18321 23366
rect 18377 23364 18401 23366
rect 18457 23364 18481 23366
rect 18537 23364 18561 23366
rect 18617 23364 18623 23366
rect 18315 23355 18623 23364
rect 18708 23118 18736 23666
rect 18880 23520 18932 23526
rect 18880 23462 18932 23468
rect 18696 23112 18748 23118
rect 18696 23054 18748 23060
rect 18236 22772 18288 22778
rect 17788 22642 17816 22766
rect 18236 22714 18288 22720
rect 18892 22642 18920 23462
rect 17776 22636 17828 22642
rect 17776 22578 17828 22584
rect 18696 22636 18748 22642
rect 18696 22578 18748 22584
rect 18880 22636 18932 22642
rect 18880 22578 18932 22584
rect 18972 22636 19024 22642
rect 18972 22578 19024 22584
rect 18315 22332 18623 22341
rect 18315 22330 18321 22332
rect 18377 22330 18401 22332
rect 18457 22330 18481 22332
rect 18537 22330 18561 22332
rect 18617 22330 18623 22332
rect 18377 22278 18379 22330
rect 18559 22278 18561 22330
rect 18315 22276 18321 22278
rect 18377 22276 18401 22278
rect 18457 22276 18481 22278
rect 18537 22276 18561 22278
rect 18617 22276 18623 22278
rect 18315 22267 18623 22276
rect 18708 22234 18736 22578
rect 18984 22420 19012 22578
rect 19064 22432 19116 22438
rect 18984 22392 19064 22420
rect 19064 22374 19116 22380
rect 18696 22228 18748 22234
rect 18696 22170 18748 22176
rect 18236 22024 18288 22030
rect 18236 21966 18288 21972
rect 18248 21350 18276 21966
rect 18236 21344 18288 21350
rect 18236 21286 18288 21292
rect 18248 20534 18276 21286
rect 18315 21244 18623 21253
rect 18315 21242 18321 21244
rect 18377 21242 18401 21244
rect 18457 21242 18481 21244
rect 18537 21242 18561 21244
rect 18617 21242 18623 21244
rect 18377 21190 18379 21242
rect 18559 21190 18561 21242
rect 18315 21188 18321 21190
rect 18377 21188 18401 21190
rect 18457 21188 18481 21190
rect 18537 21188 18561 21190
rect 18617 21188 18623 21190
rect 18315 21179 18623 21188
rect 18236 20528 18288 20534
rect 18236 20470 18288 20476
rect 18144 19168 18196 19174
rect 18144 19110 18196 19116
rect 18052 18964 18104 18970
rect 18052 18906 18104 18912
rect 17696 18834 18000 18850
rect 17696 18828 18012 18834
rect 17696 18822 17960 18828
rect 17696 18766 17724 18822
rect 17960 18770 18012 18776
rect 18064 18766 18092 18906
rect 17684 18760 17736 18766
rect 17684 18702 17736 18708
rect 18052 18760 18104 18766
rect 18052 18702 18104 18708
rect 17500 18624 17552 18630
rect 17500 18566 17552 18572
rect 17512 18290 17540 18566
rect 17500 18284 17552 18290
rect 17500 18226 17552 18232
rect 17408 17876 17460 17882
rect 17408 17818 17460 17824
rect 17316 17604 17368 17610
rect 17316 17546 17368 17552
rect 17960 17536 18012 17542
rect 17960 17478 18012 17484
rect 17316 17264 17368 17270
rect 17316 17206 17368 17212
rect 15896 17156 15976 17184
rect 15844 17138 15896 17144
rect 13268 16788 13320 16794
rect 13268 16730 13320 16736
rect 13452 16584 13504 16590
rect 13452 16526 13504 16532
rect 13728 16584 13780 16590
rect 13728 16526 13780 16532
rect 12900 15496 12952 15502
rect 12900 15438 12952 15444
rect 12912 14958 12940 15438
rect 13464 15162 13492 16526
rect 13740 16250 13768 16526
rect 13820 16448 13872 16454
rect 13820 16390 13872 16396
rect 13728 16244 13780 16250
rect 13728 16186 13780 16192
rect 13832 15706 13860 16390
rect 14842 16348 15150 16357
rect 14842 16346 14848 16348
rect 14904 16346 14928 16348
rect 14984 16346 15008 16348
rect 15064 16346 15088 16348
rect 15144 16346 15150 16348
rect 14904 16294 14906 16346
rect 15086 16294 15088 16346
rect 14842 16292 14848 16294
rect 14904 16292 14928 16294
rect 14984 16292 15008 16294
rect 15064 16292 15088 16294
rect 15144 16292 15150 16294
rect 14842 16283 15150 16292
rect 14280 16108 14332 16114
rect 14280 16050 14332 16056
rect 15200 16108 15252 16114
rect 15200 16050 15252 16056
rect 15844 16108 15896 16114
rect 15844 16050 15896 16056
rect 14292 15994 14320 16050
rect 14292 15966 14412 15994
rect 13820 15700 13872 15706
rect 13820 15642 13872 15648
rect 13728 15496 13780 15502
rect 13728 15438 13780 15444
rect 13452 15156 13504 15162
rect 13452 15098 13504 15104
rect 13360 15020 13412 15026
rect 13360 14962 13412 14968
rect 12900 14952 12952 14958
rect 12900 14894 12952 14900
rect 12912 14482 12940 14894
rect 13084 14544 13136 14550
rect 13004 14492 13084 14498
rect 13004 14486 13136 14492
rect 12900 14476 12952 14482
rect 12900 14418 12952 14424
rect 13004 14470 13124 14486
rect 13004 14362 13032 14470
rect 13372 14414 13400 14962
rect 12912 14346 13032 14362
rect 13360 14408 13412 14414
rect 13360 14350 13412 14356
rect 12900 14340 13032 14346
rect 12952 14334 13032 14340
rect 12900 14282 12952 14288
rect 13464 14278 13492 15098
rect 13740 15094 13768 15438
rect 13728 15088 13780 15094
rect 13728 15030 13780 15036
rect 13832 14346 13860 15642
rect 14384 15502 14412 15966
rect 14648 15904 14700 15910
rect 14648 15846 14700 15852
rect 14660 15502 14688 15846
rect 14372 15496 14424 15502
rect 14372 15438 14424 15444
rect 14648 15496 14700 15502
rect 14648 15438 14700 15444
rect 14384 15162 14412 15438
rect 14372 15156 14424 15162
rect 14372 15098 14424 15104
rect 14280 15020 14332 15026
rect 14280 14962 14332 14968
rect 14292 14482 14320 14962
rect 14280 14476 14332 14482
rect 14280 14418 14332 14424
rect 13820 14340 13872 14346
rect 13820 14282 13872 14288
rect 13084 14272 13136 14278
rect 13084 14214 13136 14220
rect 13452 14272 13504 14278
rect 13452 14214 13504 14220
rect 13096 14074 13124 14214
rect 13084 14068 13136 14074
rect 13084 14010 13136 14016
rect 14384 13326 14412 15098
rect 14660 14890 14688 15438
rect 14842 15260 15150 15269
rect 14842 15258 14848 15260
rect 14904 15258 14928 15260
rect 14984 15258 15008 15260
rect 15064 15258 15088 15260
rect 15144 15258 15150 15260
rect 14904 15206 14906 15258
rect 15086 15206 15088 15258
rect 14842 15204 14848 15206
rect 14904 15204 14928 15206
rect 14984 15204 15008 15206
rect 15064 15204 15088 15206
rect 15144 15204 15150 15206
rect 14842 15195 15150 15204
rect 15212 14890 15240 16050
rect 15752 15700 15804 15706
rect 15752 15642 15804 15648
rect 15292 15496 15344 15502
rect 15292 15438 15344 15444
rect 14648 14884 14700 14890
rect 14648 14826 14700 14832
rect 15200 14884 15252 14890
rect 15200 14826 15252 14832
rect 14660 14498 14688 14826
rect 15304 14822 15332 15438
rect 15476 15360 15528 15366
rect 15476 15302 15528 15308
rect 14740 14816 14792 14822
rect 14740 14758 14792 14764
rect 15292 14816 15344 14822
rect 15292 14758 15344 14764
rect 14568 14470 14688 14498
rect 14464 13864 14516 13870
rect 14464 13806 14516 13812
rect 14476 13530 14504 13806
rect 14464 13524 14516 13530
rect 14464 13466 14516 13472
rect 14568 13326 14596 14470
rect 14648 14340 14700 14346
rect 14648 14282 14700 14288
rect 14660 13870 14688 14282
rect 14648 13864 14700 13870
rect 14648 13806 14700 13812
rect 14752 13326 14780 14758
rect 14832 14544 14884 14550
rect 14832 14486 14884 14492
rect 14844 14414 14872 14486
rect 14832 14408 14884 14414
rect 14832 14350 14884 14356
rect 14842 14172 15150 14181
rect 14842 14170 14848 14172
rect 14904 14170 14928 14172
rect 14984 14170 15008 14172
rect 15064 14170 15088 14172
rect 15144 14170 15150 14172
rect 14904 14118 14906 14170
rect 15086 14118 15088 14170
rect 14842 14116 14848 14118
rect 14904 14116 14928 14118
rect 14984 14116 15008 14118
rect 15064 14116 15088 14118
rect 15144 14116 15150 14118
rect 14842 14107 15150 14116
rect 15304 14074 15332 14758
rect 15488 14414 15516 15302
rect 15764 15162 15792 15642
rect 15752 15156 15804 15162
rect 15752 15098 15804 15104
rect 15568 14816 15620 14822
rect 15568 14758 15620 14764
rect 15580 14414 15608 14758
rect 15856 14414 15884 16050
rect 15476 14408 15528 14414
rect 15476 14350 15528 14356
rect 15568 14408 15620 14414
rect 15568 14350 15620 14356
rect 15844 14408 15896 14414
rect 15844 14350 15896 14356
rect 15292 14068 15344 14074
rect 15292 14010 15344 14016
rect 15016 13932 15068 13938
rect 15016 13874 15068 13880
rect 15108 13932 15160 13938
rect 15108 13874 15160 13880
rect 13544 13320 13596 13326
rect 13544 13262 13596 13268
rect 14372 13320 14424 13326
rect 14372 13262 14424 13268
rect 14556 13320 14608 13326
rect 14556 13262 14608 13268
rect 14740 13320 14792 13326
rect 14740 13262 14792 13268
rect 13556 10742 13584 13262
rect 15028 13258 15056 13874
rect 15120 13326 15148 13874
rect 15108 13320 15160 13326
rect 15108 13262 15160 13268
rect 15016 13252 15068 13258
rect 15016 13194 15068 13200
rect 14842 13084 15150 13093
rect 14842 13082 14848 13084
rect 14904 13082 14928 13084
rect 14984 13082 15008 13084
rect 15064 13082 15088 13084
rect 15144 13082 15150 13084
rect 14904 13030 14906 13082
rect 15086 13030 15088 13082
rect 14842 13028 14848 13030
rect 14904 13028 14928 13030
rect 14984 13028 15008 13030
rect 15064 13028 15088 13030
rect 15144 13028 15150 13030
rect 14842 13019 15150 13028
rect 14842 11996 15150 12005
rect 14842 11994 14848 11996
rect 14904 11994 14928 11996
rect 14984 11994 15008 11996
rect 15064 11994 15088 11996
rect 15144 11994 15150 11996
rect 14904 11942 14906 11994
rect 15086 11942 15088 11994
rect 14842 11940 14848 11942
rect 14904 11940 14928 11942
rect 14984 11940 15008 11942
rect 15064 11940 15088 11942
rect 15144 11940 15150 11942
rect 14842 11931 15150 11940
rect 14842 10908 15150 10917
rect 14842 10906 14848 10908
rect 14904 10906 14928 10908
rect 14984 10906 15008 10908
rect 15064 10906 15088 10908
rect 15144 10906 15150 10908
rect 14904 10854 14906 10906
rect 15086 10854 15088 10906
rect 14842 10852 14848 10854
rect 14904 10852 14928 10854
rect 14984 10852 15008 10854
rect 15064 10852 15088 10854
rect 15144 10852 15150 10854
rect 14842 10843 15150 10852
rect 13544 10736 13596 10742
rect 13544 10678 13596 10684
rect 12716 8560 12768 8566
rect 12716 8502 12768 8508
rect 11369 8188 11677 8197
rect 11369 8186 11375 8188
rect 11431 8186 11455 8188
rect 11511 8186 11535 8188
rect 11591 8186 11615 8188
rect 11671 8186 11677 8188
rect 11431 8134 11433 8186
rect 11613 8134 11615 8186
rect 11369 8132 11375 8134
rect 11431 8132 11455 8134
rect 11511 8132 11535 8134
rect 11591 8132 11615 8134
rect 11671 8132 11677 8134
rect 11369 8123 11677 8132
rect 11369 7100 11677 7109
rect 11369 7098 11375 7100
rect 11431 7098 11455 7100
rect 11511 7098 11535 7100
rect 11591 7098 11615 7100
rect 11671 7098 11677 7100
rect 11431 7046 11433 7098
rect 11613 7046 11615 7098
rect 11369 7044 11375 7046
rect 11431 7044 11455 7046
rect 11511 7044 11535 7046
rect 11591 7044 11615 7046
rect 11671 7044 11677 7046
rect 11369 7035 11677 7044
rect 11369 6012 11677 6021
rect 11369 6010 11375 6012
rect 11431 6010 11455 6012
rect 11511 6010 11535 6012
rect 11591 6010 11615 6012
rect 11671 6010 11677 6012
rect 11431 5958 11433 6010
rect 11613 5958 11615 6010
rect 11369 5956 11375 5958
rect 11431 5956 11455 5958
rect 11511 5956 11535 5958
rect 11591 5956 11615 5958
rect 11671 5956 11677 5958
rect 11369 5947 11677 5956
rect 10508 5296 10560 5302
rect 10508 5238 10560 5244
rect 10520 4146 10548 5238
rect 11369 4924 11677 4933
rect 11369 4922 11375 4924
rect 11431 4922 11455 4924
rect 11511 4922 11535 4924
rect 11591 4922 11615 4924
rect 11671 4922 11677 4924
rect 11431 4870 11433 4922
rect 11613 4870 11615 4922
rect 11369 4868 11375 4870
rect 11431 4868 11455 4870
rect 11511 4868 11535 4870
rect 11591 4868 11615 4870
rect 11671 4868 11677 4870
rect 11369 4859 11677 4868
rect 10508 4140 10560 4146
rect 10508 4082 10560 4088
rect 11796 4072 11848 4078
rect 11796 4014 11848 4020
rect 12808 4072 12860 4078
rect 12808 4014 12860 4020
rect 12992 4072 13044 4078
rect 12992 4014 13044 4020
rect 10600 3936 10652 3942
rect 10600 3878 10652 3884
rect 10612 3602 10640 3878
rect 11369 3836 11677 3845
rect 11369 3834 11375 3836
rect 11431 3834 11455 3836
rect 11511 3834 11535 3836
rect 11591 3834 11615 3836
rect 11671 3834 11677 3836
rect 11431 3782 11433 3834
rect 11613 3782 11615 3834
rect 11369 3780 11375 3782
rect 11431 3780 11455 3782
rect 11511 3780 11535 3782
rect 11591 3780 11615 3782
rect 11671 3780 11677 3782
rect 11369 3771 11677 3780
rect 11808 3602 11836 4014
rect 12820 3738 12848 4014
rect 12808 3732 12860 3738
rect 12808 3674 12860 3680
rect 10600 3596 10652 3602
rect 10600 3538 10652 3544
rect 10968 3596 11020 3602
rect 10968 3538 11020 3544
rect 11796 3596 11848 3602
rect 11796 3538 11848 3544
rect 9680 2984 9732 2990
rect 9680 2926 9732 2932
rect 9496 2508 9548 2514
rect 9496 2450 9548 2456
rect 9036 2440 9088 2446
rect 9036 2382 9088 2388
rect 9048 800 9076 2382
rect 9692 800 9720 2926
rect 10980 800 11008 3538
rect 13004 3194 13032 4014
rect 13556 3534 13584 10678
rect 14842 9820 15150 9829
rect 14842 9818 14848 9820
rect 14904 9818 14928 9820
rect 14984 9818 15008 9820
rect 15064 9818 15088 9820
rect 15144 9818 15150 9820
rect 14904 9766 14906 9818
rect 15086 9766 15088 9818
rect 14842 9764 14848 9766
rect 14904 9764 14928 9766
rect 14984 9764 15008 9766
rect 15064 9764 15088 9766
rect 15144 9764 15150 9766
rect 14842 9755 15150 9764
rect 14842 8732 15150 8741
rect 14842 8730 14848 8732
rect 14904 8730 14928 8732
rect 14984 8730 15008 8732
rect 15064 8730 15088 8732
rect 15144 8730 15150 8732
rect 14904 8678 14906 8730
rect 15086 8678 15088 8730
rect 14842 8676 14848 8678
rect 14904 8676 14928 8678
rect 14984 8676 15008 8678
rect 15064 8676 15088 8678
rect 15144 8676 15150 8678
rect 14842 8667 15150 8676
rect 14842 7644 15150 7653
rect 14842 7642 14848 7644
rect 14904 7642 14928 7644
rect 14984 7642 15008 7644
rect 15064 7642 15088 7644
rect 15144 7642 15150 7644
rect 14904 7590 14906 7642
rect 15086 7590 15088 7642
rect 14842 7588 14848 7590
rect 14904 7588 14928 7590
rect 14984 7588 15008 7590
rect 15064 7588 15088 7590
rect 15144 7588 15150 7590
rect 14842 7579 15150 7588
rect 15948 6914 15976 17156
rect 16856 17196 16908 17202
rect 16856 17138 16908 17144
rect 17328 16998 17356 17206
rect 17868 17196 17920 17202
rect 17972 17184 18000 17478
rect 17920 17156 18000 17184
rect 17868 17138 17920 17144
rect 17132 16992 17184 16998
rect 17132 16934 17184 16940
rect 17316 16992 17368 16998
rect 17316 16934 17368 16940
rect 17868 16992 17920 16998
rect 17868 16934 17920 16940
rect 17144 16590 17172 16934
rect 17132 16584 17184 16590
rect 17132 16526 17184 16532
rect 16028 16516 16080 16522
rect 16028 16458 16080 16464
rect 16040 16182 16068 16458
rect 16028 16176 16080 16182
rect 16028 16118 16080 16124
rect 16040 14890 16068 16118
rect 16304 15904 16356 15910
rect 16304 15846 16356 15852
rect 16120 15360 16172 15366
rect 16120 15302 16172 15308
rect 16132 14958 16160 15302
rect 16316 15162 16344 15846
rect 16304 15156 16356 15162
rect 16304 15098 16356 15104
rect 16120 14952 16172 14958
rect 16120 14894 16172 14900
rect 16028 14884 16080 14890
rect 16028 14826 16080 14832
rect 16040 14550 16068 14826
rect 16028 14544 16080 14550
rect 16028 14486 16080 14492
rect 16040 14006 16068 14486
rect 16132 14074 16160 14894
rect 16304 14340 16356 14346
rect 16304 14282 16356 14288
rect 16316 14074 16344 14282
rect 16120 14068 16172 14074
rect 16120 14010 16172 14016
rect 16304 14068 16356 14074
rect 16304 14010 16356 14016
rect 16028 14000 16080 14006
rect 16028 13942 16080 13948
rect 16580 13932 16632 13938
rect 16580 13874 16632 13880
rect 16592 13530 16620 13874
rect 17328 13802 17356 16934
rect 17880 16726 17908 16934
rect 17868 16720 17920 16726
rect 17868 16662 17920 16668
rect 17972 16454 18000 17156
rect 17960 16448 18012 16454
rect 17960 16390 18012 16396
rect 18064 14550 18092 18702
rect 18052 14544 18104 14550
rect 18052 14486 18104 14492
rect 18064 14074 18092 14486
rect 18156 14482 18184 19110
rect 18248 18222 18276 20470
rect 18315 20156 18623 20165
rect 18315 20154 18321 20156
rect 18377 20154 18401 20156
rect 18457 20154 18481 20156
rect 18537 20154 18561 20156
rect 18617 20154 18623 20156
rect 18377 20102 18379 20154
rect 18559 20102 18561 20154
rect 18315 20100 18321 20102
rect 18377 20100 18401 20102
rect 18457 20100 18481 20102
rect 18537 20100 18561 20102
rect 18617 20100 18623 20102
rect 18315 20091 18623 20100
rect 18880 19440 18932 19446
rect 18880 19382 18932 19388
rect 18696 19236 18748 19242
rect 18696 19178 18748 19184
rect 18788 19236 18840 19242
rect 18788 19178 18840 19184
rect 18708 19145 18736 19178
rect 18694 19136 18750 19145
rect 18315 19068 18623 19077
rect 18694 19071 18750 19080
rect 18315 19066 18321 19068
rect 18377 19066 18401 19068
rect 18457 19066 18481 19068
rect 18537 19066 18561 19068
rect 18617 19066 18623 19068
rect 18377 19014 18379 19066
rect 18559 19014 18561 19066
rect 18315 19012 18321 19014
rect 18377 19012 18401 19014
rect 18457 19012 18481 19014
rect 18537 19012 18561 19014
rect 18617 19012 18623 19014
rect 18315 19003 18623 19012
rect 18800 18970 18828 19178
rect 18788 18964 18840 18970
rect 18788 18906 18840 18912
rect 18512 18624 18564 18630
rect 18512 18566 18564 18572
rect 18524 18358 18552 18566
rect 18512 18352 18564 18358
rect 18512 18294 18564 18300
rect 18236 18216 18288 18222
rect 18236 18158 18288 18164
rect 18248 16794 18276 18158
rect 18315 17980 18623 17989
rect 18315 17978 18321 17980
rect 18377 17978 18401 17980
rect 18457 17978 18481 17980
rect 18537 17978 18561 17980
rect 18617 17978 18623 17980
rect 18377 17926 18379 17978
rect 18559 17926 18561 17978
rect 18315 17924 18321 17926
rect 18377 17924 18401 17926
rect 18457 17924 18481 17926
rect 18537 17924 18561 17926
rect 18617 17924 18623 17926
rect 18315 17915 18623 17924
rect 18696 17672 18748 17678
rect 18696 17614 18748 17620
rect 18420 17536 18472 17542
rect 18420 17478 18472 17484
rect 18432 17338 18460 17478
rect 18420 17332 18472 17338
rect 18420 17274 18472 17280
rect 18708 17066 18736 17614
rect 18788 17196 18840 17202
rect 18788 17138 18840 17144
rect 18696 17060 18748 17066
rect 18696 17002 18748 17008
rect 18315 16892 18623 16901
rect 18315 16890 18321 16892
rect 18377 16890 18401 16892
rect 18457 16890 18481 16892
rect 18537 16890 18561 16892
rect 18617 16890 18623 16892
rect 18377 16838 18379 16890
rect 18559 16838 18561 16890
rect 18315 16836 18321 16838
rect 18377 16836 18401 16838
rect 18457 16836 18481 16838
rect 18537 16836 18561 16838
rect 18617 16836 18623 16838
rect 18315 16827 18623 16836
rect 18800 16794 18828 17138
rect 18236 16788 18288 16794
rect 18236 16730 18288 16736
rect 18788 16788 18840 16794
rect 18788 16730 18840 16736
rect 18144 14476 18196 14482
rect 18144 14418 18196 14424
rect 18248 14414 18276 16730
rect 18892 16572 18920 19382
rect 18972 19372 19024 19378
rect 18972 19314 19024 19320
rect 18984 18766 19012 19314
rect 18972 18760 19024 18766
rect 18972 18702 19024 18708
rect 19076 17270 19104 22374
rect 19444 22030 19472 24142
rect 19708 24132 19760 24138
rect 19708 24074 19760 24080
rect 19720 23866 19748 24074
rect 19708 23860 19760 23866
rect 19708 23802 19760 23808
rect 19800 23792 19852 23798
rect 19800 23734 19852 23740
rect 19812 23186 19840 23734
rect 19904 23730 19932 24550
rect 19892 23724 19944 23730
rect 19892 23666 19944 23672
rect 19800 23180 19852 23186
rect 19800 23122 19852 23128
rect 19812 22642 19840 23122
rect 19984 22976 20036 22982
rect 19984 22918 20036 22924
rect 19800 22636 19852 22642
rect 19800 22578 19852 22584
rect 19996 22506 20024 22918
rect 19984 22500 20036 22506
rect 19984 22442 20036 22448
rect 19432 22024 19484 22030
rect 19432 21966 19484 21972
rect 19708 21956 19760 21962
rect 19708 21898 19760 21904
rect 19720 21554 19748 21898
rect 19708 21548 19760 21554
rect 19708 21490 19760 21496
rect 19340 20868 19392 20874
rect 19340 20810 19392 20816
rect 19352 19360 19380 20810
rect 19524 20800 19576 20806
rect 19524 20742 19576 20748
rect 19536 20534 19564 20742
rect 19524 20528 19576 20534
rect 19524 20470 19576 20476
rect 19720 19378 19748 21490
rect 19708 19372 19760 19378
rect 19352 19332 19472 19360
rect 19156 19304 19208 19310
rect 19208 19264 19288 19292
rect 19156 19246 19208 19252
rect 19260 19258 19288 19264
rect 19260 19230 19380 19258
rect 19156 19168 19208 19174
rect 19154 19136 19156 19145
rect 19248 19168 19300 19174
rect 19208 19136 19210 19145
rect 19248 19110 19300 19116
rect 19154 19071 19210 19080
rect 19260 18970 19288 19110
rect 19248 18964 19300 18970
rect 19248 18906 19300 18912
rect 19352 18834 19380 19230
rect 19340 18828 19392 18834
rect 19340 18770 19392 18776
rect 19064 17264 19116 17270
rect 19064 17206 19116 17212
rect 19352 17134 19380 18770
rect 19340 17128 19392 17134
rect 19340 17070 19392 17076
rect 18972 16584 19024 16590
rect 18892 16544 18972 16572
rect 18972 16526 19024 16532
rect 19444 16454 19472 19332
rect 19708 19314 19760 19320
rect 19616 19304 19668 19310
rect 19616 19246 19668 19252
rect 19628 18766 19656 19246
rect 19720 18970 19748 19314
rect 19800 19304 19852 19310
rect 19800 19246 19852 19252
rect 19708 18964 19760 18970
rect 19708 18906 19760 18912
rect 19812 18834 19840 19246
rect 19996 19174 20024 22442
rect 20088 19310 20116 29106
rect 20180 25906 20208 32422
rect 20272 29832 20300 32778
rect 20364 31958 20392 32846
rect 20732 32298 20760 33934
rect 20824 32978 20852 36110
rect 20916 35290 20944 38898
rect 21652 38350 21680 45222
rect 23216 44878 23244 45902
rect 23204 44872 23256 44878
rect 23204 44814 23256 44820
rect 21788 44636 22096 44645
rect 21788 44634 21794 44636
rect 21850 44634 21874 44636
rect 21930 44634 21954 44636
rect 22010 44634 22034 44636
rect 22090 44634 22096 44636
rect 21850 44582 21852 44634
rect 22032 44582 22034 44634
rect 21788 44580 21794 44582
rect 21850 44580 21874 44582
rect 21930 44580 21954 44582
rect 22010 44580 22034 44582
rect 22090 44580 22096 44582
rect 21788 44571 22096 44580
rect 21788 43548 22096 43557
rect 21788 43546 21794 43548
rect 21850 43546 21874 43548
rect 21930 43546 21954 43548
rect 22010 43546 22034 43548
rect 22090 43546 22096 43548
rect 21850 43494 21852 43546
rect 22032 43494 22034 43546
rect 21788 43492 21794 43494
rect 21850 43492 21874 43494
rect 21930 43492 21954 43494
rect 22010 43492 22034 43494
rect 22090 43492 22096 43494
rect 21788 43483 22096 43492
rect 21788 42460 22096 42469
rect 21788 42458 21794 42460
rect 21850 42458 21874 42460
rect 21930 42458 21954 42460
rect 22010 42458 22034 42460
rect 22090 42458 22096 42460
rect 21850 42406 21852 42458
rect 22032 42406 22034 42458
rect 21788 42404 21794 42406
rect 21850 42404 21874 42406
rect 21930 42404 21954 42406
rect 22010 42404 22034 42406
rect 22090 42404 22096 42406
rect 21788 42395 22096 42404
rect 21788 41372 22096 41381
rect 21788 41370 21794 41372
rect 21850 41370 21874 41372
rect 21930 41370 21954 41372
rect 22010 41370 22034 41372
rect 22090 41370 22096 41372
rect 21850 41318 21852 41370
rect 22032 41318 22034 41370
rect 21788 41316 21794 41318
rect 21850 41316 21874 41318
rect 21930 41316 21954 41318
rect 22010 41316 22034 41318
rect 22090 41316 22096 41318
rect 21788 41307 22096 41316
rect 21788 40284 22096 40293
rect 21788 40282 21794 40284
rect 21850 40282 21874 40284
rect 21930 40282 21954 40284
rect 22010 40282 22034 40284
rect 22090 40282 22096 40284
rect 21850 40230 21852 40282
rect 22032 40230 22034 40282
rect 21788 40228 21794 40230
rect 21850 40228 21874 40230
rect 21930 40228 21954 40230
rect 22010 40228 22034 40230
rect 22090 40228 22096 40230
rect 21788 40219 22096 40228
rect 21788 39196 22096 39205
rect 21788 39194 21794 39196
rect 21850 39194 21874 39196
rect 21930 39194 21954 39196
rect 22010 39194 22034 39196
rect 22090 39194 22096 39196
rect 21850 39142 21852 39194
rect 22032 39142 22034 39194
rect 21788 39140 21794 39142
rect 21850 39140 21874 39142
rect 21930 39140 21954 39142
rect 22010 39140 22034 39142
rect 22090 39140 22096 39142
rect 21788 39131 22096 39140
rect 23492 38894 23520 46854
rect 22192 38888 22244 38894
rect 22192 38830 22244 38836
rect 23480 38888 23532 38894
rect 23480 38830 23532 38836
rect 22204 38554 22232 38830
rect 23112 38820 23164 38826
rect 23112 38762 23164 38768
rect 22192 38548 22244 38554
rect 22192 38490 22244 38496
rect 21640 38344 21692 38350
rect 21640 38286 21692 38292
rect 21788 38108 22096 38117
rect 21788 38106 21794 38108
rect 21850 38106 21874 38108
rect 21930 38106 21954 38108
rect 22010 38106 22034 38108
rect 22090 38106 22096 38108
rect 21850 38054 21852 38106
rect 22032 38054 22034 38106
rect 21788 38052 21794 38054
rect 21850 38052 21874 38054
rect 21930 38052 21954 38054
rect 22010 38052 22034 38054
rect 22090 38052 22096 38054
rect 21788 38043 22096 38052
rect 22376 37324 22428 37330
rect 22376 37266 22428 37272
rect 21456 37256 21508 37262
rect 21456 37198 21508 37204
rect 21468 37126 21496 37198
rect 21456 37120 21508 37126
rect 21456 37062 21508 37068
rect 21468 36854 21496 37062
rect 21788 37020 22096 37029
rect 21788 37018 21794 37020
rect 21850 37018 21874 37020
rect 21930 37018 21954 37020
rect 22010 37018 22034 37020
rect 22090 37018 22096 37020
rect 21850 36966 21852 37018
rect 22032 36966 22034 37018
rect 21788 36964 21794 36966
rect 21850 36964 21874 36966
rect 21930 36964 21954 36966
rect 22010 36964 22034 36966
rect 22090 36964 22096 36966
rect 21788 36955 22096 36964
rect 21456 36848 21508 36854
rect 21456 36790 21508 36796
rect 21272 36780 21324 36786
rect 21272 36722 21324 36728
rect 21284 36174 21312 36722
rect 21272 36168 21324 36174
rect 21272 36110 21324 36116
rect 21284 35290 21312 36110
rect 20904 35284 20956 35290
rect 20904 35226 20956 35232
rect 21272 35284 21324 35290
rect 21272 35226 21324 35232
rect 21180 34740 21232 34746
rect 21180 34682 21232 34688
rect 20904 33856 20956 33862
rect 20904 33798 20956 33804
rect 20916 33522 20944 33798
rect 20904 33516 20956 33522
rect 20904 33458 20956 33464
rect 20812 32972 20864 32978
rect 20812 32914 20864 32920
rect 20720 32292 20772 32298
rect 20720 32234 20772 32240
rect 20824 32026 20852 32914
rect 20812 32020 20864 32026
rect 20812 31962 20864 31968
rect 20352 31952 20404 31958
rect 20352 31894 20404 31900
rect 20364 31822 20392 31894
rect 20352 31816 20404 31822
rect 20352 31758 20404 31764
rect 20352 29844 20404 29850
rect 20272 29804 20352 29832
rect 20272 29306 20300 29804
rect 20352 29786 20404 29792
rect 20260 29300 20312 29306
rect 20260 29242 20312 29248
rect 20812 29232 20864 29238
rect 20812 29174 20864 29180
rect 20824 28558 20852 29174
rect 20812 28552 20864 28558
rect 20812 28494 20864 28500
rect 20260 28008 20312 28014
rect 20260 27950 20312 27956
rect 20272 27130 20300 27950
rect 20260 27124 20312 27130
rect 20260 27066 20312 27072
rect 20168 25900 20220 25906
rect 20168 25842 20220 25848
rect 20180 24750 20208 25842
rect 20168 24744 20220 24750
rect 20168 24686 20220 24692
rect 20180 23186 20208 24686
rect 20272 23798 20300 27066
rect 20720 27056 20772 27062
rect 20720 26998 20772 27004
rect 20732 25294 20760 26998
rect 20916 26908 20944 33458
rect 21192 32434 21220 34682
rect 21284 34678 21312 35226
rect 21272 34672 21324 34678
rect 21272 34614 21324 34620
rect 21272 33992 21324 33998
rect 21272 33934 21324 33940
rect 21284 33454 21312 33934
rect 21364 33924 21416 33930
rect 21364 33866 21416 33872
rect 21376 33658 21404 33866
rect 21364 33652 21416 33658
rect 21364 33594 21416 33600
rect 21468 33522 21496 36790
rect 21788 35932 22096 35941
rect 21788 35930 21794 35932
rect 21850 35930 21874 35932
rect 21930 35930 21954 35932
rect 22010 35930 22034 35932
rect 22090 35930 22096 35932
rect 21850 35878 21852 35930
rect 22032 35878 22034 35930
rect 21788 35876 21794 35878
rect 21850 35876 21874 35878
rect 21930 35876 21954 35878
rect 22010 35876 22034 35878
rect 22090 35876 22096 35878
rect 21788 35867 22096 35876
rect 22388 35086 22416 37266
rect 22744 37120 22796 37126
rect 22744 37062 22796 37068
rect 22756 36174 22784 37062
rect 22744 36168 22796 36174
rect 22744 36110 22796 36116
rect 23020 36032 23072 36038
rect 23020 35974 23072 35980
rect 23032 35698 23060 35974
rect 23020 35692 23072 35698
rect 23020 35634 23072 35640
rect 22836 35488 22888 35494
rect 22836 35430 22888 35436
rect 22376 35080 22428 35086
rect 22376 35022 22428 35028
rect 21788 34844 22096 34853
rect 21788 34842 21794 34844
rect 21850 34842 21874 34844
rect 21930 34842 21954 34844
rect 22010 34842 22034 34844
rect 22090 34842 22096 34844
rect 21850 34790 21852 34842
rect 22032 34790 22034 34842
rect 21788 34788 21794 34790
rect 21850 34788 21874 34790
rect 21930 34788 21954 34790
rect 22010 34788 22034 34790
rect 22090 34788 22096 34790
rect 21788 34779 22096 34788
rect 22848 34678 22876 35430
rect 22836 34672 22888 34678
rect 22836 34614 22888 34620
rect 22560 34536 22612 34542
rect 22560 34478 22612 34484
rect 21788 33756 22096 33765
rect 21788 33754 21794 33756
rect 21850 33754 21874 33756
rect 21930 33754 21954 33756
rect 22010 33754 22034 33756
rect 22090 33754 22096 33756
rect 21850 33702 21852 33754
rect 22032 33702 22034 33754
rect 21788 33700 21794 33702
rect 21850 33700 21874 33702
rect 21930 33700 21954 33702
rect 22010 33700 22034 33702
rect 22090 33700 22096 33702
rect 21788 33691 22096 33700
rect 21456 33516 21508 33522
rect 21456 33458 21508 33464
rect 21272 33448 21324 33454
rect 21272 33390 21324 33396
rect 21180 32428 21232 32434
rect 21180 32370 21232 32376
rect 21192 32314 21220 32370
rect 21100 32286 21220 32314
rect 21100 31346 21128 32286
rect 21284 31822 21312 33390
rect 21468 32502 21496 33458
rect 22572 33454 22600 34478
rect 22560 33448 22612 33454
rect 22560 33390 22612 33396
rect 21788 32668 22096 32677
rect 21788 32666 21794 32668
rect 21850 32666 21874 32668
rect 21930 32666 21954 32668
rect 22010 32666 22034 32668
rect 22090 32666 22096 32668
rect 21850 32614 21852 32666
rect 22032 32614 22034 32666
rect 21788 32612 21794 32614
rect 21850 32612 21874 32614
rect 21930 32612 21954 32614
rect 22010 32612 22034 32614
rect 22090 32612 22096 32614
rect 21788 32603 22096 32612
rect 21456 32496 21508 32502
rect 21456 32438 21508 32444
rect 21272 31816 21324 31822
rect 21192 31776 21272 31804
rect 21088 31340 21140 31346
rect 21088 31282 21140 31288
rect 21100 30394 21128 31282
rect 21088 30388 21140 30394
rect 21088 30330 21140 30336
rect 21100 29850 21128 30330
rect 21088 29844 21140 29850
rect 21088 29786 21140 29792
rect 21192 29646 21220 31776
rect 21272 31758 21324 31764
rect 21180 29640 21232 29646
rect 21180 29582 21232 29588
rect 21272 29504 21324 29510
rect 21272 29446 21324 29452
rect 21284 29102 21312 29446
rect 21272 29096 21324 29102
rect 21272 29038 21324 29044
rect 21088 27328 21140 27334
rect 21088 27270 21140 27276
rect 20824 26880 20944 26908
rect 20720 25288 20772 25294
rect 20720 25230 20772 25236
rect 20444 24812 20496 24818
rect 20444 24754 20496 24760
rect 20456 23866 20484 24754
rect 20444 23860 20496 23866
rect 20444 23802 20496 23808
rect 20260 23792 20312 23798
rect 20260 23734 20312 23740
rect 20168 23180 20220 23186
rect 20168 23122 20220 23128
rect 20536 23180 20588 23186
rect 20536 23122 20588 23128
rect 20548 20942 20576 23122
rect 20720 23112 20772 23118
rect 20720 23054 20772 23060
rect 20732 22778 20760 23054
rect 20720 22772 20772 22778
rect 20720 22714 20772 22720
rect 20720 21956 20772 21962
rect 20720 21898 20772 21904
rect 20732 21690 20760 21898
rect 20720 21684 20772 21690
rect 20720 21626 20772 21632
rect 20536 20936 20588 20942
rect 20536 20878 20588 20884
rect 20352 20800 20404 20806
rect 20352 20742 20404 20748
rect 20364 20262 20392 20742
rect 20352 20256 20404 20262
rect 20352 20198 20404 20204
rect 20076 19304 20128 19310
rect 20076 19246 20128 19252
rect 19984 19168 20036 19174
rect 19984 19110 20036 19116
rect 19800 18828 19852 18834
rect 19800 18770 19852 18776
rect 19616 18760 19668 18766
rect 19616 18702 19668 18708
rect 19628 17882 19656 18702
rect 19616 17876 19668 17882
rect 19616 17818 19668 17824
rect 19892 17672 19944 17678
rect 19892 17614 19944 17620
rect 19904 17338 19932 17614
rect 19892 17332 19944 17338
rect 19892 17274 19944 17280
rect 19616 17196 19668 17202
rect 19536 17156 19616 17184
rect 19432 16448 19484 16454
rect 19432 16390 19484 16396
rect 18315 15804 18623 15813
rect 18315 15802 18321 15804
rect 18377 15802 18401 15804
rect 18457 15802 18481 15804
rect 18537 15802 18561 15804
rect 18617 15802 18623 15804
rect 18377 15750 18379 15802
rect 18559 15750 18561 15802
rect 18315 15748 18321 15750
rect 18377 15748 18401 15750
rect 18457 15748 18481 15750
rect 18537 15748 18561 15750
rect 18617 15748 18623 15750
rect 18315 15739 18623 15748
rect 19340 15020 19392 15026
rect 19340 14962 19392 14968
rect 19064 14952 19116 14958
rect 19064 14894 19116 14900
rect 18315 14716 18623 14725
rect 18315 14714 18321 14716
rect 18377 14714 18401 14716
rect 18457 14714 18481 14716
rect 18537 14714 18561 14716
rect 18617 14714 18623 14716
rect 18377 14662 18379 14714
rect 18559 14662 18561 14714
rect 18315 14660 18321 14662
rect 18377 14660 18401 14662
rect 18457 14660 18481 14662
rect 18537 14660 18561 14662
rect 18617 14660 18623 14662
rect 18315 14651 18623 14660
rect 19076 14414 19104 14894
rect 18236 14408 18288 14414
rect 18236 14350 18288 14356
rect 19064 14408 19116 14414
rect 19064 14350 19116 14356
rect 18052 14068 18104 14074
rect 18052 14010 18104 14016
rect 18248 13938 18276 14350
rect 18512 14272 18564 14278
rect 18512 14214 18564 14220
rect 18524 13938 18552 14214
rect 19076 14006 19104 14350
rect 19064 14000 19116 14006
rect 19064 13942 19116 13948
rect 17592 13932 17644 13938
rect 17592 13874 17644 13880
rect 18236 13932 18288 13938
rect 18236 13874 18288 13880
rect 18512 13932 18564 13938
rect 18512 13874 18564 13880
rect 17316 13796 17368 13802
rect 17316 13738 17368 13744
rect 16764 13728 16816 13734
rect 16764 13670 16816 13676
rect 16580 13524 16632 13530
rect 16580 13466 16632 13472
rect 16776 13326 16804 13670
rect 16764 13320 16816 13326
rect 16764 13262 16816 13268
rect 15856 6886 15976 6914
rect 14842 6556 15150 6565
rect 14842 6554 14848 6556
rect 14904 6554 14928 6556
rect 14984 6554 15008 6556
rect 15064 6554 15088 6556
rect 15144 6554 15150 6556
rect 14904 6502 14906 6554
rect 15086 6502 15088 6554
rect 14842 6500 14848 6502
rect 14904 6500 14928 6502
rect 14984 6500 15008 6502
rect 15064 6500 15088 6502
rect 15144 6500 15150 6502
rect 14842 6491 15150 6500
rect 14842 5468 15150 5477
rect 14842 5466 14848 5468
rect 14904 5466 14928 5468
rect 14984 5466 15008 5468
rect 15064 5466 15088 5468
rect 15144 5466 15150 5468
rect 14904 5414 14906 5466
rect 15086 5414 15088 5466
rect 14842 5412 14848 5414
rect 14904 5412 14928 5414
rect 14984 5412 15008 5414
rect 15064 5412 15088 5414
rect 15144 5412 15150 5414
rect 14842 5403 15150 5412
rect 14842 4380 15150 4389
rect 14842 4378 14848 4380
rect 14904 4378 14928 4380
rect 14984 4378 15008 4380
rect 15064 4378 15088 4380
rect 15144 4378 15150 4380
rect 14904 4326 14906 4378
rect 15086 4326 15088 4378
rect 14842 4324 14848 4326
rect 14904 4324 14928 4326
rect 14984 4324 15008 4326
rect 15064 4324 15088 4326
rect 15144 4324 15150 4326
rect 14842 4315 15150 4324
rect 13636 4072 13688 4078
rect 13636 4014 13688 4020
rect 13544 3528 13596 3534
rect 13544 3470 13596 3476
rect 12992 3188 13044 3194
rect 12992 3130 13044 3136
rect 13556 3058 13584 3470
rect 13544 3052 13596 3058
rect 13544 2994 13596 3000
rect 11369 2748 11677 2757
rect 11369 2746 11375 2748
rect 11431 2746 11455 2748
rect 11511 2746 11535 2748
rect 11591 2746 11615 2748
rect 11671 2746 11677 2748
rect 11431 2694 11433 2746
rect 11613 2694 11615 2746
rect 11369 2692 11375 2694
rect 11431 2692 11455 2694
rect 11511 2692 11535 2694
rect 11591 2692 11615 2694
rect 11671 2692 11677 2694
rect 11369 2683 11677 2692
rect 13648 1986 13676 4014
rect 14004 3528 14056 3534
rect 14004 3470 14056 3476
rect 14016 3058 14044 3470
rect 14188 3392 14240 3398
rect 14188 3334 14240 3340
rect 14200 3126 14228 3334
rect 14842 3292 15150 3301
rect 14842 3290 14848 3292
rect 14904 3290 14928 3292
rect 14984 3290 15008 3292
rect 15064 3290 15088 3292
rect 15144 3290 15150 3292
rect 14904 3238 14906 3290
rect 15086 3238 15088 3290
rect 14842 3236 14848 3238
rect 14904 3236 14928 3238
rect 14984 3236 15008 3238
rect 15064 3236 15088 3238
rect 15144 3236 15150 3238
rect 14842 3227 15150 3236
rect 14188 3120 14240 3126
rect 14188 3062 14240 3068
rect 14004 3052 14056 3058
rect 14004 2994 14056 3000
rect 14740 2984 14792 2990
rect 14740 2926 14792 2932
rect 13556 1958 13676 1986
rect 13556 800 13584 1958
rect 14752 1714 14780 2926
rect 15856 2582 15884 6886
rect 16212 3528 16264 3534
rect 16212 3470 16264 3476
rect 16224 3058 16252 3470
rect 17040 3392 17092 3398
rect 17040 3334 17092 3340
rect 17052 3126 17080 3334
rect 17040 3120 17092 3126
rect 17040 3062 17092 3068
rect 16212 3052 16264 3058
rect 16212 2994 16264 3000
rect 16764 2984 16816 2990
rect 16764 2926 16816 2932
rect 15844 2576 15896 2582
rect 15844 2518 15896 2524
rect 16120 2372 16172 2378
rect 16120 2314 16172 2320
rect 14842 2204 15150 2213
rect 14842 2202 14848 2204
rect 14904 2202 14928 2204
rect 14984 2202 15008 2204
rect 15064 2202 15088 2204
rect 15144 2202 15150 2204
rect 14904 2150 14906 2202
rect 15086 2150 15088 2202
rect 14842 2148 14848 2150
rect 14904 2148 14928 2150
rect 14984 2148 15008 2150
rect 15064 2148 15088 2150
rect 15144 2148 15150 2150
rect 14842 2139 15150 2148
rect 14752 1686 14872 1714
rect 14844 800 14872 1686
rect 16132 800 16160 2314
rect 16776 800 16804 2926
rect 17604 2650 17632 13874
rect 18315 13628 18623 13637
rect 18315 13626 18321 13628
rect 18377 13626 18401 13628
rect 18457 13626 18481 13628
rect 18537 13626 18561 13628
rect 18617 13626 18623 13628
rect 18377 13574 18379 13626
rect 18559 13574 18561 13626
rect 18315 13572 18321 13574
rect 18377 13572 18401 13574
rect 18457 13572 18481 13574
rect 18537 13572 18561 13574
rect 18617 13572 18623 13574
rect 18315 13563 18623 13572
rect 19352 12986 19380 14962
rect 19444 13530 19472 16390
rect 19536 14074 19564 17156
rect 19616 17138 19668 17144
rect 20364 16250 20392 20198
rect 20720 19372 20772 19378
rect 20720 19314 20772 19320
rect 20732 18698 20760 19314
rect 20720 18692 20772 18698
rect 20720 18634 20772 18640
rect 20732 18290 20760 18634
rect 20720 18284 20772 18290
rect 20720 18226 20772 18232
rect 20444 16652 20496 16658
rect 20444 16594 20496 16600
rect 20352 16244 20404 16250
rect 20352 16186 20404 16192
rect 20456 15706 20484 16594
rect 20824 16590 20852 26880
rect 20904 26580 20956 26586
rect 20904 26522 20956 26528
rect 20916 23866 20944 26522
rect 21100 24886 21128 27270
rect 21180 26784 21232 26790
rect 21180 26726 21232 26732
rect 21192 26382 21220 26726
rect 21180 26376 21232 26382
rect 21180 26318 21232 26324
rect 21088 24880 21140 24886
rect 21088 24822 21140 24828
rect 21180 24744 21232 24750
rect 21180 24686 21232 24692
rect 20996 24064 21048 24070
rect 20996 24006 21048 24012
rect 20904 23860 20956 23866
rect 20904 23802 20956 23808
rect 21008 23798 21036 24006
rect 20996 23792 21048 23798
rect 20996 23734 21048 23740
rect 20904 22976 20956 22982
rect 20904 22918 20956 22924
rect 20916 21554 20944 22918
rect 20904 21548 20956 21554
rect 20904 21490 20956 21496
rect 20812 16584 20864 16590
rect 20812 16526 20864 16532
rect 20824 16232 20852 16526
rect 20732 16204 20852 16232
rect 20732 16046 20760 16204
rect 20812 16108 20864 16114
rect 20812 16050 20864 16056
rect 20720 16040 20772 16046
rect 20720 15982 20772 15988
rect 20444 15700 20496 15706
rect 20444 15642 20496 15648
rect 19616 15632 19668 15638
rect 19616 15574 19668 15580
rect 19628 15094 19656 15574
rect 20732 15502 20760 15982
rect 20720 15496 20772 15502
rect 20720 15438 20772 15444
rect 20536 15360 20588 15366
rect 20536 15302 20588 15308
rect 19616 15088 19668 15094
rect 19616 15030 19668 15036
rect 20444 14816 20496 14822
rect 20548 14804 20576 15302
rect 20496 14776 20576 14804
rect 20444 14758 20496 14764
rect 19708 14340 19760 14346
rect 19708 14282 19760 14288
rect 19524 14068 19576 14074
rect 19524 14010 19576 14016
rect 19432 13524 19484 13530
rect 19432 13466 19484 13472
rect 19340 12980 19392 12986
rect 19340 12922 19392 12928
rect 18315 12540 18623 12549
rect 18315 12538 18321 12540
rect 18377 12538 18401 12540
rect 18457 12538 18481 12540
rect 18537 12538 18561 12540
rect 18617 12538 18623 12540
rect 18377 12486 18379 12538
rect 18559 12486 18561 12538
rect 18315 12484 18321 12486
rect 18377 12484 18401 12486
rect 18457 12484 18481 12486
rect 18537 12484 18561 12486
rect 18617 12484 18623 12486
rect 18315 12475 18623 12484
rect 19432 12232 19484 12238
rect 19432 12174 19484 12180
rect 19444 11898 19472 12174
rect 19432 11892 19484 11898
rect 19432 11834 19484 11840
rect 18315 11452 18623 11461
rect 18315 11450 18321 11452
rect 18377 11450 18401 11452
rect 18457 11450 18481 11452
rect 18537 11450 18561 11452
rect 18617 11450 18623 11452
rect 18377 11398 18379 11450
rect 18559 11398 18561 11450
rect 18315 11396 18321 11398
rect 18377 11396 18401 11398
rect 18457 11396 18481 11398
rect 18537 11396 18561 11398
rect 18617 11396 18623 11398
rect 18315 11387 18623 11396
rect 19536 11234 19564 14010
rect 19616 12844 19668 12850
rect 19616 12786 19668 12792
rect 19628 11354 19656 12786
rect 19720 12442 19748 14282
rect 19800 13524 19852 13530
rect 19800 13466 19852 13472
rect 19708 12436 19760 12442
rect 19708 12378 19760 12384
rect 19812 11694 19840 13466
rect 20352 12096 20404 12102
rect 20352 12038 20404 12044
rect 20364 11762 20392 12038
rect 20456 11898 20484 14758
rect 20824 14618 20852 16050
rect 21008 15570 21036 23734
rect 21192 23662 21220 24686
rect 21180 23656 21232 23662
rect 21180 23598 21232 23604
rect 21284 23474 21312 29038
rect 21468 27606 21496 32438
rect 23124 32434 23152 38762
rect 23768 37262 23796 47126
rect 24044 47054 24072 49286
rect 25106 49200 25218 49800
rect 25750 49200 25862 49800
rect 26394 49200 26506 49800
rect 27038 49314 27150 49800
rect 26620 49286 27150 49314
rect 26146 49056 26202 49065
rect 26146 48991 26202 49000
rect 25261 47356 25569 47365
rect 25261 47354 25267 47356
rect 25323 47354 25347 47356
rect 25403 47354 25427 47356
rect 25483 47354 25507 47356
rect 25563 47354 25569 47356
rect 25323 47302 25325 47354
rect 25505 47302 25507 47354
rect 25261 47300 25267 47302
rect 25323 47300 25347 47302
rect 25403 47300 25427 47302
rect 25483 47300 25507 47302
rect 25563 47300 25569 47302
rect 25261 47291 25569 47300
rect 25044 47184 25096 47190
rect 25044 47126 25096 47132
rect 24032 47048 24084 47054
rect 24032 46990 24084 46996
rect 24952 45960 25004 45966
rect 24952 45902 25004 45908
rect 24964 44334 24992 45902
rect 25056 44470 25084 47126
rect 26054 47016 26110 47025
rect 26054 46951 26110 46960
rect 25261 46268 25569 46277
rect 25261 46266 25267 46268
rect 25323 46266 25347 46268
rect 25403 46266 25427 46268
rect 25483 46266 25507 46268
rect 25563 46266 25569 46268
rect 25323 46214 25325 46266
rect 25505 46214 25507 46266
rect 25261 46212 25267 46214
rect 25323 46212 25347 46214
rect 25403 46212 25427 46214
rect 25483 46212 25507 46214
rect 25563 46212 25569 46214
rect 25261 46203 25569 46212
rect 26068 45422 26096 46951
rect 26056 45416 26108 45422
rect 26056 45358 26108 45364
rect 25261 45180 25569 45189
rect 25261 45178 25267 45180
rect 25323 45178 25347 45180
rect 25403 45178 25427 45180
rect 25483 45178 25507 45180
rect 25563 45178 25569 45180
rect 25323 45126 25325 45178
rect 25505 45126 25507 45178
rect 25261 45124 25267 45126
rect 25323 45124 25347 45126
rect 25403 45124 25427 45126
rect 25483 45124 25507 45126
rect 25563 45124 25569 45126
rect 25261 45115 25569 45124
rect 25044 44464 25096 44470
rect 25044 44406 25096 44412
rect 26160 44334 26188 48991
rect 26620 47410 26648 49286
rect 27038 49200 27150 49286
rect 27682 49200 27794 49800
rect 28326 49200 28438 49800
rect 28970 49200 29082 49800
rect 29614 49200 29726 49800
rect 26344 47382 26648 47410
rect 26240 44872 26292 44878
rect 26240 44814 26292 44820
rect 24952 44328 25004 44334
rect 24952 44270 25004 44276
rect 26148 44328 26200 44334
rect 26148 44270 26200 44276
rect 25261 44092 25569 44101
rect 25261 44090 25267 44092
rect 25323 44090 25347 44092
rect 25403 44090 25427 44092
rect 25483 44090 25507 44092
rect 25563 44090 25569 44092
rect 25323 44038 25325 44090
rect 25505 44038 25507 44090
rect 25261 44036 25267 44038
rect 25323 44036 25347 44038
rect 25403 44036 25427 44038
rect 25483 44036 25507 44038
rect 25563 44036 25569 44038
rect 25261 44027 25569 44036
rect 26252 43858 26280 44814
rect 26240 43852 26292 43858
rect 26240 43794 26292 43800
rect 25261 43004 25569 43013
rect 25261 43002 25267 43004
rect 25323 43002 25347 43004
rect 25403 43002 25427 43004
rect 25483 43002 25507 43004
rect 25563 43002 25569 43004
rect 25323 42950 25325 43002
rect 25505 42950 25507 43002
rect 25261 42948 25267 42950
rect 25323 42948 25347 42950
rect 25403 42948 25427 42950
rect 25483 42948 25507 42950
rect 25563 42948 25569 42950
rect 25261 42939 25569 42948
rect 26054 42256 26110 42265
rect 26054 42191 26110 42200
rect 25261 41916 25569 41925
rect 25261 41914 25267 41916
rect 25323 41914 25347 41916
rect 25403 41914 25427 41916
rect 25483 41914 25507 41916
rect 25563 41914 25569 41916
rect 25323 41862 25325 41914
rect 25505 41862 25507 41914
rect 25261 41860 25267 41862
rect 25323 41860 25347 41862
rect 25403 41860 25427 41862
rect 25483 41860 25507 41862
rect 25563 41860 25569 41862
rect 25261 41851 25569 41860
rect 25261 40828 25569 40837
rect 25261 40826 25267 40828
rect 25323 40826 25347 40828
rect 25403 40826 25427 40828
rect 25483 40826 25507 40828
rect 25563 40826 25569 40828
rect 25323 40774 25325 40826
rect 25505 40774 25507 40826
rect 25261 40772 25267 40774
rect 25323 40772 25347 40774
rect 25403 40772 25427 40774
rect 25483 40772 25507 40774
rect 25563 40772 25569 40774
rect 25261 40763 25569 40772
rect 25261 39740 25569 39749
rect 25261 39738 25267 39740
rect 25323 39738 25347 39740
rect 25403 39738 25427 39740
rect 25483 39738 25507 39740
rect 25563 39738 25569 39740
rect 25323 39686 25325 39738
rect 25505 39686 25507 39738
rect 25261 39684 25267 39686
rect 25323 39684 25347 39686
rect 25403 39684 25427 39686
rect 25483 39684 25507 39686
rect 25563 39684 25569 39686
rect 25261 39675 25569 39684
rect 25261 38652 25569 38661
rect 25261 38650 25267 38652
rect 25323 38650 25347 38652
rect 25403 38650 25427 38652
rect 25483 38650 25507 38652
rect 25563 38650 25569 38652
rect 25323 38598 25325 38650
rect 25505 38598 25507 38650
rect 25261 38596 25267 38598
rect 25323 38596 25347 38598
rect 25403 38596 25427 38598
rect 25483 38596 25507 38598
rect 25563 38596 25569 38598
rect 25261 38587 25569 38596
rect 25261 37564 25569 37573
rect 25261 37562 25267 37564
rect 25323 37562 25347 37564
rect 25403 37562 25427 37564
rect 25483 37562 25507 37564
rect 25563 37562 25569 37564
rect 25323 37510 25325 37562
rect 25505 37510 25507 37562
rect 25261 37508 25267 37510
rect 25323 37508 25347 37510
rect 25403 37508 25427 37510
rect 25483 37508 25507 37510
rect 25563 37508 25569 37510
rect 25261 37499 25569 37508
rect 26068 37398 26096 42191
rect 26146 39536 26202 39545
rect 26146 39471 26202 39480
rect 26160 38894 26188 39471
rect 26148 38888 26200 38894
rect 26148 38830 26200 38836
rect 24768 37392 24820 37398
rect 24768 37334 24820 37340
rect 26056 37392 26108 37398
rect 26056 37334 26108 37340
rect 24780 37262 24808 37334
rect 26240 37324 26292 37330
rect 26240 37266 26292 37272
rect 23756 37256 23808 37262
rect 23756 37198 23808 37204
rect 24492 37256 24544 37262
rect 24492 37198 24544 37204
rect 24768 37256 24820 37262
rect 24768 37198 24820 37204
rect 23296 37120 23348 37126
rect 23348 37080 23520 37108
rect 23296 37062 23348 37068
rect 23492 36922 23520 37080
rect 23480 36916 23532 36922
rect 23480 36858 23532 36864
rect 23940 36916 23992 36922
rect 23940 36858 23992 36864
rect 23480 36780 23532 36786
rect 23480 36722 23532 36728
rect 23492 36106 23520 36722
rect 23952 36242 23980 36858
rect 23940 36236 23992 36242
rect 23940 36178 23992 36184
rect 23480 36100 23532 36106
rect 23480 36042 23532 36048
rect 23388 35012 23440 35018
rect 23388 34954 23440 34960
rect 23400 34066 23428 34954
rect 23952 34746 23980 36178
rect 24124 36100 24176 36106
rect 24124 36042 24176 36048
rect 23940 34740 23992 34746
rect 23940 34682 23992 34688
rect 23388 34060 23440 34066
rect 23388 34002 23440 34008
rect 23400 33454 23428 34002
rect 24136 33998 24164 36042
rect 23664 33992 23716 33998
rect 23664 33934 23716 33940
rect 23756 33992 23808 33998
rect 23756 33934 23808 33940
rect 24124 33992 24176 33998
rect 24124 33934 24176 33940
rect 23572 33856 23624 33862
rect 23572 33798 23624 33804
rect 23480 33516 23532 33522
rect 23480 33458 23532 33464
rect 23388 33448 23440 33454
rect 23388 33390 23440 33396
rect 23492 33114 23520 33458
rect 23480 33108 23532 33114
rect 23480 33050 23532 33056
rect 23480 32972 23532 32978
rect 23480 32914 23532 32920
rect 23112 32428 23164 32434
rect 23112 32370 23164 32376
rect 23124 32026 23152 32370
rect 22928 32020 22980 32026
rect 22928 31962 22980 31968
rect 23112 32020 23164 32026
rect 23112 31962 23164 31968
rect 22192 31816 22244 31822
rect 22192 31758 22244 31764
rect 21788 31580 22096 31589
rect 21788 31578 21794 31580
rect 21850 31578 21874 31580
rect 21930 31578 21954 31580
rect 22010 31578 22034 31580
rect 22090 31578 22096 31580
rect 21850 31526 21852 31578
rect 22032 31526 22034 31578
rect 21788 31524 21794 31526
rect 21850 31524 21874 31526
rect 21930 31524 21954 31526
rect 22010 31524 22034 31526
rect 22090 31524 22096 31526
rect 21788 31515 22096 31524
rect 22204 31482 22232 31758
rect 22560 31680 22612 31686
rect 22560 31622 22612 31628
rect 22192 31476 22244 31482
rect 22192 31418 22244 31424
rect 22468 31408 22520 31414
rect 22468 31350 22520 31356
rect 21640 31340 21692 31346
rect 21640 31282 21692 31288
rect 21652 30666 21680 31282
rect 22480 30734 22508 31350
rect 22572 31346 22600 31622
rect 22940 31414 22968 31962
rect 23204 31680 23256 31686
rect 23204 31622 23256 31628
rect 23216 31482 23244 31622
rect 23204 31476 23256 31482
rect 23204 31418 23256 31424
rect 22928 31408 22980 31414
rect 22928 31350 22980 31356
rect 22560 31340 22612 31346
rect 22560 31282 22612 31288
rect 22836 31340 22888 31346
rect 22836 31282 22888 31288
rect 23112 31340 23164 31346
rect 23112 31282 23164 31288
rect 22848 30938 22876 31282
rect 23124 30938 23152 31282
rect 23388 31272 23440 31278
rect 23388 31214 23440 31220
rect 22836 30932 22888 30938
rect 22836 30874 22888 30880
rect 23112 30932 23164 30938
rect 23112 30874 23164 30880
rect 23400 30734 23428 31214
rect 22468 30728 22520 30734
rect 22468 30670 22520 30676
rect 23388 30728 23440 30734
rect 23388 30670 23440 30676
rect 21640 30660 21692 30666
rect 21640 30602 21692 30608
rect 21652 30326 21680 30602
rect 21788 30492 22096 30501
rect 21788 30490 21794 30492
rect 21850 30490 21874 30492
rect 21930 30490 21954 30492
rect 22010 30490 22034 30492
rect 22090 30490 22096 30492
rect 21850 30438 21852 30490
rect 22032 30438 22034 30490
rect 21788 30436 21794 30438
rect 21850 30436 21874 30438
rect 21930 30436 21954 30438
rect 22010 30436 22034 30438
rect 22090 30436 22096 30438
rect 21788 30427 22096 30436
rect 21640 30320 21692 30326
rect 21640 30262 21692 30268
rect 21456 27600 21508 27606
rect 21456 27542 21508 27548
rect 21652 27130 21680 30262
rect 22480 30258 22508 30670
rect 23112 30592 23164 30598
rect 23112 30534 23164 30540
rect 22284 30252 22336 30258
rect 22284 30194 22336 30200
rect 22468 30252 22520 30258
rect 22468 30194 22520 30200
rect 22008 30048 22060 30054
rect 22008 29990 22060 29996
rect 22020 29578 22048 29990
rect 22008 29572 22060 29578
rect 22008 29514 22060 29520
rect 22192 29504 22244 29510
rect 22192 29446 22244 29452
rect 21788 29404 22096 29413
rect 21788 29402 21794 29404
rect 21850 29402 21874 29404
rect 21930 29402 21954 29404
rect 22010 29402 22034 29404
rect 22090 29402 22096 29404
rect 21850 29350 21852 29402
rect 22032 29350 22034 29402
rect 21788 29348 21794 29350
rect 21850 29348 21874 29350
rect 21930 29348 21954 29350
rect 22010 29348 22034 29350
rect 22090 29348 22096 29350
rect 21788 29339 22096 29348
rect 22204 29170 22232 29446
rect 22296 29306 22324 30194
rect 22744 30116 22796 30122
rect 22744 30058 22796 30064
rect 22652 29640 22704 29646
rect 22652 29582 22704 29588
rect 22284 29300 22336 29306
rect 22284 29242 22336 29248
rect 22192 29164 22244 29170
rect 22192 29106 22244 29112
rect 22284 29164 22336 29170
rect 22284 29106 22336 29112
rect 22192 29028 22244 29034
rect 22192 28970 22244 28976
rect 21788 28316 22096 28325
rect 21788 28314 21794 28316
rect 21850 28314 21874 28316
rect 21930 28314 21954 28316
rect 22010 28314 22034 28316
rect 22090 28314 22096 28316
rect 21850 28262 21852 28314
rect 22032 28262 22034 28314
rect 21788 28260 21794 28262
rect 21850 28260 21874 28262
rect 21930 28260 21954 28262
rect 22010 28260 22034 28262
rect 22090 28260 22096 28262
rect 21788 28251 22096 28260
rect 22204 28082 22232 28970
rect 22296 28082 22324 29106
rect 22664 28626 22692 29582
rect 22756 29102 22784 30058
rect 23124 29186 23152 30534
rect 23296 30320 23348 30326
rect 23296 30262 23348 30268
rect 23204 30184 23256 30190
rect 23204 30126 23256 30132
rect 23216 29306 23244 30126
rect 23308 30054 23336 30262
rect 23296 30048 23348 30054
rect 23296 29990 23348 29996
rect 23204 29300 23256 29306
rect 23204 29242 23256 29248
rect 23124 29170 23244 29186
rect 23124 29164 23256 29170
rect 23124 29158 23204 29164
rect 23204 29106 23256 29112
rect 22744 29096 22796 29102
rect 22744 29038 22796 29044
rect 22652 28620 22704 28626
rect 22652 28562 22704 28568
rect 22560 28552 22612 28558
rect 22560 28494 22612 28500
rect 22468 28484 22520 28490
rect 22468 28426 22520 28432
rect 22480 28218 22508 28426
rect 22468 28212 22520 28218
rect 22468 28154 22520 28160
rect 22192 28076 22244 28082
rect 22192 28018 22244 28024
rect 22284 28076 22336 28082
rect 22284 28018 22336 28024
rect 22204 27690 22232 28018
rect 22296 27826 22324 28018
rect 22296 27798 22416 27826
rect 22204 27662 22324 27690
rect 22192 27600 22244 27606
rect 22192 27542 22244 27548
rect 21788 27228 22096 27237
rect 21788 27226 21794 27228
rect 21850 27226 21874 27228
rect 21930 27226 21954 27228
rect 22010 27226 22034 27228
rect 22090 27226 22096 27228
rect 21850 27174 21852 27226
rect 22032 27174 22034 27226
rect 21788 27172 21794 27174
rect 21850 27172 21874 27174
rect 21930 27172 21954 27174
rect 22010 27172 22034 27174
rect 22090 27172 22096 27174
rect 21788 27163 22096 27172
rect 21640 27124 21692 27130
rect 21640 27066 21692 27072
rect 22008 26920 22060 26926
rect 22008 26862 22060 26868
rect 22020 26586 22048 26862
rect 22204 26858 22232 27542
rect 22296 27334 22324 27662
rect 22284 27328 22336 27334
rect 22284 27270 22336 27276
rect 22192 26852 22244 26858
rect 22192 26794 22244 26800
rect 22008 26580 22060 26586
rect 22008 26522 22060 26528
rect 21788 26140 22096 26149
rect 21788 26138 21794 26140
rect 21850 26138 21874 26140
rect 21930 26138 21954 26140
rect 22010 26138 22034 26140
rect 22090 26138 22096 26140
rect 21850 26086 21852 26138
rect 22032 26086 22034 26138
rect 21788 26084 21794 26086
rect 21850 26084 21874 26086
rect 21930 26084 21954 26086
rect 22010 26084 22034 26086
rect 22090 26084 22096 26086
rect 21788 26075 22096 26084
rect 21732 25696 21784 25702
rect 21732 25638 21784 25644
rect 21744 25294 21772 25638
rect 21456 25288 21508 25294
rect 21456 25230 21508 25236
rect 21732 25288 21784 25294
rect 21732 25230 21784 25236
rect 21192 23446 21312 23474
rect 21192 22778 21220 23446
rect 21180 22772 21232 22778
rect 21180 22714 21232 22720
rect 21272 22704 21324 22710
rect 21272 22646 21324 22652
rect 21284 21894 21312 22646
rect 21468 22030 21496 25230
rect 21788 25052 22096 25061
rect 21788 25050 21794 25052
rect 21850 25050 21874 25052
rect 21930 25050 21954 25052
rect 22010 25050 22034 25052
rect 22090 25050 22096 25052
rect 21850 24998 21852 25050
rect 22032 24998 22034 25050
rect 21788 24996 21794 24998
rect 21850 24996 21874 24998
rect 21930 24996 21954 24998
rect 22010 24996 22034 24998
rect 22090 24996 22096 24998
rect 21788 24987 22096 24996
rect 21548 24880 21600 24886
rect 21548 24822 21600 24828
rect 21456 22024 21508 22030
rect 21456 21966 21508 21972
rect 21272 21888 21324 21894
rect 21272 21830 21324 21836
rect 21180 19780 21232 19786
rect 21180 19722 21232 19728
rect 21192 19378 21220 19722
rect 21180 19372 21232 19378
rect 21180 19314 21232 19320
rect 20996 15564 21048 15570
rect 20996 15506 21048 15512
rect 20812 14612 20864 14618
rect 20812 14554 20864 14560
rect 20824 12238 20852 14554
rect 21192 12434 21220 19314
rect 21284 16658 21312 21830
rect 21456 19848 21508 19854
rect 21456 19790 21508 19796
rect 21468 18426 21496 19790
rect 21456 18420 21508 18426
rect 21456 18362 21508 18368
rect 21468 17610 21496 18362
rect 21456 17604 21508 17610
rect 21456 17546 21508 17552
rect 21272 16652 21324 16658
rect 21272 16594 21324 16600
rect 21560 15502 21588 24822
rect 21640 24812 21692 24818
rect 21640 24754 21692 24760
rect 21652 24410 21680 24754
rect 21640 24404 21692 24410
rect 21640 24346 21692 24352
rect 21788 23964 22096 23973
rect 21788 23962 21794 23964
rect 21850 23962 21874 23964
rect 21930 23962 21954 23964
rect 22010 23962 22034 23964
rect 22090 23962 22096 23964
rect 21850 23910 21852 23962
rect 22032 23910 22034 23962
rect 21788 23908 21794 23910
rect 21850 23908 21874 23910
rect 21930 23908 21954 23910
rect 22010 23908 22034 23910
rect 22090 23908 22096 23910
rect 21788 23899 22096 23908
rect 21640 23656 21692 23662
rect 21640 23598 21692 23604
rect 21652 22574 21680 23598
rect 21788 22876 22096 22885
rect 21788 22874 21794 22876
rect 21850 22874 21874 22876
rect 21930 22874 21954 22876
rect 22010 22874 22034 22876
rect 22090 22874 22096 22876
rect 21850 22822 21852 22874
rect 22032 22822 22034 22874
rect 21788 22820 21794 22822
rect 21850 22820 21874 22822
rect 21930 22820 21954 22822
rect 22010 22820 22034 22822
rect 22090 22820 22096 22822
rect 21788 22811 22096 22820
rect 21640 22568 21692 22574
rect 21640 22510 21692 22516
rect 21652 21010 21680 22510
rect 21788 21788 22096 21797
rect 21788 21786 21794 21788
rect 21850 21786 21874 21788
rect 21930 21786 21954 21788
rect 22010 21786 22034 21788
rect 22090 21786 22096 21788
rect 21850 21734 21852 21786
rect 22032 21734 22034 21786
rect 21788 21732 21794 21734
rect 21850 21732 21874 21734
rect 21930 21732 21954 21734
rect 22010 21732 22034 21734
rect 22090 21732 22096 21734
rect 21788 21723 22096 21732
rect 22008 21480 22060 21486
rect 22008 21422 22060 21428
rect 21640 21004 21692 21010
rect 21640 20946 21692 20952
rect 21652 19836 21680 20946
rect 22020 20806 22048 21422
rect 22008 20800 22060 20806
rect 22008 20742 22060 20748
rect 21788 20700 22096 20709
rect 21788 20698 21794 20700
rect 21850 20698 21874 20700
rect 21930 20698 21954 20700
rect 22010 20698 22034 20700
rect 22090 20698 22096 20700
rect 21850 20646 21852 20698
rect 22032 20646 22034 20698
rect 21788 20644 21794 20646
rect 21850 20644 21874 20646
rect 21930 20644 21954 20646
rect 22010 20644 22034 20646
rect 22090 20644 22096 20646
rect 21788 20635 22096 20644
rect 21824 19848 21876 19854
rect 21652 19808 21824 19836
rect 21824 19790 21876 19796
rect 21788 19612 22096 19621
rect 21788 19610 21794 19612
rect 21850 19610 21874 19612
rect 21930 19610 21954 19612
rect 22010 19610 22034 19612
rect 22090 19610 22096 19612
rect 21850 19558 21852 19610
rect 22032 19558 22034 19610
rect 21788 19556 21794 19558
rect 21850 19556 21874 19558
rect 21930 19556 21954 19558
rect 22010 19556 22034 19558
rect 22090 19556 22096 19558
rect 21788 19547 22096 19556
rect 22100 19372 22152 19378
rect 22100 19314 22152 19320
rect 22112 18834 22140 19314
rect 22100 18828 22152 18834
rect 22100 18770 22152 18776
rect 21788 18524 22096 18533
rect 21788 18522 21794 18524
rect 21850 18522 21874 18524
rect 21930 18522 21954 18524
rect 22010 18522 22034 18524
rect 22090 18522 22096 18524
rect 21850 18470 21852 18522
rect 22032 18470 22034 18522
rect 21788 18468 21794 18470
rect 21850 18468 21874 18470
rect 21930 18468 21954 18470
rect 22010 18468 22034 18470
rect 22090 18468 22096 18470
rect 21788 18459 22096 18468
rect 22204 18290 22232 26794
rect 22296 19446 22324 27270
rect 22388 26926 22416 27798
rect 22376 26920 22428 26926
rect 22428 26880 22508 26908
rect 22376 26862 22428 26868
rect 22376 25424 22428 25430
rect 22376 25366 22428 25372
rect 22388 24206 22416 25366
rect 22480 24818 22508 26880
rect 22572 25158 22600 28494
rect 22652 28416 22704 28422
rect 22652 28358 22704 28364
rect 22664 25906 22692 28358
rect 22756 26926 22784 29038
rect 23216 28422 23244 29106
rect 23204 28416 23256 28422
rect 23204 28358 23256 28364
rect 23204 27396 23256 27402
rect 23204 27338 23256 27344
rect 23216 27130 23244 27338
rect 23204 27124 23256 27130
rect 23204 27066 23256 27072
rect 22928 27056 22980 27062
rect 22928 26998 22980 27004
rect 22744 26920 22796 26926
rect 22744 26862 22796 26868
rect 22652 25900 22704 25906
rect 22652 25842 22704 25848
rect 22560 25152 22612 25158
rect 22560 25094 22612 25100
rect 22468 24812 22520 24818
rect 22468 24754 22520 24760
rect 22376 24200 22428 24206
rect 22376 24142 22428 24148
rect 22480 24018 22508 24754
rect 22388 23990 22508 24018
rect 22388 21554 22416 23990
rect 22468 22432 22520 22438
rect 22468 22374 22520 22380
rect 22480 22030 22508 22374
rect 22468 22024 22520 22030
rect 22468 21966 22520 21972
rect 22376 21548 22428 21554
rect 22376 21490 22428 21496
rect 22388 19786 22416 21490
rect 22468 19848 22520 19854
rect 22468 19790 22520 19796
rect 22376 19780 22428 19786
rect 22376 19722 22428 19728
rect 22284 19440 22336 19446
rect 22284 19382 22336 19388
rect 22296 18834 22324 19382
rect 22284 18828 22336 18834
rect 22284 18770 22336 18776
rect 22192 18284 22244 18290
rect 22192 18226 22244 18232
rect 22296 18222 22324 18770
rect 22388 18698 22416 19722
rect 22480 19514 22508 19790
rect 22468 19508 22520 19514
rect 22468 19450 22520 19456
rect 22376 18692 22428 18698
rect 22376 18634 22428 18640
rect 22284 18216 22336 18222
rect 22284 18158 22336 18164
rect 22480 18170 22508 19450
rect 22572 18358 22600 25094
rect 22664 22642 22692 25842
rect 22756 24750 22784 26862
rect 22940 26042 22968 26998
rect 23308 26994 23336 29990
rect 23400 28558 23428 30670
rect 23492 29170 23520 32914
rect 23584 32910 23612 33798
rect 23676 32910 23704 33934
rect 23768 33318 23796 33934
rect 24136 33590 24164 33934
rect 24124 33584 24176 33590
rect 24124 33526 24176 33532
rect 23756 33312 23808 33318
rect 23756 33254 23808 33260
rect 23768 32978 23796 33254
rect 23756 32972 23808 32978
rect 23756 32914 23808 32920
rect 23572 32904 23624 32910
rect 23572 32846 23624 32852
rect 23664 32904 23716 32910
rect 23664 32846 23716 32852
rect 23664 32224 23716 32230
rect 23664 32166 23716 32172
rect 23676 31890 23704 32166
rect 23664 31884 23716 31890
rect 23664 31826 23716 31832
rect 23572 31816 23624 31822
rect 23572 31758 23624 31764
rect 23584 31482 23612 31758
rect 23940 31748 23992 31754
rect 23940 31690 23992 31696
rect 23572 31476 23624 31482
rect 23572 31418 23624 31424
rect 23584 30734 23612 31418
rect 23952 31346 23980 31690
rect 23940 31340 23992 31346
rect 23940 31282 23992 31288
rect 23952 30802 23980 31282
rect 23940 30796 23992 30802
rect 23940 30738 23992 30744
rect 23572 30728 23624 30734
rect 23572 30670 23624 30676
rect 23664 30660 23716 30666
rect 23664 30602 23716 30608
rect 23756 30660 23808 30666
rect 23756 30602 23808 30608
rect 23676 30122 23704 30602
rect 23664 30116 23716 30122
rect 23664 30058 23716 30064
rect 23676 29306 23704 30058
rect 23768 30054 23796 30602
rect 23756 30048 23808 30054
rect 23756 29990 23808 29996
rect 23768 29782 23796 29990
rect 23756 29776 23808 29782
rect 23756 29718 23808 29724
rect 23664 29300 23716 29306
rect 23664 29242 23716 29248
rect 23480 29164 23532 29170
rect 23480 29106 23532 29112
rect 23388 28552 23440 28558
rect 23388 28494 23440 28500
rect 23400 28218 23428 28494
rect 23388 28212 23440 28218
rect 23388 28154 23440 28160
rect 23296 26988 23348 26994
rect 23296 26930 23348 26936
rect 22928 26036 22980 26042
rect 22928 25978 22980 25984
rect 22836 25288 22888 25294
rect 22836 25230 22888 25236
rect 22848 24818 22876 25230
rect 22836 24812 22888 24818
rect 22836 24754 22888 24760
rect 22744 24744 22796 24750
rect 22744 24686 22796 24692
rect 22652 22636 22704 22642
rect 22652 22578 22704 22584
rect 22756 21486 22784 24686
rect 22928 22024 22980 22030
rect 22928 21966 22980 21972
rect 22940 21690 22968 21966
rect 23112 21888 23164 21894
rect 23112 21830 23164 21836
rect 22928 21684 22980 21690
rect 22928 21626 22980 21632
rect 22744 21480 22796 21486
rect 22744 21422 22796 21428
rect 23124 20942 23152 21830
rect 23112 20936 23164 20942
rect 23112 20878 23164 20884
rect 23204 19712 23256 19718
rect 23204 19654 23256 19660
rect 23216 19446 23244 19654
rect 23204 19440 23256 19446
rect 23204 19382 23256 19388
rect 23308 18902 23336 26930
rect 23388 24200 23440 24206
rect 23388 24142 23440 24148
rect 23400 22710 23428 24142
rect 23492 24138 23520 29106
rect 23756 28960 23808 28966
rect 23756 28902 23808 28908
rect 23768 28150 23796 28902
rect 23952 28490 23980 30738
rect 24032 29708 24084 29714
rect 24032 29650 24084 29656
rect 23940 28484 23992 28490
rect 23940 28426 23992 28432
rect 23664 28144 23716 28150
rect 23664 28086 23716 28092
rect 23756 28144 23808 28150
rect 23756 28086 23808 28092
rect 23676 26994 23704 28086
rect 23768 27062 23796 28086
rect 23756 27056 23808 27062
rect 23756 26998 23808 27004
rect 23664 26988 23716 26994
rect 23664 26930 23716 26936
rect 23952 26382 23980 28426
rect 24044 26586 24072 29650
rect 24136 28082 24164 33526
rect 24216 32768 24268 32774
rect 24216 32710 24268 32716
rect 24228 31414 24256 32710
rect 24308 31952 24360 31958
rect 24308 31894 24360 31900
rect 24216 31408 24268 31414
rect 24216 31350 24268 31356
rect 24216 30388 24268 30394
rect 24216 30330 24268 30336
rect 24228 30258 24256 30330
rect 24216 30252 24268 30258
rect 24216 30194 24268 30200
rect 24320 30122 24348 31894
rect 24308 30116 24360 30122
rect 24308 30058 24360 30064
rect 24320 28098 24348 30058
rect 24504 28506 24532 37198
rect 26056 37188 26108 37194
rect 26056 37130 26108 37136
rect 26068 36922 26096 37130
rect 26056 36916 26108 36922
rect 26056 36858 26108 36864
rect 25964 36780 26016 36786
rect 25964 36722 26016 36728
rect 25261 36476 25569 36485
rect 25261 36474 25267 36476
rect 25323 36474 25347 36476
rect 25403 36474 25427 36476
rect 25483 36474 25507 36476
rect 25563 36474 25569 36476
rect 25323 36422 25325 36474
rect 25505 36422 25507 36474
rect 25261 36420 25267 36422
rect 25323 36420 25347 36422
rect 25403 36420 25427 36422
rect 25483 36420 25507 36422
rect 25563 36420 25569 36422
rect 25261 36411 25569 36420
rect 25688 35624 25740 35630
rect 25688 35566 25740 35572
rect 24952 35488 25004 35494
rect 24952 35430 25004 35436
rect 24860 34740 24912 34746
rect 24860 34682 24912 34688
rect 24872 33114 24900 34682
rect 24964 33998 24992 35430
rect 25261 35388 25569 35397
rect 25261 35386 25267 35388
rect 25323 35386 25347 35388
rect 25403 35386 25427 35388
rect 25483 35386 25507 35388
rect 25563 35386 25569 35388
rect 25323 35334 25325 35386
rect 25505 35334 25507 35386
rect 25261 35332 25267 35334
rect 25323 35332 25347 35334
rect 25403 35332 25427 35334
rect 25483 35332 25507 35334
rect 25563 35332 25569 35334
rect 25261 35323 25569 35332
rect 25044 34944 25096 34950
rect 25044 34886 25096 34892
rect 24952 33992 25004 33998
rect 24952 33934 25004 33940
rect 25056 33658 25084 34886
rect 25700 34746 25728 35566
rect 25688 34740 25740 34746
rect 25688 34682 25740 34688
rect 25261 34300 25569 34309
rect 25261 34298 25267 34300
rect 25323 34298 25347 34300
rect 25403 34298 25427 34300
rect 25483 34298 25507 34300
rect 25563 34298 25569 34300
rect 25323 34246 25325 34298
rect 25505 34246 25507 34298
rect 25261 34244 25267 34246
rect 25323 34244 25347 34246
rect 25403 34244 25427 34246
rect 25483 34244 25507 34246
rect 25563 34244 25569 34246
rect 25261 34235 25569 34244
rect 25136 33924 25188 33930
rect 25136 33866 25188 33872
rect 25044 33652 25096 33658
rect 25044 33594 25096 33600
rect 24860 33108 24912 33114
rect 24860 33050 24912 33056
rect 25044 32836 25096 32842
rect 25044 32778 25096 32784
rect 24952 31748 25004 31754
rect 24952 31690 25004 31696
rect 24964 30938 24992 31690
rect 24952 30932 25004 30938
rect 24952 30874 25004 30880
rect 24860 30728 24912 30734
rect 24860 30670 24912 30676
rect 24584 30592 24636 30598
rect 24584 30534 24636 30540
rect 24768 30592 24820 30598
rect 24768 30534 24820 30540
rect 24596 30258 24624 30534
rect 24584 30252 24636 30258
rect 24584 30194 24636 30200
rect 24596 29646 24624 30194
rect 24780 30190 24808 30534
rect 24872 30326 24900 30670
rect 24860 30320 24912 30326
rect 24860 30262 24912 30268
rect 24768 30184 24820 30190
rect 24768 30126 24820 30132
rect 24952 30048 25004 30054
rect 24952 29990 25004 29996
rect 24964 29850 24992 29990
rect 24952 29844 25004 29850
rect 24952 29786 25004 29792
rect 24584 29640 24636 29646
rect 25056 29594 25084 32778
rect 25148 30666 25176 33866
rect 25780 33856 25832 33862
rect 25780 33798 25832 33804
rect 25872 33856 25924 33862
rect 25872 33798 25924 33804
rect 25261 33212 25569 33221
rect 25261 33210 25267 33212
rect 25323 33210 25347 33212
rect 25403 33210 25427 33212
rect 25483 33210 25507 33212
rect 25563 33210 25569 33212
rect 25323 33158 25325 33210
rect 25505 33158 25507 33210
rect 25261 33156 25267 33158
rect 25323 33156 25347 33158
rect 25403 33156 25427 33158
rect 25483 33156 25507 33158
rect 25563 33156 25569 33158
rect 25261 33147 25569 33156
rect 25261 32124 25569 32133
rect 25261 32122 25267 32124
rect 25323 32122 25347 32124
rect 25403 32122 25427 32124
rect 25483 32122 25507 32124
rect 25563 32122 25569 32124
rect 25323 32070 25325 32122
rect 25505 32070 25507 32122
rect 25261 32068 25267 32070
rect 25323 32068 25347 32070
rect 25403 32068 25427 32070
rect 25483 32068 25507 32070
rect 25563 32068 25569 32070
rect 25261 32059 25569 32068
rect 25792 31890 25820 33798
rect 25884 32910 25912 33798
rect 25872 32904 25924 32910
rect 25872 32846 25924 32852
rect 25976 32756 26004 36722
rect 26252 35894 26280 37266
rect 26344 37126 26372 47382
rect 26608 47048 26660 47054
rect 26608 46990 26660 46996
rect 27344 47048 27396 47054
rect 27344 46990 27396 46996
rect 26424 46980 26476 46986
rect 26424 46922 26476 46928
rect 26436 46714 26464 46922
rect 26424 46708 26476 46714
rect 26424 46650 26476 46656
rect 26620 46510 26648 46990
rect 26608 46504 26660 46510
rect 26608 46446 26660 46452
rect 26516 46368 26568 46374
rect 26516 46310 26568 46316
rect 27252 46368 27304 46374
rect 27252 46310 27304 46316
rect 26528 46034 26556 46310
rect 26516 46028 26568 46034
rect 26516 45970 26568 45976
rect 27264 45558 27292 46310
rect 27252 45552 27304 45558
rect 27252 45494 27304 45500
rect 27356 45286 27384 46990
rect 27436 46572 27488 46578
rect 27436 46514 27488 46520
rect 27448 46102 27476 46514
rect 27526 46336 27582 46345
rect 27526 46271 27582 46280
rect 27436 46096 27488 46102
rect 27436 46038 27488 46044
rect 27344 45280 27396 45286
rect 27344 45222 27396 45228
rect 27160 44396 27212 44402
rect 27160 44338 27212 44344
rect 26424 44192 26476 44198
rect 26424 44134 26476 44140
rect 26436 43858 26464 44134
rect 26424 43852 26476 43858
rect 26424 43794 26476 43800
rect 27172 43314 27200 44338
rect 27160 43308 27212 43314
rect 27160 43250 27212 43256
rect 26700 43104 26752 43110
rect 26700 43046 26752 43052
rect 27160 43104 27212 43110
rect 27160 43046 27212 43052
rect 26712 42634 26740 43046
rect 27172 42770 27200 43046
rect 27160 42764 27212 42770
rect 27160 42706 27212 42712
rect 26700 42628 26752 42634
rect 26700 42570 26752 42576
rect 27448 41138 27476 46038
rect 27540 44946 27568 46271
rect 27724 46034 27752 49200
rect 28262 47696 28318 47705
rect 28262 47631 28318 47640
rect 27896 47048 27948 47054
rect 27896 46990 27948 46996
rect 27712 46028 27764 46034
rect 27712 45970 27764 45976
rect 27712 45620 27764 45626
rect 27712 45562 27764 45568
rect 27528 44940 27580 44946
rect 27528 44882 27580 44888
rect 27724 42226 27752 45562
rect 27908 45490 27936 46990
rect 27896 45484 27948 45490
rect 27896 45426 27948 45432
rect 27988 45348 28040 45354
rect 27988 45290 28040 45296
rect 27896 44804 27948 44810
rect 27896 44746 27948 44752
rect 27908 44538 27936 44746
rect 27896 44532 27948 44538
rect 27896 44474 27948 44480
rect 28000 44402 28028 45290
rect 28078 44976 28134 44985
rect 28078 44911 28134 44920
rect 27988 44396 28040 44402
rect 27988 44338 28040 44344
rect 27712 42220 27764 42226
rect 27712 42162 27764 42168
rect 27528 41676 27580 41682
rect 27528 41618 27580 41624
rect 27540 41585 27568 41618
rect 27526 41576 27582 41585
rect 27526 41511 27582 41520
rect 27436 41132 27488 41138
rect 27436 41074 27488 41080
rect 26516 39840 26568 39846
rect 26516 39782 26568 39788
rect 26528 39506 26556 39782
rect 26516 39500 26568 39506
rect 26516 39442 26568 39448
rect 26516 38344 26568 38350
rect 26516 38286 26568 38292
rect 26528 37874 26556 38286
rect 26700 38276 26752 38282
rect 26700 38218 26752 38224
rect 26516 37868 26568 37874
rect 26516 37810 26568 37816
rect 26332 37120 26384 37126
rect 26332 37062 26384 37068
rect 26712 36922 26740 38218
rect 26700 36916 26752 36922
rect 26700 36858 26752 36864
rect 26976 36780 27028 36786
rect 26976 36722 27028 36728
rect 26700 36100 26752 36106
rect 26700 36042 26752 36048
rect 26252 35866 26372 35894
rect 26240 35488 26292 35494
rect 26240 35430 26292 35436
rect 26252 35018 26280 35430
rect 26240 35012 26292 35018
rect 26240 34954 26292 34960
rect 26344 33522 26372 35866
rect 26712 35834 26740 36042
rect 26988 35894 27016 36722
rect 27448 35894 27476 41074
rect 27526 40624 27582 40633
rect 27526 40559 27528 40568
rect 27580 40559 27582 40568
rect 27528 40530 27580 40536
rect 27528 39840 27580 39846
rect 27528 39782 27580 39788
rect 27540 38962 27568 39782
rect 27896 39364 27948 39370
rect 27896 39306 27948 39312
rect 27528 38956 27580 38962
rect 27528 38898 27580 38904
rect 27712 38956 27764 38962
rect 27712 38898 27764 38904
rect 27724 38418 27752 38898
rect 27712 38412 27764 38418
rect 27712 38354 27764 38360
rect 27908 38010 27936 39306
rect 27896 38004 27948 38010
rect 27896 37946 27948 37952
rect 27804 37868 27856 37874
rect 27804 37810 27856 37816
rect 27816 36854 27844 37810
rect 27804 36848 27856 36854
rect 27804 36790 27856 36796
rect 27896 36576 27948 36582
rect 27896 36518 27948 36524
rect 27804 36304 27856 36310
rect 27804 36246 27856 36252
rect 27816 35894 27844 36246
rect 27908 36242 27936 36518
rect 27896 36236 27948 36242
rect 27896 36178 27948 36184
rect 28000 35894 28028 44338
rect 28092 43858 28120 44911
rect 28080 43852 28132 43858
rect 28080 43794 28132 43800
rect 28080 43104 28132 43110
rect 28080 43046 28132 43052
rect 28092 41750 28120 43046
rect 28172 42016 28224 42022
rect 28172 41958 28224 41964
rect 28080 41744 28132 41750
rect 28080 41686 28132 41692
rect 28184 41682 28212 41958
rect 28172 41676 28224 41682
rect 28172 41618 28224 41624
rect 28172 40928 28224 40934
rect 28172 40870 28224 40876
rect 28184 40594 28212 40870
rect 28172 40588 28224 40594
rect 28172 40530 28224 40536
rect 28276 38418 28304 47631
rect 28368 47122 28396 49200
rect 28356 47116 28408 47122
rect 28356 47058 28408 47064
rect 28734 46812 29042 46821
rect 28734 46810 28740 46812
rect 28796 46810 28820 46812
rect 28876 46810 28900 46812
rect 28956 46810 28980 46812
rect 29036 46810 29042 46812
rect 28796 46758 28798 46810
rect 28978 46758 28980 46810
rect 28734 46756 28740 46758
rect 28796 46756 28820 46758
rect 28876 46756 28900 46758
rect 28956 46756 28980 46758
rect 29036 46756 29042 46758
rect 28734 46747 29042 46756
rect 28540 46436 28592 46442
rect 28540 46378 28592 46384
rect 28356 45280 28408 45286
rect 28356 45222 28408 45228
rect 28368 44946 28396 45222
rect 28356 44940 28408 44946
rect 28356 44882 28408 44888
rect 28354 42936 28410 42945
rect 28354 42871 28410 42880
rect 28368 42770 28396 42871
rect 28356 42764 28408 42770
rect 28356 42706 28408 42712
rect 28356 40928 28408 40934
rect 28356 40870 28408 40876
rect 28368 40594 28396 40870
rect 28356 40588 28408 40594
rect 28356 40530 28408 40536
rect 28264 38412 28316 38418
rect 28264 38354 28316 38360
rect 28356 37256 28408 37262
rect 28356 37198 28408 37204
rect 28172 37120 28224 37126
rect 28172 37062 28224 37068
rect 26896 35866 27016 35894
rect 27172 35866 27476 35894
rect 27632 35866 27844 35894
rect 27908 35866 28028 35894
rect 26700 35828 26752 35834
rect 26700 35770 26752 35776
rect 26896 35766 26924 35866
rect 26884 35760 26936 35766
rect 26884 35702 26936 35708
rect 26608 34944 26660 34950
rect 26608 34886 26660 34892
rect 26620 34610 26648 34886
rect 26608 34604 26660 34610
rect 26608 34546 26660 34552
rect 26332 33516 26384 33522
rect 26332 33458 26384 33464
rect 25884 32728 26004 32756
rect 25884 32434 25912 32728
rect 25872 32428 25924 32434
rect 25872 32370 25924 32376
rect 25884 32026 25912 32370
rect 25964 32224 26016 32230
rect 25964 32166 26016 32172
rect 26608 32224 26660 32230
rect 26608 32166 26660 32172
rect 25872 32020 25924 32026
rect 25872 31962 25924 31968
rect 25976 31890 26004 32166
rect 25780 31884 25832 31890
rect 25780 31826 25832 31832
rect 25964 31884 26016 31890
rect 25964 31826 26016 31832
rect 26620 31346 26648 32166
rect 26608 31340 26660 31346
rect 26608 31282 26660 31288
rect 26148 31272 26200 31278
rect 26148 31214 26200 31220
rect 25261 31036 25569 31045
rect 25261 31034 25267 31036
rect 25323 31034 25347 31036
rect 25403 31034 25427 31036
rect 25483 31034 25507 31036
rect 25563 31034 25569 31036
rect 25323 30982 25325 31034
rect 25505 30982 25507 31034
rect 25261 30980 25267 30982
rect 25323 30980 25347 30982
rect 25403 30980 25427 30982
rect 25483 30980 25507 30982
rect 25563 30980 25569 30982
rect 25261 30971 25569 30980
rect 26160 30705 26188 31214
rect 26332 30728 26384 30734
rect 26146 30696 26202 30705
rect 25136 30660 25188 30666
rect 26332 30670 26384 30676
rect 26146 30631 26202 30640
rect 25136 30602 25188 30608
rect 25964 30252 26016 30258
rect 25964 30194 26016 30200
rect 26148 30252 26200 30258
rect 26148 30194 26200 30200
rect 25261 29948 25569 29957
rect 25261 29946 25267 29948
rect 25323 29946 25347 29948
rect 25403 29946 25427 29948
rect 25483 29946 25507 29948
rect 25563 29946 25569 29948
rect 25323 29894 25325 29946
rect 25505 29894 25507 29946
rect 25261 29892 25267 29894
rect 25323 29892 25347 29894
rect 25403 29892 25427 29894
rect 25483 29892 25507 29894
rect 25563 29892 25569 29894
rect 25261 29883 25569 29892
rect 24584 29582 24636 29588
rect 24964 29566 25084 29594
rect 25872 29640 25924 29646
rect 25872 29582 25924 29588
rect 24964 29170 24992 29566
rect 25044 29504 25096 29510
rect 25044 29446 25096 29452
rect 24952 29164 25004 29170
rect 24952 29106 25004 29112
rect 24858 29064 24914 29073
rect 24858 28999 24914 29008
rect 24676 28756 24728 28762
rect 24676 28698 24728 28704
rect 24504 28478 24624 28506
rect 24492 28416 24544 28422
rect 24492 28358 24544 28364
rect 24124 28076 24176 28082
rect 24320 28070 24440 28098
rect 24504 28082 24532 28358
rect 24124 28018 24176 28024
rect 24412 28014 24440 28070
rect 24492 28076 24544 28082
rect 24492 28018 24544 28024
rect 24400 28008 24452 28014
rect 24400 27950 24452 27956
rect 24492 27872 24544 27878
rect 24492 27814 24544 27820
rect 24504 27674 24532 27814
rect 24492 27668 24544 27674
rect 24492 27610 24544 27616
rect 24504 27130 24532 27610
rect 24492 27124 24544 27130
rect 24492 27066 24544 27072
rect 24124 26988 24176 26994
rect 24124 26930 24176 26936
rect 24492 26988 24544 26994
rect 24492 26930 24544 26936
rect 24032 26580 24084 26586
rect 24032 26522 24084 26528
rect 24136 26518 24164 26930
rect 24124 26512 24176 26518
rect 24124 26454 24176 26460
rect 24136 26382 24164 26454
rect 23940 26376 23992 26382
rect 23940 26318 23992 26324
rect 24124 26376 24176 26382
rect 24124 26318 24176 26324
rect 23664 25764 23716 25770
rect 23664 25706 23716 25712
rect 23676 24138 23704 25706
rect 23756 24404 23808 24410
rect 23756 24346 23808 24352
rect 23480 24132 23532 24138
rect 23480 24074 23532 24080
rect 23664 24132 23716 24138
rect 23664 24074 23716 24080
rect 23492 22982 23520 24074
rect 23572 23248 23624 23254
rect 23572 23190 23624 23196
rect 23480 22976 23532 22982
rect 23480 22918 23532 22924
rect 23388 22704 23440 22710
rect 23388 22646 23440 22652
rect 23400 21010 23428 22646
rect 23584 22506 23612 23190
rect 23676 23118 23704 24074
rect 23664 23112 23716 23118
rect 23664 23054 23716 23060
rect 23768 23050 23796 24346
rect 23756 23044 23808 23050
rect 23756 22986 23808 22992
rect 23768 22642 23796 22986
rect 23952 22642 23980 26318
rect 24032 24812 24084 24818
rect 24032 24754 24084 24760
rect 24044 24070 24072 24754
rect 24136 24682 24164 26318
rect 24216 25220 24268 25226
rect 24216 25162 24268 25168
rect 24124 24676 24176 24682
rect 24124 24618 24176 24624
rect 24032 24064 24084 24070
rect 24032 24006 24084 24012
rect 24044 22642 24072 24006
rect 23756 22636 23808 22642
rect 23756 22578 23808 22584
rect 23940 22636 23992 22642
rect 23940 22578 23992 22584
rect 24032 22636 24084 22642
rect 24032 22578 24084 22584
rect 23572 22500 23624 22506
rect 23572 22442 23624 22448
rect 23768 22094 23796 22578
rect 23848 22432 23900 22438
rect 23848 22374 23900 22380
rect 23676 22066 23796 22094
rect 23676 21554 23704 22066
rect 23860 22030 23888 22374
rect 23952 22234 23980 22578
rect 24124 22568 24176 22574
rect 24124 22510 24176 22516
rect 23940 22228 23992 22234
rect 23940 22170 23992 22176
rect 23848 22024 23900 22030
rect 23848 21966 23900 21972
rect 24136 21554 24164 22510
rect 24228 22030 24256 25162
rect 24308 22636 24360 22642
rect 24308 22578 24360 22584
rect 24216 22024 24268 22030
rect 24216 21966 24268 21972
rect 23664 21548 23716 21554
rect 23664 21490 23716 21496
rect 24124 21548 24176 21554
rect 24124 21490 24176 21496
rect 24032 21344 24084 21350
rect 24032 21286 24084 21292
rect 23388 21004 23440 21010
rect 23388 20946 23440 20952
rect 23400 20754 23428 20946
rect 23400 20726 23520 20754
rect 23492 20398 23520 20726
rect 23480 20392 23532 20398
rect 23480 20334 23532 20340
rect 23492 19378 23520 20334
rect 23480 19372 23532 19378
rect 23480 19314 23532 19320
rect 23296 18896 23348 18902
rect 23296 18838 23348 18844
rect 23204 18828 23256 18834
rect 23204 18770 23256 18776
rect 22560 18352 22612 18358
rect 22560 18294 22612 18300
rect 22480 18142 22600 18170
rect 22284 17536 22336 17542
rect 22284 17478 22336 17484
rect 21788 17436 22096 17445
rect 21788 17434 21794 17436
rect 21850 17434 21874 17436
rect 21930 17434 21954 17436
rect 22010 17434 22034 17436
rect 22090 17434 22096 17436
rect 21850 17382 21852 17434
rect 22032 17382 22034 17434
rect 21788 17380 21794 17382
rect 21850 17380 21874 17382
rect 21930 17380 21954 17382
rect 22010 17380 22034 17382
rect 22090 17380 22096 17382
rect 21788 17371 22096 17380
rect 22192 17196 22244 17202
rect 22192 17138 22244 17144
rect 21788 16348 22096 16357
rect 21788 16346 21794 16348
rect 21850 16346 21874 16348
rect 21930 16346 21954 16348
rect 22010 16346 22034 16348
rect 22090 16346 22096 16348
rect 21850 16294 21852 16346
rect 22032 16294 22034 16346
rect 21788 16292 21794 16294
rect 21850 16292 21874 16294
rect 21930 16292 21954 16294
rect 22010 16292 22034 16294
rect 22090 16292 22096 16294
rect 21788 16283 22096 16292
rect 22204 16250 22232 17138
rect 22192 16244 22244 16250
rect 22192 16186 22244 16192
rect 21548 15496 21600 15502
rect 21548 15438 21600 15444
rect 21788 15260 22096 15269
rect 21788 15258 21794 15260
rect 21850 15258 21874 15260
rect 21930 15258 21954 15260
rect 22010 15258 22034 15260
rect 22090 15258 22096 15260
rect 21850 15206 21852 15258
rect 22032 15206 22034 15258
rect 21788 15204 21794 15206
rect 21850 15204 21874 15206
rect 21930 15204 21954 15206
rect 22010 15204 22034 15206
rect 22090 15204 22096 15206
rect 21788 15195 22096 15204
rect 21272 14408 21324 14414
rect 21272 14350 21324 14356
rect 21284 13938 21312 14350
rect 21548 14340 21600 14346
rect 21548 14282 21600 14288
rect 21272 13932 21324 13938
rect 21272 13874 21324 13880
rect 21560 12442 21588 14282
rect 21788 14172 22096 14181
rect 21788 14170 21794 14172
rect 21850 14170 21874 14172
rect 21930 14170 21954 14172
rect 22010 14170 22034 14172
rect 22090 14170 22096 14172
rect 21850 14118 21852 14170
rect 22032 14118 22034 14170
rect 21788 14116 21794 14118
rect 21850 14116 21874 14118
rect 21930 14116 21954 14118
rect 22010 14116 22034 14118
rect 22090 14116 22096 14118
rect 21788 14107 22096 14116
rect 21640 14000 21692 14006
rect 21640 13942 21692 13948
rect 21548 12436 21600 12442
rect 21192 12406 21404 12434
rect 20996 12300 21048 12306
rect 20996 12242 21048 12248
rect 20812 12232 20864 12238
rect 20812 12174 20864 12180
rect 20444 11892 20496 11898
rect 20444 11834 20496 11840
rect 20352 11756 20404 11762
rect 20352 11698 20404 11704
rect 21008 11694 21036 12242
rect 21088 12232 21140 12238
rect 21088 12174 21140 12180
rect 19800 11688 19852 11694
rect 19800 11630 19852 11636
rect 20996 11688 21048 11694
rect 20996 11630 21048 11636
rect 19708 11552 19760 11558
rect 19708 11494 19760 11500
rect 19616 11348 19668 11354
rect 19616 11290 19668 11296
rect 19536 11206 19656 11234
rect 18315 10364 18623 10373
rect 18315 10362 18321 10364
rect 18377 10362 18401 10364
rect 18457 10362 18481 10364
rect 18537 10362 18561 10364
rect 18617 10362 18623 10364
rect 18377 10310 18379 10362
rect 18559 10310 18561 10362
rect 18315 10308 18321 10310
rect 18377 10308 18401 10310
rect 18457 10308 18481 10310
rect 18537 10308 18561 10310
rect 18617 10308 18623 10310
rect 18315 10299 18623 10308
rect 18315 9276 18623 9285
rect 18315 9274 18321 9276
rect 18377 9274 18401 9276
rect 18457 9274 18481 9276
rect 18537 9274 18561 9276
rect 18617 9274 18623 9276
rect 18377 9222 18379 9274
rect 18559 9222 18561 9274
rect 18315 9220 18321 9222
rect 18377 9220 18401 9222
rect 18457 9220 18481 9222
rect 18537 9220 18561 9222
rect 18617 9220 18623 9222
rect 18315 9211 18623 9220
rect 18315 8188 18623 8197
rect 18315 8186 18321 8188
rect 18377 8186 18401 8188
rect 18457 8186 18481 8188
rect 18537 8186 18561 8188
rect 18617 8186 18623 8188
rect 18377 8134 18379 8186
rect 18559 8134 18561 8186
rect 18315 8132 18321 8134
rect 18377 8132 18401 8134
rect 18457 8132 18481 8134
rect 18537 8132 18561 8134
rect 18617 8132 18623 8134
rect 18315 8123 18623 8132
rect 18315 7100 18623 7109
rect 18315 7098 18321 7100
rect 18377 7098 18401 7100
rect 18457 7098 18481 7100
rect 18537 7098 18561 7100
rect 18617 7098 18623 7100
rect 18377 7046 18379 7098
rect 18559 7046 18561 7098
rect 18315 7044 18321 7046
rect 18377 7044 18401 7046
rect 18457 7044 18481 7046
rect 18537 7044 18561 7046
rect 18617 7044 18623 7046
rect 18315 7035 18623 7044
rect 19628 6866 19656 11206
rect 19720 11150 19748 11494
rect 19812 11150 19840 11630
rect 21008 11218 21036 11630
rect 20996 11212 21048 11218
rect 20996 11154 21048 11160
rect 19708 11144 19760 11150
rect 19708 11086 19760 11092
rect 19800 11144 19852 11150
rect 19800 11086 19852 11092
rect 20720 11144 20772 11150
rect 20720 11086 20772 11092
rect 20732 10674 20760 11086
rect 20904 11008 20956 11014
rect 20904 10950 20956 10956
rect 20916 10674 20944 10950
rect 21100 10810 21128 12174
rect 21088 10804 21140 10810
rect 21088 10746 21140 10752
rect 20720 10668 20772 10674
rect 20720 10610 20772 10616
rect 20904 10668 20956 10674
rect 20904 10610 20956 10616
rect 21376 9586 21404 12406
rect 21548 12378 21600 12384
rect 21652 11898 21680 13942
rect 21788 13084 22096 13093
rect 21788 13082 21794 13084
rect 21850 13082 21874 13084
rect 21930 13082 21954 13084
rect 22010 13082 22034 13084
rect 22090 13082 22096 13084
rect 21850 13030 21852 13082
rect 22032 13030 22034 13082
rect 21788 13028 21794 13030
rect 21850 13028 21874 13030
rect 21930 13028 21954 13030
rect 22010 13028 22034 13030
rect 22090 13028 22096 13030
rect 21788 13019 22096 13028
rect 22296 12850 22324 17478
rect 22376 16448 22428 16454
rect 22376 16390 22428 16396
rect 22388 16250 22416 16390
rect 22376 16244 22428 16250
rect 22376 16186 22428 16192
rect 22572 16046 22600 18142
rect 23216 17678 23244 18770
rect 23388 18692 23440 18698
rect 23388 18634 23440 18640
rect 23400 17678 23428 18634
rect 23492 18426 23520 19314
rect 23664 18624 23716 18630
rect 23716 18572 23796 18578
rect 23664 18566 23796 18572
rect 23676 18550 23796 18566
rect 23480 18420 23532 18426
rect 23480 18362 23532 18368
rect 23204 17672 23256 17678
rect 23204 17614 23256 17620
rect 23388 17672 23440 17678
rect 23388 17614 23440 17620
rect 23492 17202 23520 18362
rect 23664 18080 23716 18086
rect 23664 18022 23716 18028
rect 23676 17202 23704 18022
rect 23480 17196 23532 17202
rect 23480 17138 23532 17144
rect 23664 17196 23716 17202
rect 23664 17138 23716 17144
rect 23020 16992 23072 16998
rect 23020 16934 23072 16940
rect 23032 16590 23060 16934
rect 23492 16658 23520 17138
rect 23480 16652 23532 16658
rect 23480 16594 23532 16600
rect 23020 16584 23072 16590
rect 23020 16526 23072 16532
rect 23492 16046 23520 16594
rect 23768 16590 23796 18550
rect 23848 18284 23900 18290
rect 23848 18226 23900 18232
rect 23756 16584 23808 16590
rect 23756 16526 23808 16532
rect 22560 16040 22612 16046
rect 22560 15982 22612 15988
rect 23480 16040 23532 16046
rect 23480 15982 23532 15988
rect 22376 14816 22428 14822
rect 22376 14758 22428 14764
rect 22284 12844 22336 12850
rect 22284 12786 22336 12792
rect 22296 12238 22324 12786
rect 22284 12232 22336 12238
rect 22284 12174 22336 12180
rect 22388 12102 22416 14758
rect 22572 12306 22600 15982
rect 22836 15972 22888 15978
rect 22836 15914 22888 15920
rect 22652 15360 22704 15366
rect 22652 15302 22704 15308
rect 22664 14278 22692 15302
rect 22652 14272 22704 14278
rect 22652 14214 22704 14220
rect 22560 12300 22612 12306
rect 22560 12242 22612 12248
rect 22468 12232 22520 12238
rect 22468 12174 22520 12180
rect 22192 12096 22244 12102
rect 22192 12038 22244 12044
rect 22376 12096 22428 12102
rect 22376 12038 22428 12044
rect 21788 11996 22096 12005
rect 21788 11994 21794 11996
rect 21850 11994 21874 11996
rect 21930 11994 21954 11996
rect 22010 11994 22034 11996
rect 22090 11994 22096 11996
rect 21850 11942 21852 11994
rect 22032 11942 22034 11994
rect 21788 11940 21794 11942
rect 21850 11940 21874 11942
rect 21930 11940 21954 11942
rect 22010 11940 22034 11942
rect 22090 11940 22096 11942
rect 21788 11931 22096 11940
rect 21640 11892 21692 11898
rect 21640 11834 21692 11840
rect 22204 11150 22232 12038
rect 22376 11892 22428 11898
rect 22376 11834 22428 11840
rect 22388 11354 22416 11834
rect 22376 11348 22428 11354
rect 22376 11290 22428 11296
rect 22480 11218 22508 12174
rect 22560 12096 22612 12102
rect 22560 12038 22612 12044
rect 22468 11212 22520 11218
rect 22468 11154 22520 11160
rect 22192 11144 22244 11150
rect 22192 11086 22244 11092
rect 21788 10908 22096 10917
rect 21788 10906 21794 10908
rect 21850 10906 21874 10908
rect 21930 10906 21954 10908
rect 22010 10906 22034 10908
rect 22090 10906 22096 10908
rect 21850 10854 21852 10906
rect 22032 10854 22034 10906
rect 21788 10852 21794 10854
rect 21850 10852 21874 10854
rect 21930 10852 21954 10854
rect 22010 10852 22034 10854
rect 22090 10852 22096 10854
rect 21788 10843 22096 10852
rect 22376 10736 22428 10742
rect 22376 10678 22428 10684
rect 22388 10606 22416 10678
rect 22572 10606 22600 12038
rect 22664 11082 22692 14214
rect 22744 12844 22796 12850
rect 22744 12786 22796 12792
rect 22756 12306 22784 12786
rect 22848 12434 22876 15914
rect 23112 15020 23164 15026
rect 23112 14962 23164 14968
rect 22848 12406 22968 12434
rect 22744 12300 22796 12306
rect 22744 12242 22796 12248
rect 22652 11076 22704 11082
rect 22652 11018 22704 11024
rect 22756 10810 22784 12242
rect 22940 12238 22968 12406
rect 22928 12232 22980 12238
rect 22928 12174 22980 12180
rect 23020 12096 23072 12102
rect 23020 12038 23072 12044
rect 23032 11778 23060 12038
rect 23124 11898 23152 14962
rect 23388 13728 23440 13734
rect 23388 13670 23440 13676
rect 23400 12374 23428 13670
rect 23480 12640 23532 12646
rect 23480 12582 23532 12588
rect 23388 12368 23440 12374
rect 23388 12310 23440 12316
rect 23388 12232 23440 12238
rect 23388 12174 23440 12180
rect 23296 12096 23348 12102
rect 23296 12038 23348 12044
rect 23112 11892 23164 11898
rect 23112 11834 23164 11840
rect 23204 11892 23256 11898
rect 23204 11834 23256 11840
rect 23032 11750 23152 11778
rect 23124 11558 23152 11750
rect 23216 11626 23244 11834
rect 23308 11830 23336 12038
rect 23296 11824 23348 11830
rect 23296 11766 23348 11772
rect 23204 11620 23256 11626
rect 23204 11562 23256 11568
rect 23112 11552 23164 11558
rect 23112 11494 23164 11500
rect 23124 11286 23152 11494
rect 23400 11370 23428 12174
rect 23492 11728 23520 12582
rect 23572 12436 23624 12442
rect 23572 12378 23624 12384
rect 23584 12170 23612 12378
rect 23768 12374 23796 16526
rect 23860 16522 23888 18226
rect 23940 18148 23992 18154
rect 23940 18090 23992 18096
rect 23952 17270 23980 18090
rect 23940 17264 23992 17270
rect 23940 17206 23992 17212
rect 24044 16658 24072 21286
rect 24136 17542 24164 21490
rect 24320 21486 24348 22578
rect 24400 22228 24452 22234
rect 24400 22170 24452 22176
rect 24412 21622 24440 22170
rect 24400 21616 24452 21622
rect 24400 21558 24452 21564
rect 24308 21480 24360 21486
rect 24308 21422 24360 21428
rect 24504 19922 24532 26930
rect 24492 19916 24544 19922
rect 24492 19858 24544 19864
rect 24596 18986 24624 28478
rect 24688 26858 24716 28698
rect 24768 27872 24820 27878
rect 24768 27814 24820 27820
rect 24676 26852 24728 26858
rect 24676 26794 24728 26800
rect 24676 26580 24728 26586
rect 24676 26522 24728 26528
rect 24688 24750 24716 26522
rect 24676 24744 24728 24750
rect 24676 24686 24728 24692
rect 24676 24608 24728 24614
rect 24676 24550 24728 24556
rect 24688 24206 24716 24550
rect 24676 24200 24728 24206
rect 24676 24142 24728 24148
rect 24676 23112 24728 23118
rect 24676 23054 24728 23060
rect 24688 22982 24716 23054
rect 24676 22976 24728 22982
rect 24676 22918 24728 22924
rect 24676 22024 24728 22030
rect 24676 21966 24728 21972
rect 24688 19990 24716 21966
rect 24676 19984 24728 19990
rect 24676 19926 24728 19932
rect 24688 19378 24716 19926
rect 24780 19854 24808 27814
rect 24872 25294 24900 28999
rect 24952 27464 25004 27470
rect 24952 27406 25004 27412
rect 24964 27282 24992 27406
rect 25056 27402 25084 29446
rect 25884 29102 25912 29582
rect 25976 29306 26004 30194
rect 26056 30116 26108 30122
rect 26056 30058 26108 30064
rect 26068 29646 26096 30058
rect 26160 29782 26188 30194
rect 26240 30048 26292 30054
rect 26240 29990 26292 29996
rect 26148 29776 26200 29782
rect 26148 29718 26200 29724
rect 26056 29640 26108 29646
rect 26056 29582 26108 29588
rect 25964 29300 26016 29306
rect 25964 29242 26016 29248
rect 25872 29096 25924 29102
rect 25872 29038 25924 29044
rect 26068 29034 26096 29582
rect 26056 29028 26108 29034
rect 26056 28970 26108 28976
rect 25261 28860 25569 28869
rect 25261 28858 25267 28860
rect 25323 28858 25347 28860
rect 25403 28858 25427 28860
rect 25483 28858 25507 28860
rect 25563 28858 25569 28860
rect 25323 28806 25325 28858
rect 25505 28806 25507 28858
rect 25261 28804 25267 28806
rect 25323 28804 25347 28806
rect 25403 28804 25427 28806
rect 25483 28804 25507 28806
rect 25563 28804 25569 28806
rect 25261 28795 25569 28804
rect 25136 28620 25188 28626
rect 25136 28562 25188 28568
rect 25148 28014 25176 28562
rect 25780 28076 25832 28082
rect 25780 28018 25832 28024
rect 25136 28008 25188 28014
rect 25136 27950 25188 27956
rect 25148 27606 25176 27950
rect 25596 27872 25648 27878
rect 25596 27814 25648 27820
rect 25261 27772 25569 27781
rect 25261 27770 25267 27772
rect 25323 27770 25347 27772
rect 25403 27770 25427 27772
rect 25483 27770 25507 27772
rect 25563 27770 25569 27772
rect 25323 27718 25325 27770
rect 25505 27718 25507 27770
rect 25261 27716 25267 27718
rect 25323 27716 25347 27718
rect 25403 27716 25427 27718
rect 25483 27716 25507 27718
rect 25563 27716 25569 27718
rect 25261 27707 25569 27716
rect 25136 27600 25188 27606
rect 25136 27542 25188 27548
rect 25608 27554 25636 27814
rect 25792 27674 25820 28018
rect 25780 27668 25832 27674
rect 25780 27610 25832 27616
rect 25044 27396 25096 27402
rect 25044 27338 25096 27344
rect 24964 27254 25084 27282
rect 24952 25356 25004 25362
rect 24952 25298 25004 25304
rect 24860 25288 24912 25294
rect 24860 25230 24912 25236
rect 24964 24410 24992 25298
rect 25056 25294 25084 27254
rect 25148 26382 25176 27542
rect 25608 27526 25728 27554
rect 25596 27396 25648 27402
rect 25596 27338 25648 27344
rect 25261 26684 25569 26693
rect 25261 26682 25267 26684
rect 25323 26682 25347 26684
rect 25403 26682 25427 26684
rect 25483 26682 25507 26684
rect 25563 26682 25569 26684
rect 25323 26630 25325 26682
rect 25505 26630 25507 26682
rect 25261 26628 25267 26630
rect 25323 26628 25347 26630
rect 25403 26628 25427 26630
rect 25483 26628 25507 26630
rect 25563 26628 25569 26630
rect 25261 26619 25569 26628
rect 25136 26376 25188 26382
rect 25136 26318 25188 26324
rect 25504 26240 25556 26246
rect 25504 26182 25556 26188
rect 25516 25906 25544 26182
rect 25608 26042 25636 27338
rect 25596 26036 25648 26042
rect 25596 25978 25648 25984
rect 25504 25900 25556 25906
rect 25504 25842 25556 25848
rect 25700 25702 25728 27526
rect 25964 26240 26016 26246
rect 25964 26182 26016 26188
rect 25976 25906 26004 26182
rect 26068 25974 26096 28970
rect 26252 28150 26280 29990
rect 26240 28144 26292 28150
rect 26240 28086 26292 28092
rect 26240 26308 26292 26314
rect 26240 26250 26292 26256
rect 26056 25968 26108 25974
rect 26056 25910 26108 25916
rect 25964 25900 26016 25906
rect 25964 25842 26016 25848
rect 25872 25764 25924 25770
rect 25872 25706 25924 25712
rect 25688 25696 25740 25702
rect 25688 25638 25740 25644
rect 25780 25696 25832 25702
rect 25780 25638 25832 25644
rect 25261 25596 25569 25605
rect 25261 25594 25267 25596
rect 25323 25594 25347 25596
rect 25403 25594 25427 25596
rect 25483 25594 25507 25596
rect 25563 25594 25569 25596
rect 25323 25542 25325 25594
rect 25505 25542 25507 25594
rect 25261 25540 25267 25542
rect 25323 25540 25347 25542
rect 25403 25540 25427 25542
rect 25483 25540 25507 25542
rect 25563 25540 25569 25542
rect 25261 25531 25569 25540
rect 25700 25362 25728 25638
rect 25688 25356 25740 25362
rect 25688 25298 25740 25304
rect 25044 25288 25096 25294
rect 25044 25230 25096 25236
rect 25228 25288 25280 25294
rect 25228 25230 25280 25236
rect 25596 25288 25648 25294
rect 25596 25230 25648 25236
rect 25240 24954 25268 25230
rect 25228 24948 25280 24954
rect 25228 24890 25280 24896
rect 25608 24818 25636 25230
rect 25596 24812 25648 24818
rect 25596 24754 25648 24760
rect 25261 24508 25569 24517
rect 25261 24506 25267 24508
rect 25323 24506 25347 24508
rect 25403 24506 25427 24508
rect 25483 24506 25507 24508
rect 25563 24506 25569 24508
rect 25323 24454 25325 24506
rect 25505 24454 25507 24506
rect 25261 24452 25267 24454
rect 25323 24452 25347 24454
rect 25403 24452 25427 24454
rect 25483 24452 25507 24454
rect 25563 24452 25569 24454
rect 25261 24443 25569 24452
rect 24952 24404 25004 24410
rect 24952 24346 25004 24352
rect 25700 24206 25728 25298
rect 25792 24750 25820 25638
rect 25884 24818 25912 25706
rect 25976 25294 26004 25842
rect 26148 25832 26200 25838
rect 26148 25774 26200 25780
rect 25964 25288 26016 25294
rect 25964 25230 26016 25236
rect 26160 24886 26188 25774
rect 26252 25498 26280 26250
rect 26240 25492 26292 25498
rect 26240 25434 26292 25440
rect 26148 24880 26200 24886
rect 26148 24822 26200 24828
rect 25872 24812 25924 24818
rect 25872 24754 25924 24760
rect 25780 24744 25832 24750
rect 25780 24686 25832 24692
rect 24860 24200 24912 24206
rect 24860 24142 24912 24148
rect 25688 24200 25740 24206
rect 25688 24142 25740 24148
rect 24872 21894 24900 24142
rect 25261 23420 25569 23429
rect 25261 23418 25267 23420
rect 25323 23418 25347 23420
rect 25403 23418 25427 23420
rect 25483 23418 25507 23420
rect 25563 23418 25569 23420
rect 25323 23366 25325 23418
rect 25505 23366 25507 23418
rect 25261 23364 25267 23366
rect 25323 23364 25347 23366
rect 25403 23364 25427 23366
rect 25483 23364 25507 23366
rect 25563 23364 25569 23366
rect 25261 23355 25569 23364
rect 25792 23186 25820 24686
rect 25044 23180 25096 23186
rect 25044 23122 25096 23128
rect 25780 23180 25832 23186
rect 25780 23122 25832 23128
rect 25056 22094 25084 23122
rect 26160 23050 26188 24822
rect 26148 23044 26200 23050
rect 26148 22986 26200 22992
rect 25596 22976 25648 22982
rect 25596 22918 25648 22924
rect 25228 22636 25280 22642
rect 25228 22578 25280 22584
rect 25240 22522 25268 22578
rect 25148 22494 25268 22522
rect 25148 22234 25176 22494
rect 25261 22332 25569 22341
rect 25261 22330 25267 22332
rect 25323 22330 25347 22332
rect 25403 22330 25427 22332
rect 25483 22330 25507 22332
rect 25563 22330 25569 22332
rect 25323 22278 25325 22330
rect 25505 22278 25507 22330
rect 25261 22276 25267 22278
rect 25323 22276 25347 22278
rect 25403 22276 25427 22278
rect 25483 22276 25507 22278
rect 25563 22276 25569 22278
rect 25261 22267 25569 22276
rect 25136 22228 25188 22234
rect 25136 22170 25188 22176
rect 25056 22066 25360 22094
rect 24860 21888 24912 21894
rect 24860 21830 24912 21836
rect 24872 21554 24900 21830
rect 25332 21554 25360 22066
rect 25608 21622 25636 22918
rect 26160 22778 26188 22986
rect 26148 22772 26200 22778
rect 26148 22714 26200 22720
rect 26160 22030 26188 22714
rect 26148 22024 26200 22030
rect 26148 21966 26200 21972
rect 25596 21616 25648 21622
rect 25596 21558 25648 21564
rect 24860 21548 24912 21554
rect 24860 21490 24912 21496
rect 25044 21548 25096 21554
rect 25044 21490 25096 21496
rect 25320 21548 25372 21554
rect 25320 21490 25372 21496
rect 25688 21548 25740 21554
rect 25688 21490 25740 21496
rect 25056 19854 25084 21490
rect 25332 21418 25360 21490
rect 25320 21412 25372 21418
rect 25320 21354 25372 21360
rect 25136 21344 25188 21350
rect 25136 21286 25188 21292
rect 24768 19848 24820 19854
rect 24768 19790 24820 19796
rect 25044 19848 25096 19854
rect 25044 19790 25096 19796
rect 24860 19712 24912 19718
rect 24860 19654 24912 19660
rect 24676 19372 24728 19378
rect 24676 19314 24728 19320
rect 24504 18958 24624 18986
rect 24124 17536 24176 17542
rect 24124 17478 24176 17484
rect 24032 16652 24084 16658
rect 24032 16594 24084 16600
rect 23848 16516 23900 16522
rect 23848 16458 23900 16464
rect 23860 16130 23888 16458
rect 23860 16102 23980 16130
rect 23848 16040 23900 16046
rect 23848 15982 23900 15988
rect 23860 15026 23888 15982
rect 23848 15020 23900 15026
rect 23848 14962 23900 14968
rect 23860 14482 23888 14962
rect 23848 14476 23900 14482
rect 23848 14418 23900 14424
rect 23952 14362 23980 16102
rect 23860 14334 23980 14362
rect 23860 12646 23888 14334
rect 23848 12640 23900 12646
rect 23848 12582 23900 12588
rect 23756 12368 23808 12374
rect 23756 12310 23808 12316
rect 23664 12232 23716 12238
rect 23664 12174 23716 12180
rect 23572 12164 23624 12170
rect 23572 12106 23624 12112
rect 23572 11756 23624 11762
rect 23480 11722 23532 11728
rect 23572 11698 23624 11704
rect 23480 11664 23532 11670
rect 23308 11354 23428 11370
rect 23584 11354 23612 11698
rect 23308 11348 23440 11354
rect 23308 11342 23388 11348
rect 23112 11280 23164 11286
rect 23112 11222 23164 11228
rect 22744 10804 22796 10810
rect 22744 10746 22796 10752
rect 22376 10600 22428 10606
rect 22376 10542 22428 10548
rect 22560 10600 22612 10606
rect 22560 10542 22612 10548
rect 23124 10470 23152 11222
rect 23308 11014 23336 11342
rect 23388 11290 23440 11296
rect 23572 11348 23624 11354
rect 23572 11290 23624 11296
rect 23388 11212 23440 11218
rect 23388 11154 23440 11160
rect 23296 11008 23348 11014
rect 23296 10950 23348 10956
rect 23308 10742 23336 10950
rect 23296 10736 23348 10742
rect 23296 10678 23348 10684
rect 23400 10606 23428 11154
rect 23676 11082 23704 12174
rect 23860 11830 23888 12582
rect 24044 12306 24072 16594
rect 24504 16182 24532 18958
rect 24584 18828 24636 18834
rect 24584 18770 24636 18776
rect 24596 18426 24624 18770
rect 24584 18420 24636 18426
rect 24584 18362 24636 18368
rect 24596 17746 24624 18362
rect 24584 17740 24636 17746
rect 24584 17682 24636 17688
rect 24688 17338 24716 19314
rect 24872 17678 24900 19654
rect 25056 19446 25084 19790
rect 25044 19440 25096 19446
rect 25044 19382 25096 19388
rect 25148 19378 25176 21286
rect 25261 21244 25569 21253
rect 25261 21242 25267 21244
rect 25323 21242 25347 21244
rect 25403 21242 25427 21244
rect 25483 21242 25507 21244
rect 25563 21242 25569 21244
rect 25323 21190 25325 21242
rect 25505 21190 25507 21242
rect 25261 21188 25267 21190
rect 25323 21188 25347 21190
rect 25403 21188 25427 21190
rect 25483 21188 25507 21190
rect 25563 21188 25569 21190
rect 25261 21179 25569 21188
rect 25700 20602 25728 21490
rect 25688 20596 25740 20602
rect 25688 20538 25740 20544
rect 25596 20528 25648 20534
rect 25596 20470 25648 20476
rect 25261 20156 25569 20165
rect 25261 20154 25267 20156
rect 25323 20154 25347 20156
rect 25403 20154 25427 20156
rect 25483 20154 25507 20156
rect 25563 20154 25569 20156
rect 25323 20102 25325 20154
rect 25505 20102 25507 20154
rect 25261 20100 25267 20102
rect 25323 20100 25347 20102
rect 25403 20100 25427 20102
rect 25483 20100 25507 20102
rect 25563 20100 25569 20102
rect 25261 20091 25569 20100
rect 25228 19848 25280 19854
rect 25228 19790 25280 19796
rect 25136 19372 25188 19378
rect 25136 19314 25188 19320
rect 25240 19258 25268 19790
rect 25608 19514 25636 20470
rect 25596 19508 25648 19514
rect 25596 19450 25648 19456
rect 25700 19378 25728 20538
rect 26146 19816 26202 19825
rect 26146 19751 26202 19760
rect 25688 19372 25740 19378
rect 25688 19314 25740 19320
rect 25056 19230 25268 19258
rect 24952 18760 25004 18766
rect 24952 18702 25004 18708
rect 24860 17672 24912 17678
rect 24860 17614 24912 17620
rect 24676 17332 24728 17338
rect 24676 17274 24728 17280
rect 24688 16454 24716 17274
rect 24964 16998 24992 18702
rect 25056 17542 25084 19230
rect 25261 19068 25569 19077
rect 25261 19066 25267 19068
rect 25323 19066 25347 19068
rect 25403 19066 25427 19068
rect 25483 19066 25507 19068
rect 25563 19066 25569 19068
rect 25323 19014 25325 19066
rect 25505 19014 25507 19066
rect 25261 19012 25267 19014
rect 25323 19012 25347 19014
rect 25403 19012 25427 19014
rect 25483 19012 25507 19014
rect 25563 19012 25569 19014
rect 25261 19003 25569 19012
rect 25261 17980 25569 17989
rect 25261 17978 25267 17980
rect 25323 17978 25347 17980
rect 25403 17978 25427 17980
rect 25483 17978 25507 17980
rect 25563 17978 25569 17980
rect 25323 17926 25325 17978
rect 25505 17926 25507 17978
rect 25261 17924 25267 17926
rect 25323 17924 25347 17926
rect 25403 17924 25427 17926
rect 25483 17924 25507 17926
rect 25563 17924 25569 17926
rect 25261 17915 25569 17924
rect 26160 17746 26188 19751
rect 26148 17740 26200 17746
rect 26148 17682 26200 17688
rect 25044 17536 25096 17542
rect 25044 17478 25096 17484
rect 24952 16992 25004 16998
rect 24952 16934 25004 16940
rect 24676 16448 24728 16454
rect 24676 16390 24728 16396
rect 24860 16448 24912 16454
rect 24860 16390 24912 16396
rect 24492 16176 24544 16182
rect 24492 16118 24544 16124
rect 24216 14476 24268 14482
rect 24216 14418 24268 14424
rect 24228 13938 24256 14418
rect 24584 14340 24636 14346
rect 24584 14282 24636 14288
rect 24216 13932 24268 13938
rect 24216 13874 24268 13880
rect 24308 12844 24360 12850
rect 24308 12786 24360 12792
rect 24492 12844 24544 12850
rect 24492 12786 24544 12792
rect 24216 12776 24268 12782
rect 24216 12718 24268 12724
rect 24032 12300 24084 12306
rect 24032 12242 24084 12248
rect 24044 11830 24072 12242
rect 24228 12170 24256 12718
rect 24216 12164 24268 12170
rect 24216 12106 24268 12112
rect 23848 11824 23900 11830
rect 23848 11766 23900 11772
rect 24032 11824 24084 11830
rect 24032 11766 24084 11772
rect 24228 11762 24256 12106
rect 24320 11898 24348 12786
rect 24504 12646 24532 12786
rect 24492 12640 24544 12646
rect 24492 12582 24544 12588
rect 24400 12368 24452 12374
rect 24400 12310 24452 12316
rect 24308 11892 24360 11898
rect 24308 11834 24360 11840
rect 24216 11756 24268 11762
rect 24216 11698 24268 11704
rect 24412 11694 24440 12310
rect 24504 12306 24532 12582
rect 24596 12442 24624 14282
rect 24688 12918 24716 16390
rect 24872 16114 24900 16390
rect 24860 16108 24912 16114
rect 24860 16050 24912 16056
rect 24768 13932 24820 13938
rect 24768 13874 24820 13880
rect 24780 12986 24808 13874
rect 24768 12980 24820 12986
rect 24768 12922 24820 12928
rect 24676 12912 24728 12918
rect 24676 12854 24728 12860
rect 24584 12436 24636 12442
rect 24584 12378 24636 12384
rect 24492 12300 24544 12306
rect 24492 12242 24544 12248
rect 24860 12232 24912 12238
rect 24860 12174 24912 12180
rect 24872 11898 24900 12174
rect 24860 11892 24912 11898
rect 24860 11834 24912 11840
rect 24860 11756 24912 11762
rect 24860 11698 24912 11704
rect 24400 11688 24452 11694
rect 24400 11630 24452 11636
rect 24412 11150 24440 11630
rect 24768 11620 24820 11626
rect 24768 11562 24820 11568
rect 24400 11144 24452 11150
rect 24400 11086 24452 11092
rect 24780 11098 24808 11562
rect 24872 11286 24900 11698
rect 24964 11286 24992 16934
rect 24860 11280 24912 11286
rect 24860 11222 24912 11228
rect 24952 11280 25004 11286
rect 24952 11222 25004 11228
rect 24952 11144 25004 11150
rect 24780 11092 24952 11098
rect 24780 11086 25004 11092
rect 23664 11076 23716 11082
rect 24780 11070 24992 11086
rect 23664 11018 23716 11024
rect 23388 10600 23440 10606
rect 23388 10542 23440 10548
rect 23112 10464 23164 10470
rect 23112 10406 23164 10412
rect 21788 9820 22096 9829
rect 21788 9818 21794 9820
rect 21850 9818 21874 9820
rect 21930 9818 21954 9820
rect 22010 9818 22034 9820
rect 22090 9818 22096 9820
rect 21850 9766 21852 9818
rect 22032 9766 22034 9818
rect 21788 9764 21794 9766
rect 21850 9764 21874 9766
rect 21930 9764 21954 9766
rect 22010 9764 22034 9766
rect 22090 9764 22096 9766
rect 21788 9755 22096 9764
rect 21364 9580 21416 9586
rect 21364 9522 21416 9528
rect 21788 8732 22096 8741
rect 21788 8730 21794 8732
rect 21850 8730 21874 8732
rect 21930 8730 21954 8732
rect 22010 8730 22034 8732
rect 22090 8730 22096 8732
rect 21850 8678 21852 8730
rect 22032 8678 22034 8730
rect 21788 8676 21794 8678
rect 21850 8676 21874 8678
rect 21930 8676 21954 8678
rect 22010 8676 22034 8678
rect 22090 8676 22096 8678
rect 21788 8667 22096 8676
rect 21788 7644 22096 7653
rect 21788 7642 21794 7644
rect 21850 7642 21874 7644
rect 21930 7642 21954 7644
rect 22010 7642 22034 7644
rect 22090 7642 22096 7644
rect 21850 7590 21852 7642
rect 22032 7590 22034 7642
rect 21788 7588 21794 7590
rect 21850 7588 21874 7590
rect 21930 7588 21954 7590
rect 22010 7588 22034 7590
rect 22090 7588 22096 7590
rect 21788 7579 22096 7588
rect 19616 6860 19668 6866
rect 19616 6802 19668 6808
rect 23848 6656 23900 6662
rect 23848 6598 23900 6604
rect 21788 6556 22096 6565
rect 21788 6554 21794 6556
rect 21850 6554 21874 6556
rect 21930 6554 21954 6556
rect 22010 6554 22034 6556
rect 22090 6554 22096 6556
rect 21850 6502 21852 6554
rect 22032 6502 22034 6554
rect 21788 6500 21794 6502
rect 21850 6500 21874 6502
rect 21930 6500 21954 6502
rect 22010 6500 22034 6502
rect 22090 6500 22096 6502
rect 21788 6491 22096 6500
rect 18315 6012 18623 6021
rect 18315 6010 18321 6012
rect 18377 6010 18401 6012
rect 18457 6010 18481 6012
rect 18537 6010 18561 6012
rect 18617 6010 18623 6012
rect 18377 5958 18379 6010
rect 18559 5958 18561 6010
rect 18315 5956 18321 5958
rect 18377 5956 18401 5958
rect 18457 5956 18481 5958
rect 18537 5956 18561 5958
rect 18617 5956 18623 5958
rect 18315 5947 18623 5956
rect 21788 5468 22096 5477
rect 21788 5466 21794 5468
rect 21850 5466 21874 5468
rect 21930 5466 21954 5468
rect 22010 5466 22034 5468
rect 22090 5466 22096 5468
rect 21850 5414 21852 5466
rect 22032 5414 22034 5466
rect 21788 5412 21794 5414
rect 21850 5412 21874 5414
rect 21930 5412 21954 5414
rect 22010 5412 22034 5414
rect 22090 5412 22096 5414
rect 21788 5403 22096 5412
rect 18315 4924 18623 4933
rect 18315 4922 18321 4924
rect 18377 4922 18401 4924
rect 18457 4922 18481 4924
rect 18537 4922 18561 4924
rect 18617 4922 18623 4924
rect 18377 4870 18379 4922
rect 18559 4870 18561 4922
rect 18315 4868 18321 4870
rect 18377 4868 18401 4870
rect 18457 4868 18481 4870
rect 18537 4868 18561 4870
rect 18617 4868 18623 4870
rect 18315 4859 18623 4868
rect 22192 4548 22244 4554
rect 22192 4490 22244 4496
rect 23756 4548 23808 4554
rect 23756 4490 23808 4496
rect 21788 4380 22096 4389
rect 21788 4378 21794 4380
rect 21850 4378 21874 4380
rect 21930 4378 21954 4380
rect 22010 4378 22034 4380
rect 22090 4378 22096 4380
rect 21850 4326 21852 4378
rect 22032 4326 22034 4378
rect 21788 4324 21794 4326
rect 21850 4324 21874 4326
rect 21930 4324 21954 4326
rect 22010 4324 22034 4326
rect 22090 4324 22096 4326
rect 21788 4315 22096 4324
rect 21180 4140 21232 4146
rect 21180 4082 21232 4088
rect 22100 4140 22152 4146
rect 22100 4082 22152 4088
rect 18144 4004 18196 4010
rect 18144 3946 18196 3952
rect 18156 3534 18184 3946
rect 19616 3936 19668 3942
rect 19616 3878 19668 3884
rect 20352 3936 20404 3942
rect 20352 3878 20404 3884
rect 20536 3936 20588 3942
rect 20536 3878 20588 3884
rect 18315 3836 18623 3845
rect 18315 3834 18321 3836
rect 18377 3834 18401 3836
rect 18457 3834 18481 3836
rect 18537 3834 18561 3836
rect 18617 3834 18623 3836
rect 18377 3782 18379 3834
rect 18559 3782 18561 3834
rect 18315 3780 18321 3782
rect 18377 3780 18401 3782
rect 18457 3780 18481 3782
rect 18537 3780 18561 3782
rect 18617 3780 18623 3782
rect 18315 3771 18623 3780
rect 18144 3528 18196 3534
rect 18144 3470 18196 3476
rect 19432 3528 19484 3534
rect 19432 3470 19484 3476
rect 19156 3460 19208 3466
rect 19156 3402 19208 3408
rect 19168 3058 19196 3402
rect 19340 3392 19392 3398
rect 19340 3334 19392 3340
rect 19352 3126 19380 3334
rect 19340 3120 19392 3126
rect 19340 3062 19392 3068
rect 19156 3052 19208 3058
rect 19156 2994 19208 3000
rect 18052 2916 18104 2922
rect 18052 2858 18104 2864
rect 17592 2644 17644 2650
rect 17592 2586 17644 2592
rect 17408 2440 17460 2446
rect 17408 2382 17460 2388
rect 17420 800 17448 2382
rect 18064 800 18092 2858
rect 18315 2748 18623 2757
rect 18315 2746 18321 2748
rect 18377 2746 18401 2748
rect 18457 2746 18481 2748
rect 18537 2746 18561 2748
rect 18617 2746 18623 2748
rect 18377 2694 18379 2746
rect 18559 2694 18561 2746
rect 18315 2692 18321 2694
rect 18377 2692 18401 2694
rect 18457 2692 18481 2694
rect 18537 2692 18561 2694
rect 18617 2692 18623 2694
rect 18315 2683 18623 2692
rect 19444 2514 19472 3470
rect 19628 2514 19656 3878
rect 20364 3602 20392 3878
rect 20548 3602 20576 3878
rect 21192 3670 21220 4082
rect 21180 3664 21232 3670
rect 21180 3606 21232 3612
rect 20352 3596 20404 3602
rect 20352 3538 20404 3544
rect 20536 3596 20588 3602
rect 20536 3538 20588 3544
rect 21272 3596 21324 3602
rect 21272 3538 21324 3544
rect 19432 2508 19484 2514
rect 19432 2450 19484 2456
rect 19616 2508 19668 2514
rect 19616 2450 19668 2456
rect 19984 2508 20036 2514
rect 19984 2450 20036 2456
rect 19996 800 20024 2450
rect 21284 800 21312 3538
rect 22112 3466 22140 4082
rect 22100 3460 22152 3466
rect 22100 3402 22152 3408
rect 21788 3292 22096 3301
rect 21788 3290 21794 3292
rect 21850 3290 21874 3292
rect 21930 3290 21954 3292
rect 22010 3290 22034 3292
rect 22090 3290 22096 3292
rect 21850 3238 21852 3290
rect 22032 3238 22034 3290
rect 21788 3236 21794 3238
rect 21850 3236 21874 3238
rect 21930 3236 21954 3238
rect 22010 3236 22034 3238
rect 22090 3236 22096 3238
rect 21788 3227 22096 3236
rect 21788 2204 22096 2213
rect 21788 2202 21794 2204
rect 21850 2202 21874 2204
rect 21930 2202 21954 2204
rect 22010 2202 22034 2204
rect 22090 2202 22096 2204
rect 21850 2150 21852 2202
rect 22032 2150 22034 2202
rect 21788 2148 21794 2150
rect 21850 2148 21874 2150
rect 21930 2148 21954 2150
rect 22010 2148 22034 2150
rect 22090 2148 22096 2150
rect 21788 2139 22096 2148
rect 22204 1986 22232 4490
rect 23768 4146 23796 4490
rect 23756 4140 23808 4146
rect 23756 4082 23808 4088
rect 23860 3466 23888 6598
rect 24952 5704 25004 5710
rect 24952 5646 25004 5652
rect 24964 4078 24992 5646
rect 25056 4690 25084 17478
rect 25872 17060 25924 17066
rect 25872 17002 25924 17008
rect 25261 16892 25569 16901
rect 25261 16890 25267 16892
rect 25323 16890 25347 16892
rect 25403 16890 25427 16892
rect 25483 16890 25507 16892
rect 25563 16890 25569 16892
rect 25323 16838 25325 16890
rect 25505 16838 25507 16890
rect 25261 16836 25267 16838
rect 25323 16836 25347 16838
rect 25403 16836 25427 16838
rect 25483 16836 25507 16838
rect 25563 16836 25569 16838
rect 25261 16827 25569 16836
rect 25884 16794 25912 17002
rect 25872 16788 25924 16794
rect 25872 16730 25924 16736
rect 25596 16584 25648 16590
rect 25596 16526 25648 16532
rect 25261 15804 25569 15813
rect 25261 15802 25267 15804
rect 25323 15802 25347 15804
rect 25403 15802 25427 15804
rect 25483 15802 25507 15804
rect 25563 15802 25569 15804
rect 25323 15750 25325 15802
rect 25505 15750 25507 15802
rect 25261 15748 25267 15750
rect 25323 15748 25347 15750
rect 25403 15748 25427 15750
rect 25483 15748 25507 15750
rect 25563 15748 25569 15750
rect 25261 15739 25569 15748
rect 25608 15706 25636 16526
rect 25596 15700 25648 15706
rect 25596 15642 25648 15648
rect 25884 15570 25912 16730
rect 25872 15564 25924 15570
rect 25872 15506 25924 15512
rect 25872 15360 25924 15366
rect 25872 15302 25924 15308
rect 25261 14716 25569 14725
rect 25261 14714 25267 14716
rect 25323 14714 25347 14716
rect 25403 14714 25427 14716
rect 25483 14714 25507 14716
rect 25563 14714 25569 14716
rect 25323 14662 25325 14714
rect 25505 14662 25507 14714
rect 25261 14660 25267 14662
rect 25323 14660 25347 14662
rect 25403 14660 25427 14662
rect 25483 14660 25507 14662
rect 25563 14660 25569 14662
rect 25261 14651 25569 14660
rect 25596 13728 25648 13734
rect 25596 13670 25648 13676
rect 25261 13628 25569 13637
rect 25261 13626 25267 13628
rect 25323 13626 25347 13628
rect 25403 13626 25427 13628
rect 25483 13626 25507 13628
rect 25563 13626 25569 13628
rect 25323 13574 25325 13626
rect 25505 13574 25507 13626
rect 25261 13572 25267 13574
rect 25323 13572 25347 13574
rect 25403 13572 25427 13574
rect 25483 13572 25507 13574
rect 25563 13572 25569 13574
rect 25261 13563 25569 13572
rect 25261 12540 25569 12549
rect 25261 12538 25267 12540
rect 25323 12538 25347 12540
rect 25403 12538 25427 12540
rect 25483 12538 25507 12540
rect 25563 12538 25569 12540
rect 25323 12486 25325 12538
rect 25505 12486 25507 12538
rect 25261 12484 25267 12486
rect 25323 12484 25347 12486
rect 25403 12484 25427 12486
rect 25483 12484 25507 12486
rect 25563 12484 25569 12486
rect 25261 12475 25569 12484
rect 25608 12238 25636 13670
rect 25688 12776 25740 12782
rect 25688 12718 25740 12724
rect 25700 12442 25728 12718
rect 25688 12436 25740 12442
rect 25688 12378 25740 12384
rect 25136 12232 25188 12238
rect 25136 12174 25188 12180
rect 25596 12232 25648 12238
rect 25596 12174 25648 12180
rect 25148 11354 25176 12174
rect 25608 11694 25636 12174
rect 25596 11688 25648 11694
rect 25596 11630 25648 11636
rect 25261 11452 25569 11461
rect 25261 11450 25267 11452
rect 25323 11450 25347 11452
rect 25403 11450 25427 11452
rect 25483 11450 25507 11452
rect 25563 11450 25569 11452
rect 25323 11398 25325 11450
rect 25505 11398 25507 11450
rect 25261 11396 25267 11398
rect 25323 11396 25347 11398
rect 25403 11396 25427 11398
rect 25483 11396 25507 11398
rect 25563 11396 25569 11398
rect 25261 11387 25569 11396
rect 25136 11348 25188 11354
rect 25136 11290 25188 11296
rect 25596 11212 25648 11218
rect 25596 11154 25648 11160
rect 25261 10364 25569 10373
rect 25261 10362 25267 10364
rect 25323 10362 25347 10364
rect 25403 10362 25427 10364
rect 25483 10362 25507 10364
rect 25563 10362 25569 10364
rect 25323 10310 25325 10362
rect 25505 10310 25507 10362
rect 25261 10308 25267 10310
rect 25323 10308 25347 10310
rect 25403 10308 25427 10310
rect 25483 10308 25507 10310
rect 25563 10308 25569 10310
rect 25261 10299 25569 10308
rect 25261 9276 25569 9285
rect 25261 9274 25267 9276
rect 25323 9274 25347 9276
rect 25403 9274 25427 9276
rect 25483 9274 25507 9276
rect 25563 9274 25569 9276
rect 25323 9222 25325 9274
rect 25505 9222 25507 9274
rect 25261 9220 25267 9222
rect 25323 9220 25347 9222
rect 25403 9220 25427 9222
rect 25483 9220 25507 9222
rect 25563 9220 25569 9222
rect 25261 9211 25569 9220
rect 25608 9042 25636 11154
rect 25688 9648 25740 9654
rect 25688 9590 25740 9596
rect 25596 9036 25648 9042
rect 25596 8978 25648 8984
rect 25261 8188 25569 8197
rect 25261 8186 25267 8188
rect 25323 8186 25347 8188
rect 25403 8186 25427 8188
rect 25483 8186 25507 8188
rect 25563 8186 25569 8188
rect 25323 8134 25325 8186
rect 25505 8134 25507 8186
rect 25261 8132 25267 8134
rect 25323 8132 25347 8134
rect 25403 8132 25427 8134
rect 25483 8132 25507 8134
rect 25563 8132 25569 8134
rect 25261 8123 25569 8132
rect 25261 7100 25569 7109
rect 25261 7098 25267 7100
rect 25323 7098 25347 7100
rect 25403 7098 25427 7100
rect 25483 7098 25507 7100
rect 25563 7098 25569 7100
rect 25323 7046 25325 7098
rect 25505 7046 25507 7098
rect 25261 7044 25267 7046
rect 25323 7044 25347 7046
rect 25403 7044 25427 7046
rect 25483 7044 25507 7046
rect 25563 7044 25569 7046
rect 25261 7035 25569 7044
rect 25136 6860 25188 6866
rect 25136 6802 25188 6808
rect 25044 4684 25096 4690
rect 25044 4626 25096 4632
rect 24952 4072 25004 4078
rect 24952 4014 25004 4020
rect 23848 3460 23900 3466
rect 23848 3402 23900 3408
rect 21928 1958 22232 1986
rect 21928 800 21956 1958
rect 25148 800 25176 6802
rect 25261 6012 25569 6021
rect 25261 6010 25267 6012
rect 25323 6010 25347 6012
rect 25403 6010 25427 6012
rect 25483 6010 25507 6012
rect 25563 6010 25569 6012
rect 25323 5958 25325 6010
rect 25505 5958 25507 6010
rect 25261 5956 25267 5958
rect 25323 5956 25347 5958
rect 25403 5956 25427 5958
rect 25483 5956 25507 5958
rect 25563 5956 25569 5958
rect 25261 5947 25569 5956
rect 25700 5846 25728 9590
rect 25780 9376 25832 9382
rect 25780 9318 25832 9324
rect 25792 9042 25820 9318
rect 25780 9036 25832 9042
rect 25780 8978 25832 8984
rect 25688 5840 25740 5846
rect 25688 5782 25740 5788
rect 25261 4924 25569 4933
rect 25261 4922 25267 4924
rect 25323 4922 25347 4924
rect 25403 4922 25427 4924
rect 25483 4922 25507 4924
rect 25563 4922 25569 4924
rect 25323 4870 25325 4922
rect 25505 4870 25507 4922
rect 25261 4868 25267 4870
rect 25323 4868 25347 4870
rect 25403 4868 25427 4870
rect 25483 4868 25507 4870
rect 25563 4868 25569 4870
rect 25261 4859 25569 4868
rect 25261 3836 25569 3845
rect 25261 3834 25267 3836
rect 25323 3834 25347 3836
rect 25403 3834 25427 3836
rect 25483 3834 25507 3836
rect 25563 3834 25569 3836
rect 25323 3782 25325 3834
rect 25505 3782 25507 3834
rect 25261 3780 25267 3782
rect 25323 3780 25347 3782
rect 25403 3780 25427 3782
rect 25483 3780 25507 3782
rect 25563 3780 25569 3782
rect 25261 3771 25569 3780
rect 25261 2748 25569 2757
rect 25261 2746 25267 2748
rect 25323 2746 25347 2748
rect 25403 2746 25427 2748
rect 25483 2746 25507 2748
rect 25563 2746 25569 2748
rect 25323 2694 25325 2746
rect 25505 2694 25507 2746
rect 25261 2692 25267 2694
rect 25323 2692 25347 2694
rect 25403 2692 25427 2694
rect 25483 2692 25507 2694
rect 25563 2692 25569 2694
rect 25261 2683 25569 2692
rect 25884 2650 25912 15302
rect 26344 14618 26372 30670
rect 26608 30660 26660 30666
rect 26608 30602 26660 30608
rect 26620 30394 26648 30602
rect 26608 30388 26660 30394
rect 26608 30330 26660 30336
rect 26516 30184 26568 30190
rect 26516 30126 26568 30132
rect 26528 29850 26556 30126
rect 26516 29844 26568 29850
rect 26516 29786 26568 29792
rect 26528 29646 26556 29786
rect 26516 29640 26568 29646
rect 26516 29582 26568 29588
rect 26528 29186 26556 29582
rect 26528 29170 26648 29186
rect 26528 29164 26660 29170
rect 26528 29158 26608 29164
rect 26608 29106 26660 29112
rect 26516 29028 26568 29034
rect 26516 28970 26568 28976
rect 26528 28626 26556 28970
rect 26516 28620 26568 28626
rect 26516 28562 26568 28568
rect 26620 27878 26648 29106
rect 26608 27872 26660 27878
rect 26608 27814 26660 27820
rect 26620 27674 26648 27814
rect 26608 27668 26660 27674
rect 26608 27610 26660 27616
rect 26700 25220 26752 25226
rect 26700 25162 26752 25168
rect 26712 24954 26740 25162
rect 26700 24948 26752 24954
rect 26700 24890 26752 24896
rect 26896 24818 26924 35702
rect 27068 32020 27120 32026
rect 27068 31962 27120 31968
rect 27080 30274 27108 31962
rect 27172 31754 27200 35866
rect 27252 35692 27304 35698
rect 27252 35634 27304 35640
rect 27264 33658 27292 35634
rect 27526 34096 27582 34105
rect 27526 34031 27528 34040
rect 27580 34031 27582 34040
rect 27528 34002 27580 34008
rect 27252 33652 27304 33658
rect 27252 33594 27304 33600
rect 27526 33008 27582 33017
rect 27526 32943 27528 32952
rect 27580 32943 27582 32952
rect 27528 32914 27580 32920
rect 27528 31884 27580 31890
rect 27528 31826 27580 31832
rect 27172 31726 27292 31754
rect 27080 30258 27200 30274
rect 26976 30252 27028 30258
rect 27080 30252 27212 30258
rect 27080 30246 27160 30252
rect 26976 30194 27028 30200
rect 27160 30194 27212 30200
rect 26988 25906 27016 30194
rect 27068 29504 27120 29510
rect 27068 29446 27120 29452
rect 27080 29170 27108 29446
rect 27068 29164 27120 29170
rect 27068 29106 27120 29112
rect 27080 26042 27108 29106
rect 27068 26036 27120 26042
rect 27068 25978 27120 25984
rect 26976 25900 27028 25906
rect 26976 25842 27028 25848
rect 26884 24812 26936 24818
rect 26884 24754 26936 24760
rect 26516 24200 26568 24206
rect 26516 24142 26568 24148
rect 26528 23798 26556 24142
rect 26516 23792 26568 23798
rect 26516 23734 26568 23740
rect 26884 23724 26936 23730
rect 26884 23666 26936 23672
rect 26516 23520 26568 23526
rect 26516 23462 26568 23468
rect 26528 23186 26556 23462
rect 26516 23180 26568 23186
rect 26516 23122 26568 23128
rect 26700 21344 26752 21350
rect 26700 21286 26752 21292
rect 26712 19786 26740 21286
rect 26700 19780 26752 19786
rect 26700 19722 26752 19728
rect 26516 18216 26568 18222
rect 26516 18158 26568 18164
rect 26424 17196 26476 17202
rect 26424 17138 26476 17144
rect 26436 16794 26464 17138
rect 26528 16998 26556 18158
rect 26516 16992 26568 16998
rect 26516 16934 26568 16940
rect 26424 16788 26476 16794
rect 26424 16730 26476 16736
rect 26528 16658 26556 16934
rect 26516 16652 26568 16658
rect 26516 16594 26568 16600
rect 26608 15904 26660 15910
rect 26608 15846 26660 15852
rect 26620 15502 26648 15846
rect 26608 15496 26660 15502
rect 26608 15438 26660 15444
rect 26896 15026 26924 23666
rect 26988 21486 27016 25842
rect 27068 24812 27120 24818
rect 27068 24754 27120 24760
rect 26976 21480 27028 21486
rect 26976 21422 27028 21428
rect 26884 15020 26936 15026
rect 26884 14962 26936 14968
rect 26700 14816 26752 14822
rect 26700 14758 26752 14764
rect 26332 14612 26384 14618
rect 26332 14554 26384 14560
rect 26712 14482 26740 14758
rect 26700 14476 26752 14482
rect 26700 14418 26752 14424
rect 25964 14272 26016 14278
rect 25964 14214 26016 14220
rect 25976 12238 26004 14214
rect 26700 13728 26752 13734
rect 26700 13670 26752 13676
rect 26712 13394 26740 13670
rect 26700 13388 26752 13394
rect 26700 13330 26752 13336
rect 26516 12708 26568 12714
rect 26516 12650 26568 12656
rect 26528 12306 26556 12650
rect 26700 12640 26752 12646
rect 26700 12582 26752 12588
rect 26712 12306 26740 12582
rect 26516 12300 26568 12306
rect 26516 12242 26568 12248
rect 26700 12300 26752 12306
rect 26700 12242 26752 12248
rect 25964 12232 26016 12238
rect 25964 12174 26016 12180
rect 25976 11762 26004 12174
rect 25964 11756 26016 11762
rect 25964 11698 26016 11704
rect 26700 10464 26752 10470
rect 26700 10406 26752 10412
rect 26712 10130 26740 10406
rect 26700 10124 26752 10130
rect 26700 10066 26752 10072
rect 26608 8288 26660 8294
rect 26146 8256 26202 8265
rect 26608 8230 26660 8236
rect 26146 8191 26202 8200
rect 26160 7342 26188 8191
rect 26620 7410 26648 8230
rect 26608 7404 26660 7410
rect 26608 7346 26660 7352
rect 26148 7336 26200 7342
rect 26148 7278 26200 7284
rect 26146 6896 26202 6905
rect 26146 6831 26202 6840
rect 26160 6254 26188 6831
rect 26608 6792 26660 6798
rect 26608 6734 26660 6740
rect 26620 6322 26648 6734
rect 26608 6316 26660 6322
rect 26608 6258 26660 6264
rect 26148 6248 26200 6254
rect 26148 6190 26200 6196
rect 26240 5704 26292 5710
rect 26240 5646 26292 5652
rect 26424 5704 26476 5710
rect 26424 5646 26476 5652
rect 26252 5302 26280 5646
rect 26240 5296 26292 5302
rect 26240 5238 26292 5244
rect 26436 5234 26464 5646
rect 26608 5636 26660 5642
rect 26608 5578 26660 5584
rect 26620 5370 26648 5578
rect 26608 5364 26660 5370
rect 26608 5306 26660 5312
rect 27080 5302 27108 24754
rect 27172 16114 27200 30194
rect 27264 28082 27292 31726
rect 27540 31385 27568 31826
rect 27526 31376 27582 31385
rect 27632 31346 27660 35866
rect 27712 34944 27764 34950
rect 27712 34886 27764 34892
rect 27724 34610 27752 34886
rect 27712 34604 27764 34610
rect 27712 34546 27764 34552
rect 27804 34536 27856 34542
rect 27804 34478 27856 34484
rect 27816 31754 27844 34478
rect 27908 31822 27936 35866
rect 27988 35488 28040 35494
rect 27988 35430 28040 35436
rect 28000 34066 28028 35430
rect 28080 35284 28132 35290
rect 28080 35226 28132 35232
rect 28092 34542 28120 35226
rect 28184 35018 28212 37062
rect 28368 36825 28396 37198
rect 28354 36816 28410 36825
rect 28354 36751 28410 36760
rect 28356 36168 28408 36174
rect 28354 36136 28356 36145
rect 28408 36136 28410 36145
rect 28354 36071 28410 36080
rect 28448 35692 28500 35698
rect 28448 35634 28500 35640
rect 28172 35012 28224 35018
rect 28172 34954 28224 34960
rect 28080 34536 28132 34542
rect 28080 34478 28132 34484
rect 27988 34060 28040 34066
rect 27988 34002 28040 34008
rect 28080 33924 28132 33930
rect 28080 33866 28132 33872
rect 28092 33658 28120 33866
rect 28080 33652 28132 33658
rect 28080 33594 28132 33600
rect 28080 33448 28132 33454
rect 28080 33390 28132 33396
rect 27896 31816 27948 31822
rect 27896 31758 27948 31764
rect 27724 31726 27844 31754
rect 27526 31311 27582 31320
rect 27620 31340 27672 31346
rect 27620 31282 27672 31288
rect 27528 29708 27580 29714
rect 27528 29650 27580 29656
rect 27344 29572 27396 29578
rect 27344 29514 27396 29520
rect 27356 29306 27384 29514
rect 27344 29300 27396 29306
rect 27344 29242 27396 29248
rect 27540 28665 27568 29650
rect 27526 28656 27582 28665
rect 27436 28620 27488 28626
rect 27526 28591 27582 28600
rect 27436 28562 27488 28568
rect 27344 28484 27396 28490
rect 27344 28426 27396 28432
rect 27356 28218 27384 28426
rect 27344 28212 27396 28218
rect 27344 28154 27396 28160
rect 27252 28076 27304 28082
rect 27252 28018 27304 28024
rect 27448 26625 27476 28562
rect 27526 27568 27582 27577
rect 27526 27503 27528 27512
rect 27580 27503 27582 27512
rect 27528 27474 27580 27480
rect 27434 26616 27490 26625
rect 27434 26551 27490 26560
rect 27436 26036 27488 26042
rect 27436 25978 27488 25984
rect 27344 24132 27396 24138
rect 27344 24074 27396 24080
rect 27356 23866 27384 24074
rect 27344 23860 27396 23866
rect 27344 23802 27396 23808
rect 27252 23044 27304 23050
rect 27252 22986 27304 22992
rect 27264 22778 27292 22986
rect 27252 22772 27304 22778
rect 27252 22714 27304 22720
rect 27448 21554 27476 25978
rect 27632 23730 27660 31282
rect 27724 26994 27752 31726
rect 28092 30122 28120 33390
rect 28356 32904 28408 32910
rect 28356 32846 28408 32852
rect 28172 32836 28224 32842
rect 28172 32778 28224 32784
rect 28184 32026 28212 32778
rect 28368 32434 28396 32846
rect 28356 32428 28408 32434
rect 28356 32370 28408 32376
rect 28262 32056 28318 32065
rect 28172 32020 28224 32026
rect 28262 31991 28318 32000
rect 28172 31962 28224 31968
rect 28172 31816 28224 31822
rect 28172 31758 28224 31764
rect 28080 30116 28132 30122
rect 28080 30058 28132 30064
rect 27988 28076 28040 28082
rect 27988 28018 28040 28024
rect 27804 27396 27856 27402
rect 27804 27338 27856 27344
rect 27816 27130 27844 27338
rect 27804 27124 27856 27130
rect 27804 27066 27856 27072
rect 27712 26988 27764 26994
rect 27712 26930 27764 26936
rect 27712 25356 27764 25362
rect 27712 25298 27764 25304
rect 27724 24818 27752 25298
rect 27712 24812 27764 24818
rect 27712 24754 27764 24760
rect 27620 23724 27672 23730
rect 27620 23666 27672 23672
rect 27528 22092 27580 22098
rect 27528 22034 27580 22040
rect 27540 22001 27568 22034
rect 27526 21992 27582 22001
rect 27526 21927 27582 21936
rect 27896 21956 27948 21962
rect 27896 21898 27948 21904
rect 27908 21690 27936 21898
rect 27896 21684 27948 21690
rect 27896 21626 27948 21632
rect 27436 21548 27488 21554
rect 27436 21490 27488 21496
rect 27804 21548 27856 21554
rect 27804 21490 27856 21496
rect 27344 20868 27396 20874
rect 27344 20810 27396 20816
rect 27356 19514 27384 20810
rect 27344 19508 27396 19514
rect 27344 19450 27396 19456
rect 27252 19372 27304 19378
rect 27252 19314 27304 19320
rect 27160 16108 27212 16114
rect 27160 16050 27212 16056
rect 27172 13938 27200 16050
rect 27160 13932 27212 13938
rect 27160 13874 27212 13880
rect 27264 12850 27292 19314
rect 27344 18284 27396 18290
rect 27344 18226 27396 18232
rect 27356 17338 27384 18226
rect 27344 17332 27396 17338
rect 27344 17274 27396 17280
rect 27344 16584 27396 16590
rect 27342 16552 27344 16561
rect 27396 16552 27398 16561
rect 27342 16487 27398 16496
rect 27252 12844 27304 12850
rect 27252 12786 27304 12792
rect 27448 12434 27476 21490
rect 27712 21004 27764 21010
rect 27712 20946 27764 20952
rect 27724 19310 27752 20946
rect 27816 19378 27844 21490
rect 27896 20256 27948 20262
rect 27896 20198 27948 20204
rect 27908 19922 27936 20198
rect 27896 19916 27948 19922
rect 27896 19858 27948 19864
rect 28000 19394 28028 28018
rect 28080 27872 28132 27878
rect 28080 27814 28132 27820
rect 28092 27538 28120 27814
rect 28080 27532 28132 27538
rect 28080 27474 28132 27480
rect 28080 22432 28132 22438
rect 28080 22374 28132 22380
rect 28092 22098 28120 22374
rect 28080 22092 28132 22098
rect 28080 22034 28132 22040
rect 28184 21554 28212 31758
rect 28276 30802 28304 31991
rect 28460 31754 28488 35634
rect 28552 33522 28580 46378
rect 28734 45724 29042 45733
rect 28734 45722 28740 45724
rect 28796 45722 28820 45724
rect 28876 45722 28900 45724
rect 28956 45722 28980 45724
rect 29036 45722 29042 45724
rect 28796 45670 28798 45722
rect 28978 45670 28980 45722
rect 28734 45668 28740 45670
rect 28796 45668 28820 45670
rect 28876 45668 28900 45670
rect 28956 45668 28980 45670
rect 29036 45668 29042 45670
rect 28734 45659 29042 45668
rect 28734 44636 29042 44645
rect 28734 44634 28740 44636
rect 28796 44634 28820 44636
rect 28876 44634 28900 44636
rect 28956 44634 28980 44636
rect 29036 44634 29042 44636
rect 28796 44582 28798 44634
rect 28978 44582 28980 44634
rect 28734 44580 28740 44582
rect 28796 44580 28820 44582
rect 28876 44580 28900 44582
rect 28956 44580 28980 44582
rect 29036 44580 29042 44582
rect 28734 44571 29042 44580
rect 28734 43548 29042 43557
rect 28734 43546 28740 43548
rect 28796 43546 28820 43548
rect 28876 43546 28900 43548
rect 28956 43546 28980 43548
rect 29036 43546 29042 43548
rect 28796 43494 28798 43546
rect 28978 43494 28980 43546
rect 28734 43492 28740 43494
rect 28796 43492 28820 43494
rect 28876 43492 28900 43494
rect 28956 43492 28980 43494
rect 29036 43492 29042 43494
rect 28734 43483 29042 43492
rect 28734 42460 29042 42469
rect 28734 42458 28740 42460
rect 28796 42458 28820 42460
rect 28876 42458 28900 42460
rect 28956 42458 28980 42460
rect 29036 42458 29042 42460
rect 28796 42406 28798 42458
rect 28978 42406 28980 42458
rect 28734 42404 28740 42406
rect 28796 42404 28820 42406
rect 28876 42404 28900 42406
rect 28956 42404 28980 42406
rect 29036 42404 29042 42406
rect 28734 42395 29042 42404
rect 28734 41372 29042 41381
rect 28734 41370 28740 41372
rect 28796 41370 28820 41372
rect 28876 41370 28900 41372
rect 28956 41370 28980 41372
rect 29036 41370 29042 41372
rect 28796 41318 28798 41370
rect 28978 41318 28980 41370
rect 28734 41316 28740 41318
rect 28796 41316 28820 41318
rect 28876 41316 28900 41318
rect 28956 41316 28980 41318
rect 29036 41316 29042 41318
rect 28734 41307 29042 41316
rect 28630 40896 28686 40905
rect 28630 40831 28686 40840
rect 28644 39506 28672 40831
rect 28734 40284 29042 40293
rect 28734 40282 28740 40284
rect 28796 40282 28820 40284
rect 28876 40282 28900 40284
rect 28956 40282 28980 40284
rect 29036 40282 29042 40284
rect 28796 40230 28798 40282
rect 28978 40230 28980 40282
rect 28734 40228 28740 40230
rect 28796 40228 28820 40230
rect 28876 40228 28900 40230
rect 28956 40228 28980 40230
rect 29036 40228 29042 40230
rect 28734 40219 29042 40228
rect 28632 39500 28684 39506
rect 28632 39442 28684 39448
rect 28734 39196 29042 39205
rect 28734 39194 28740 39196
rect 28796 39194 28820 39196
rect 28876 39194 28900 39196
rect 28956 39194 28980 39196
rect 29036 39194 29042 39196
rect 28796 39142 28798 39194
rect 28978 39142 28980 39194
rect 28734 39140 28740 39142
rect 28796 39140 28820 39142
rect 28876 39140 28900 39142
rect 28956 39140 28980 39142
rect 29036 39140 29042 39142
rect 28734 39131 29042 39140
rect 28632 38956 28684 38962
rect 28632 38898 28684 38904
rect 28540 33516 28592 33522
rect 28540 33458 28592 33464
rect 28460 31726 28580 31754
rect 28264 30796 28316 30802
rect 28264 30738 28316 30744
rect 28356 30252 28408 30258
rect 28356 30194 28408 30200
rect 28368 30025 28396 30194
rect 28354 30016 28410 30025
rect 28354 29951 28410 29960
rect 28264 26988 28316 26994
rect 28264 26930 28316 26936
rect 28172 21548 28224 21554
rect 28172 21490 28224 21496
rect 27804 19372 27856 19378
rect 27804 19314 27856 19320
rect 27908 19366 28028 19394
rect 27712 19304 27764 19310
rect 27712 19246 27764 19252
rect 27528 18964 27580 18970
rect 27528 18906 27580 18912
rect 27540 17338 27568 18906
rect 27528 17332 27580 17338
rect 27528 17274 27580 17280
rect 27620 17128 27672 17134
rect 27620 17070 27672 17076
rect 27526 15736 27582 15745
rect 27526 15671 27582 15680
rect 27540 15570 27568 15671
rect 27528 15564 27580 15570
rect 27528 15506 27580 15512
rect 27528 15020 27580 15026
rect 27528 14962 27580 14968
rect 27540 13954 27568 14962
rect 27632 14074 27660 17070
rect 27908 16658 27936 19366
rect 27988 18692 28040 18698
rect 27988 18634 28040 18640
rect 28000 18426 28028 18634
rect 27988 18420 28040 18426
rect 27988 18362 28040 18368
rect 28172 17604 28224 17610
rect 28172 17546 28224 17552
rect 28184 16794 28212 17546
rect 28172 16788 28224 16794
rect 28172 16730 28224 16736
rect 27896 16652 27948 16658
rect 27896 16594 27948 16600
rect 28172 15904 28224 15910
rect 28172 15846 28224 15852
rect 28184 15570 28212 15846
rect 28172 15564 28224 15570
rect 28172 15506 28224 15512
rect 27896 14816 27948 14822
rect 27896 14758 27948 14764
rect 27908 14550 27936 14758
rect 27896 14544 27948 14550
rect 27896 14486 27948 14492
rect 27620 14068 27672 14074
rect 27620 14010 27672 14016
rect 27540 13926 27660 13954
rect 27356 12406 27476 12434
rect 27160 10464 27212 10470
rect 27160 10406 27212 10412
rect 27172 10198 27200 10406
rect 27160 10192 27212 10198
rect 27160 10134 27212 10140
rect 27356 6662 27384 12406
rect 27528 11212 27580 11218
rect 27528 11154 27580 11160
rect 27540 10305 27568 11154
rect 27526 10296 27582 10305
rect 27526 10231 27582 10240
rect 27632 9586 27660 13926
rect 28080 13388 28132 13394
rect 28080 13330 28132 13336
rect 27712 11076 27764 11082
rect 27712 11018 27764 11024
rect 27724 9654 27752 11018
rect 27712 9648 27764 9654
rect 27712 9590 27764 9596
rect 27620 9580 27672 9586
rect 27620 9522 27672 9528
rect 27526 8936 27582 8945
rect 27526 8871 27582 8880
rect 27540 7954 27568 8871
rect 27528 7948 27580 7954
rect 27528 7890 27580 7896
rect 27344 6656 27396 6662
rect 27344 6598 27396 6604
rect 27356 6322 27384 6598
rect 27344 6316 27396 6322
rect 27344 6258 27396 6264
rect 27068 5296 27120 5302
rect 27068 5238 27120 5244
rect 26424 5228 26476 5234
rect 26424 5170 26476 5176
rect 26608 5024 26660 5030
rect 26608 4966 26660 4972
rect 26620 3058 26648 4966
rect 27436 4684 27488 4690
rect 27436 4626 27488 4632
rect 27448 3505 27476 4626
rect 27632 3942 27660 9522
rect 27712 8492 27764 8498
rect 27712 8434 27764 8440
rect 27724 5846 27752 8434
rect 27712 5840 27764 5846
rect 27712 5782 27764 5788
rect 27724 4146 27752 5782
rect 27712 4140 27764 4146
rect 27712 4082 27764 4088
rect 27620 3936 27672 3942
rect 27620 3878 27672 3884
rect 27528 3596 27580 3602
rect 27528 3538 27580 3544
rect 27434 3496 27490 3505
rect 27252 3460 27304 3466
rect 27434 3431 27490 3440
rect 27252 3402 27304 3408
rect 27264 3194 27292 3402
rect 27252 3188 27304 3194
rect 27252 3130 27304 3136
rect 26608 3052 26660 3058
rect 26608 2994 26660 3000
rect 26148 2984 26200 2990
rect 26148 2926 26200 2932
rect 26160 2825 26188 2926
rect 26146 2816 26202 2825
rect 26146 2751 26202 2760
rect 25872 2644 25924 2650
rect 25872 2586 25924 2592
rect 27068 2440 27120 2446
rect 27068 2382 27120 2388
rect 27080 800 27108 2382
rect 27540 1465 27568 3538
rect 27632 3058 27660 3878
rect 27620 3052 27672 3058
rect 27620 2994 27672 3000
rect 27724 2774 27752 4082
rect 27804 3120 27856 3126
rect 27804 3062 27856 3068
rect 27632 2746 27752 2774
rect 27632 2446 27660 2746
rect 27816 2650 27844 3062
rect 27804 2644 27856 2650
rect 27804 2586 27856 2592
rect 28092 2553 28120 13330
rect 28172 8288 28224 8294
rect 28172 8230 28224 8236
rect 28184 7954 28212 8230
rect 28172 7948 28224 7954
rect 28172 7890 28224 7896
rect 28276 7410 28304 26930
rect 28354 25256 28410 25265
rect 28354 25191 28356 25200
rect 28408 25191 28410 25200
rect 28356 25162 28408 25168
rect 28354 24576 28410 24585
rect 28354 24511 28410 24520
rect 28368 24274 28396 24511
rect 28356 24268 28408 24274
rect 28356 24210 28408 24216
rect 28354 21176 28410 21185
rect 28354 21111 28410 21120
rect 28368 21010 28396 21111
rect 28356 21004 28408 21010
rect 28356 20946 28408 20952
rect 28354 20496 28410 20505
rect 28354 20431 28410 20440
rect 28368 19922 28396 20431
rect 28356 19916 28408 19922
rect 28356 19858 28408 19864
rect 28356 18760 28408 18766
rect 28356 18702 28408 18708
rect 28368 17746 28396 18702
rect 28356 17740 28408 17746
rect 28356 17682 28408 17688
rect 28356 15904 28408 15910
rect 28356 15846 28408 15852
rect 28368 15570 28396 15846
rect 28356 15564 28408 15570
rect 28356 15506 28408 15512
rect 28446 15056 28502 15065
rect 28446 14991 28502 15000
rect 28356 14408 28408 14414
rect 28354 14376 28356 14385
rect 28408 14376 28410 14385
rect 28354 14311 28410 14320
rect 28460 13938 28488 14991
rect 28448 13932 28500 13938
rect 28448 13874 28500 13880
rect 28354 12336 28410 12345
rect 28354 12271 28356 12280
rect 28408 12271 28410 12280
rect 28356 12242 28408 12248
rect 28356 11144 28408 11150
rect 28356 11086 28408 11092
rect 28368 10674 28396 11086
rect 28356 10668 28408 10674
rect 28356 10610 28408 10616
rect 28356 8968 28408 8974
rect 28356 8910 28408 8916
rect 28368 7954 28396 8910
rect 28552 8498 28580 31726
rect 28644 22642 28672 38898
rect 28734 38108 29042 38117
rect 28734 38106 28740 38108
rect 28796 38106 28820 38108
rect 28876 38106 28900 38108
rect 28956 38106 28980 38108
rect 29036 38106 29042 38108
rect 28796 38054 28798 38106
rect 28978 38054 28980 38106
rect 28734 38052 28740 38054
rect 28796 38052 28820 38054
rect 28876 38052 28900 38054
rect 28956 38052 28980 38054
rect 29036 38052 29042 38054
rect 28734 38043 29042 38052
rect 28734 37020 29042 37029
rect 28734 37018 28740 37020
rect 28796 37018 28820 37020
rect 28876 37018 28900 37020
rect 28956 37018 28980 37020
rect 29036 37018 29042 37020
rect 28796 36966 28798 37018
rect 28978 36966 28980 37018
rect 28734 36964 28740 36966
rect 28796 36964 28820 36966
rect 28876 36964 28900 36966
rect 28956 36964 28980 36966
rect 29036 36964 29042 36966
rect 28734 36955 29042 36964
rect 28734 35932 29042 35941
rect 28734 35930 28740 35932
rect 28796 35930 28820 35932
rect 28876 35930 28900 35932
rect 28956 35930 28980 35932
rect 29036 35930 29042 35932
rect 28796 35878 28798 35930
rect 28978 35878 28980 35930
rect 28734 35876 28740 35878
rect 28796 35876 28820 35878
rect 28876 35876 28900 35878
rect 28956 35876 28980 35878
rect 29036 35876 29042 35878
rect 28734 35867 29042 35876
rect 28734 34844 29042 34853
rect 28734 34842 28740 34844
rect 28796 34842 28820 34844
rect 28876 34842 28900 34844
rect 28956 34842 28980 34844
rect 29036 34842 29042 34844
rect 28796 34790 28798 34842
rect 28978 34790 28980 34842
rect 28734 34788 28740 34790
rect 28796 34788 28820 34790
rect 28876 34788 28900 34790
rect 28956 34788 28980 34790
rect 29036 34788 29042 34790
rect 28734 34779 29042 34788
rect 28734 33756 29042 33765
rect 28734 33754 28740 33756
rect 28796 33754 28820 33756
rect 28876 33754 28900 33756
rect 28956 33754 28980 33756
rect 29036 33754 29042 33756
rect 28796 33702 28798 33754
rect 28978 33702 28980 33754
rect 28734 33700 28740 33702
rect 28796 33700 28820 33702
rect 28876 33700 28900 33702
rect 28956 33700 28980 33702
rect 29036 33700 29042 33702
rect 28734 33691 29042 33700
rect 28734 32668 29042 32677
rect 28734 32666 28740 32668
rect 28796 32666 28820 32668
rect 28876 32666 28900 32668
rect 28956 32666 28980 32668
rect 29036 32666 29042 32668
rect 28796 32614 28798 32666
rect 28978 32614 28980 32666
rect 28734 32612 28740 32614
rect 28796 32612 28820 32614
rect 28876 32612 28900 32614
rect 28956 32612 28980 32614
rect 29036 32612 29042 32614
rect 28734 32603 29042 32612
rect 28734 31580 29042 31589
rect 28734 31578 28740 31580
rect 28796 31578 28820 31580
rect 28876 31578 28900 31580
rect 28956 31578 28980 31580
rect 29036 31578 29042 31580
rect 28796 31526 28798 31578
rect 28978 31526 28980 31578
rect 28734 31524 28740 31526
rect 28796 31524 28820 31526
rect 28876 31524 28900 31526
rect 28956 31524 28980 31526
rect 29036 31524 29042 31526
rect 28734 31515 29042 31524
rect 28734 30492 29042 30501
rect 28734 30490 28740 30492
rect 28796 30490 28820 30492
rect 28876 30490 28900 30492
rect 28956 30490 28980 30492
rect 29036 30490 29042 30492
rect 28796 30438 28798 30490
rect 28978 30438 28980 30490
rect 28734 30436 28740 30438
rect 28796 30436 28820 30438
rect 28876 30436 28900 30438
rect 28956 30436 28980 30438
rect 29036 30436 29042 30438
rect 28734 30427 29042 30436
rect 28734 29404 29042 29413
rect 28734 29402 28740 29404
rect 28796 29402 28820 29404
rect 28876 29402 28900 29404
rect 28956 29402 28980 29404
rect 29036 29402 29042 29404
rect 28796 29350 28798 29402
rect 28978 29350 28980 29402
rect 28734 29348 28740 29350
rect 28796 29348 28820 29350
rect 28876 29348 28900 29350
rect 28956 29348 28980 29350
rect 29036 29348 29042 29350
rect 28734 29339 29042 29348
rect 28734 28316 29042 28325
rect 28734 28314 28740 28316
rect 28796 28314 28820 28316
rect 28876 28314 28900 28316
rect 28956 28314 28980 28316
rect 29036 28314 29042 28316
rect 28796 28262 28798 28314
rect 28978 28262 28980 28314
rect 28734 28260 28740 28262
rect 28796 28260 28820 28262
rect 28876 28260 28900 28262
rect 28956 28260 28980 28262
rect 29036 28260 29042 28262
rect 28734 28251 29042 28260
rect 28734 27228 29042 27237
rect 28734 27226 28740 27228
rect 28796 27226 28820 27228
rect 28876 27226 28900 27228
rect 28956 27226 28980 27228
rect 29036 27226 29042 27228
rect 28796 27174 28798 27226
rect 28978 27174 28980 27226
rect 28734 27172 28740 27174
rect 28796 27172 28820 27174
rect 28876 27172 28900 27174
rect 28956 27172 28980 27174
rect 29036 27172 29042 27174
rect 28734 27163 29042 27172
rect 28734 26140 29042 26149
rect 28734 26138 28740 26140
rect 28796 26138 28820 26140
rect 28876 26138 28900 26140
rect 28956 26138 28980 26140
rect 29036 26138 29042 26140
rect 28796 26086 28798 26138
rect 28978 26086 28980 26138
rect 28734 26084 28740 26086
rect 28796 26084 28820 26086
rect 28876 26084 28900 26086
rect 28956 26084 28980 26086
rect 29036 26084 29042 26086
rect 28734 26075 29042 26084
rect 28734 25052 29042 25061
rect 28734 25050 28740 25052
rect 28796 25050 28820 25052
rect 28876 25050 28900 25052
rect 28956 25050 28980 25052
rect 29036 25050 29042 25052
rect 28796 24998 28798 25050
rect 28978 24998 28980 25050
rect 28734 24996 28740 24998
rect 28796 24996 28820 24998
rect 28876 24996 28900 24998
rect 28956 24996 28980 24998
rect 29036 24996 29042 24998
rect 28734 24987 29042 24996
rect 28734 23964 29042 23973
rect 28734 23962 28740 23964
rect 28796 23962 28820 23964
rect 28876 23962 28900 23964
rect 28956 23962 28980 23964
rect 29036 23962 29042 23964
rect 28796 23910 28798 23962
rect 28978 23910 28980 23962
rect 28734 23908 28740 23910
rect 28796 23908 28820 23910
rect 28876 23908 28900 23910
rect 28956 23908 28980 23910
rect 29036 23908 29042 23910
rect 28734 23899 29042 23908
rect 29918 23896 29974 23905
rect 29918 23831 29974 23840
rect 29932 23186 29960 23831
rect 29920 23180 29972 23186
rect 29920 23122 29972 23128
rect 28734 22876 29042 22885
rect 28734 22874 28740 22876
rect 28796 22874 28820 22876
rect 28876 22874 28900 22876
rect 28956 22874 28980 22876
rect 29036 22874 29042 22876
rect 28796 22822 28798 22874
rect 28978 22822 28980 22874
rect 28734 22820 28740 22822
rect 28796 22820 28820 22822
rect 28876 22820 28900 22822
rect 28956 22820 28980 22822
rect 29036 22820 29042 22822
rect 28734 22811 29042 22820
rect 28632 22636 28684 22642
rect 28632 22578 28684 22584
rect 28734 21788 29042 21797
rect 28734 21786 28740 21788
rect 28796 21786 28820 21788
rect 28876 21786 28900 21788
rect 28956 21786 28980 21788
rect 29036 21786 29042 21788
rect 28796 21734 28798 21786
rect 28978 21734 28980 21786
rect 28734 21732 28740 21734
rect 28796 21732 28820 21734
rect 28876 21732 28900 21734
rect 28956 21732 28980 21734
rect 29036 21732 29042 21734
rect 28734 21723 29042 21732
rect 28734 20700 29042 20709
rect 28734 20698 28740 20700
rect 28796 20698 28820 20700
rect 28876 20698 28900 20700
rect 28956 20698 28980 20700
rect 29036 20698 29042 20700
rect 28796 20646 28798 20698
rect 28978 20646 28980 20698
rect 28734 20644 28740 20646
rect 28796 20644 28820 20646
rect 28876 20644 28900 20646
rect 28956 20644 28980 20646
rect 29036 20644 29042 20646
rect 28734 20635 29042 20644
rect 28734 19612 29042 19621
rect 28734 19610 28740 19612
rect 28796 19610 28820 19612
rect 28876 19610 28900 19612
rect 28956 19610 28980 19612
rect 29036 19610 29042 19612
rect 28796 19558 28798 19610
rect 28978 19558 28980 19610
rect 28734 19556 28740 19558
rect 28796 19556 28820 19558
rect 28876 19556 28900 19558
rect 28956 19556 28980 19558
rect 29036 19556 29042 19558
rect 28734 19547 29042 19556
rect 28734 18524 29042 18533
rect 28734 18522 28740 18524
rect 28796 18522 28820 18524
rect 28876 18522 28900 18524
rect 28956 18522 28980 18524
rect 29036 18522 29042 18524
rect 28796 18470 28798 18522
rect 28978 18470 28980 18522
rect 28734 18468 28740 18470
rect 28796 18468 28820 18470
rect 28876 18468 28900 18470
rect 28956 18468 28980 18470
rect 29036 18468 29042 18470
rect 28734 18459 29042 18468
rect 28734 17436 29042 17445
rect 28734 17434 28740 17436
rect 28796 17434 28820 17436
rect 28876 17434 28900 17436
rect 28956 17434 28980 17436
rect 29036 17434 29042 17436
rect 28796 17382 28798 17434
rect 28978 17382 28980 17434
rect 28734 17380 28740 17382
rect 28796 17380 28820 17382
rect 28876 17380 28900 17382
rect 28956 17380 28980 17382
rect 29036 17380 29042 17382
rect 28734 17371 29042 17380
rect 28734 16348 29042 16357
rect 28734 16346 28740 16348
rect 28796 16346 28820 16348
rect 28876 16346 28900 16348
rect 28956 16346 28980 16348
rect 29036 16346 29042 16348
rect 28796 16294 28798 16346
rect 28978 16294 28980 16346
rect 28734 16292 28740 16294
rect 28796 16292 28820 16294
rect 28876 16292 28900 16294
rect 28956 16292 28980 16294
rect 29036 16292 29042 16294
rect 28734 16283 29042 16292
rect 28734 15260 29042 15269
rect 28734 15258 28740 15260
rect 28796 15258 28820 15260
rect 28876 15258 28900 15260
rect 28956 15258 28980 15260
rect 29036 15258 29042 15260
rect 28796 15206 28798 15258
rect 28978 15206 28980 15258
rect 28734 15204 28740 15206
rect 28796 15204 28820 15206
rect 28876 15204 28900 15206
rect 28956 15204 28980 15206
rect 29036 15204 29042 15206
rect 28734 15195 29042 15204
rect 28734 14172 29042 14181
rect 28734 14170 28740 14172
rect 28796 14170 28820 14172
rect 28876 14170 28900 14172
rect 28956 14170 28980 14172
rect 29036 14170 29042 14172
rect 28796 14118 28798 14170
rect 28978 14118 28980 14170
rect 28734 14116 28740 14118
rect 28796 14116 28820 14118
rect 28876 14116 28900 14118
rect 28956 14116 28980 14118
rect 29036 14116 29042 14118
rect 28734 14107 29042 14116
rect 28734 13084 29042 13093
rect 28734 13082 28740 13084
rect 28796 13082 28820 13084
rect 28876 13082 28900 13084
rect 28956 13082 28980 13084
rect 29036 13082 29042 13084
rect 28796 13030 28798 13082
rect 28978 13030 28980 13082
rect 28734 13028 28740 13030
rect 28796 13028 28820 13030
rect 28876 13028 28900 13030
rect 28956 13028 28980 13030
rect 29036 13028 29042 13030
rect 28734 13019 29042 13028
rect 28734 11996 29042 12005
rect 28734 11994 28740 11996
rect 28796 11994 28820 11996
rect 28876 11994 28900 11996
rect 28956 11994 28980 11996
rect 29036 11994 29042 11996
rect 28796 11942 28798 11994
rect 28978 11942 28980 11994
rect 28734 11940 28740 11942
rect 28796 11940 28820 11942
rect 28876 11940 28900 11942
rect 28956 11940 28980 11942
rect 29036 11940 29042 11942
rect 28734 11931 29042 11940
rect 29918 10976 29974 10985
rect 28734 10908 29042 10917
rect 29918 10911 29974 10920
rect 28734 10906 28740 10908
rect 28796 10906 28820 10908
rect 28876 10906 28900 10908
rect 28956 10906 28980 10908
rect 29036 10906 29042 10908
rect 28796 10854 28798 10906
rect 28978 10854 28980 10906
rect 28734 10852 28740 10854
rect 28796 10852 28820 10854
rect 28876 10852 28900 10854
rect 28956 10852 28980 10854
rect 29036 10852 29042 10854
rect 28734 10843 29042 10852
rect 29932 10130 29960 10911
rect 29920 10124 29972 10130
rect 29920 10066 29972 10072
rect 28734 9820 29042 9829
rect 28734 9818 28740 9820
rect 28796 9818 28820 9820
rect 28876 9818 28900 9820
rect 28956 9818 28980 9820
rect 29036 9818 29042 9820
rect 28796 9766 28798 9818
rect 28978 9766 28980 9818
rect 28734 9764 28740 9766
rect 28796 9764 28820 9766
rect 28876 9764 28900 9766
rect 28956 9764 28980 9766
rect 29036 9764 29042 9766
rect 28734 9755 29042 9764
rect 29920 8900 29972 8906
rect 29920 8842 29972 8848
rect 28734 8732 29042 8741
rect 28734 8730 28740 8732
rect 28796 8730 28820 8732
rect 28876 8730 28900 8732
rect 28956 8730 28980 8732
rect 29036 8730 29042 8732
rect 28796 8678 28798 8730
rect 28978 8678 28980 8730
rect 28734 8676 28740 8678
rect 28796 8676 28820 8678
rect 28876 8676 28900 8678
rect 28956 8676 28980 8678
rect 29036 8676 29042 8678
rect 28734 8667 29042 8676
rect 28540 8492 28592 8498
rect 28540 8434 28592 8440
rect 28356 7948 28408 7954
rect 28356 7890 28408 7896
rect 28734 7644 29042 7653
rect 28734 7642 28740 7644
rect 28796 7642 28820 7644
rect 28876 7642 28900 7644
rect 28956 7642 28980 7644
rect 29036 7642 29042 7644
rect 28796 7590 28798 7642
rect 28978 7590 28980 7642
rect 28734 7588 28740 7590
rect 28796 7588 28820 7590
rect 28876 7588 28900 7590
rect 28956 7588 28980 7590
rect 29036 7588 29042 7590
rect 28734 7579 29042 7588
rect 29932 7585 29960 8842
rect 29918 7576 29974 7585
rect 29918 7511 29974 7520
rect 28264 7404 28316 7410
rect 28264 7346 28316 7352
rect 28734 6556 29042 6565
rect 28734 6554 28740 6556
rect 28796 6554 28820 6556
rect 28876 6554 28900 6556
rect 28956 6554 28980 6556
rect 29036 6554 29042 6556
rect 28796 6502 28798 6554
rect 28978 6502 28980 6554
rect 28734 6500 28740 6502
rect 28796 6500 28820 6502
rect 28876 6500 28900 6502
rect 28956 6500 28980 6502
rect 29036 6500 29042 6502
rect 28734 6491 29042 6500
rect 29920 5636 29972 5642
rect 29920 5578 29972 5584
rect 29932 5545 29960 5578
rect 29918 5536 29974 5545
rect 28734 5468 29042 5477
rect 29918 5471 29974 5480
rect 28734 5466 28740 5468
rect 28796 5466 28820 5468
rect 28876 5466 28900 5468
rect 28956 5466 28980 5468
rect 29036 5466 29042 5468
rect 28796 5414 28798 5466
rect 28978 5414 28980 5466
rect 28734 5412 28740 5414
rect 28796 5412 28820 5414
rect 28876 5412 28900 5414
rect 28956 5412 28980 5414
rect 29036 5412 29042 5414
rect 28734 5403 29042 5412
rect 28356 4616 28408 4622
rect 28356 4558 28408 4564
rect 28172 4548 28224 4554
rect 28172 4490 28224 4496
rect 28184 4282 28212 4490
rect 28172 4276 28224 4282
rect 28172 4218 28224 4224
rect 28368 3058 28396 4558
rect 28734 4380 29042 4389
rect 28734 4378 28740 4380
rect 28796 4378 28820 4380
rect 28876 4378 28900 4380
rect 28956 4378 28980 4380
rect 29036 4378 29042 4380
rect 28796 4326 28798 4378
rect 28978 4326 28980 4378
rect 28734 4324 28740 4326
rect 28796 4324 28820 4326
rect 28876 4324 28900 4326
rect 28956 4324 28980 4326
rect 29036 4324 29042 4326
rect 28734 4315 29042 4324
rect 28734 3292 29042 3301
rect 28734 3290 28740 3292
rect 28796 3290 28820 3292
rect 28876 3290 28900 3292
rect 28956 3290 28980 3292
rect 29036 3290 29042 3292
rect 28796 3238 28798 3290
rect 28978 3238 28980 3290
rect 28734 3236 28740 3238
rect 28796 3236 28820 3238
rect 28876 3236 28900 3238
rect 28956 3236 28980 3238
rect 29036 3236 29042 3238
rect 28734 3227 29042 3236
rect 28356 3052 28408 3058
rect 28356 2994 28408 3000
rect 28078 2544 28134 2553
rect 28078 2479 28134 2488
rect 27620 2440 27672 2446
rect 27620 2382 27672 2388
rect 28734 2204 29042 2213
rect 28734 2202 28740 2204
rect 28796 2202 28820 2204
rect 28876 2202 28900 2204
rect 28956 2202 28980 2204
rect 29036 2202 29042 2204
rect 28796 2150 28798 2202
rect 28978 2150 28980 2202
rect 28734 2148 28740 2150
rect 28796 2148 28820 2150
rect 28876 2148 28900 2150
rect 28956 2148 28980 2150
rect 29036 2148 29042 2150
rect 28734 2139 29042 2148
rect 27526 1456 27582 1465
rect 27526 1391 27582 1400
rect -10 200 102 800
rect 634 200 746 800
rect 1278 200 1390 800
rect 1922 200 2034 800
rect 2566 200 2678 800
rect 3210 200 3322 800
rect 3854 200 3966 800
rect 4498 200 4610 800
rect 5786 200 5898 800
rect 6430 200 6542 800
rect 7074 200 7186 800
rect 7718 200 7830 800
rect 8362 200 8474 800
rect 9006 200 9118 800
rect 9650 200 9762 800
rect 10938 200 11050 800
rect 11582 200 11694 800
rect 12226 200 12338 800
rect 12870 200 12982 800
rect 13514 200 13626 800
rect 14158 200 14270 800
rect 14802 200 14914 800
rect 16090 200 16202 800
rect 16734 200 16846 800
rect 17378 200 17490 800
rect 18022 200 18134 800
rect 18666 200 18778 800
rect 19310 200 19422 800
rect 19954 200 20066 800
rect 21242 200 21354 800
rect 21886 200 21998 800
rect 22530 200 22642 800
rect 23174 200 23286 800
rect 23818 200 23930 800
rect 24462 200 24574 800
rect 25106 200 25218 800
rect 26394 200 26506 800
rect 27038 200 27150 800
rect 27682 200 27794 800
rect 28326 200 28438 800
rect 28970 200 29082 800
rect 29614 200 29726 800
<< via2 >>
rect 3514 49680 3570 49736
rect 2778 44920 2834 44976
rect 1582 41556 1584 41576
rect 1584 41556 1636 41576
rect 1636 41556 1638 41576
rect 1582 41520 1638 41556
rect 1582 37440 1638 37496
rect 1582 29960 1638 30016
rect 1582 27920 1638 27976
rect 1582 25200 1638 25256
rect 2778 42200 2834 42256
rect 2778 38800 2834 38856
rect 2870 36760 2926 36816
rect 1582 18400 1638 18456
rect 1582 13640 1638 13696
rect 2778 36080 2834 36136
rect 4429 47354 4485 47356
rect 4509 47354 4565 47356
rect 4589 47354 4645 47356
rect 4669 47354 4725 47356
rect 4429 47302 4475 47354
rect 4475 47302 4485 47354
rect 4509 47302 4539 47354
rect 4539 47302 4551 47354
rect 4551 47302 4565 47354
rect 4589 47302 4603 47354
rect 4603 47302 4615 47354
rect 4615 47302 4645 47354
rect 4669 47302 4679 47354
rect 4679 47302 4725 47354
rect 4429 47300 4485 47302
rect 4509 47300 4565 47302
rect 4589 47300 4645 47302
rect 4669 47300 4725 47302
rect 4429 46266 4485 46268
rect 4509 46266 4565 46268
rect 4589 46266 4645 46268
rect 4669 46266 4725 46268
rect 4429 46214 4475 46266
rect 4475 46214 4485 46266
rect 4509 46214 4539 46266
rect 4539 46214 4551 46266
rect 4551 46214 4565 46266
rect 4589 46214 4603 46266
rect 4603 46214 4615 46266
rect 4615 46214 4645 46266
rect 4669 46214 4679 46266
rect 4679 46214 4725 46266
rect 4429 46212 4485 46214
rect 4509 46212 4565 46214
rect 4589 46212 4645 46214
rect 4669 46212 4725 46214
rect 4429 45178 4485 45180
rect 4509 45178 4565 45180
rect 4589 45178 4645 45180
rect 4669 45178 4725 45180
rect 4429 45126 4475 45178
rect 4475 45126 4485 45178
rect 4509 45126 4539 45178
rect 4539 45126 4551 45178
rect 4551 45126 4565 45178
rect 4589 45126 4603 45178
rect 4603 45126 4615 45178
rect 4615 45126 4645 45178
rect 4669 45126 4679 45178
rect 4679 45126 4725 45178
rect 4429 45124 4485 45126
rect 4509 45124 4565 45126
rect 4589 45124 4645 45126
rect 4669 45124 4725 45126
rect 4158 44240 4214 44296
rect 4429 44090 4485 44092
rect 4509 44090 4565 44092
rect 4589 44090 4645 44092
rect 4669 44090 4725 44092
rect 4429 44038 4475 44090
rect 4475 44038 4485 44090
rect 4509 44038 4539 44090
rect 4539 44038 4551 44090
rect 4551 44038 4565 44090
rect 4589 44038 4603 44090
rect 4603 44038 4615 44090
rect 4615 44038 4645 44090
rect 4669 44038 4679 44090
rect 4679 44038 4725 44090
rect 4429 44036 4485 44038
rect 4509 44036 4565 44038
rect 4589 44036 4645 44038
rect 4669 44036 4725 44038
rect 4429 43002 4485 43004
rect 4509 43002 4565 43004
rect 4589 43002 4645 43004
rect 4669 43002 4725 43004
rect 4429 42950 4475 43002
rect 4475 42950 4485 43002
rect 4509 42950 4539 43002
rect 4539 42950 4551 43002
rect 4551 42950 4565 43002
rect 4589 42950 4603 43002
rect 4603 42950 4615 43002
rect 4615 42950 4645 43002
rect 4669 42950 4679 43002
rect 4679 42950 4725 43002
rect 4429 42948 4485 42950
rect 4509 42948 4565 42950
rect 4589 42948 4645 42950
rect 4669 42948 4725 42950
rect 4429 41914 4485 41916
rect 4509 41914 4565 41916
rect 4589 41914 4645 41916
rect 4669 41914 4725 41916
rect 4429 41862 4475 41914
rect 4475 41862 4485 41914
rect 4509 41862 4539 41914
rect 4539 41862 4551 41914
rect 4551 41862 4565 41914
rect 4589 41862 4603 41914
rect 4603 41862 4615 41914
rect 4615 41862 4645 41914
rect 4669 41862 4679 41914
rect 4679 41862 4725 41914
rect 4429 41860 4485 41862
rect 4509 41860 4565 41862
rect 4589 41860 4645 41862
rect 4669 41860 4725 41862
rect 4429 40826 4485 40828
rect 4509 40826 4565 40828
rect 4589 40826 4645 40828
rect 4669 40826 4725 40828
rect 4429 40774 4475 40826
rect 4475 40774 4485 40826
rect 4509 40774 4539 40826
rect 4539 40774 4551 40826
rect 4551 40774 4565 40826
rect 4589 40774 4603 40826
rect 4603 40774 4615 40826
rect 4615 40774 4645 40826
rect 4669 40774 4679 40826
rect 4679 40774 4725 40826
rect 4429 40772 4485 40774
rect 4509 40772 4565 40774
rect 4589 40772 4645 40774
rect 4669 40772 4725 40774
rect 4429 39738 4485 39740
rect 4509 39738 4565 39740
rect 4589 39738 4645 39740
rect 4669 39738 4725 39740
rect 4429 39686 4475 39738
rect 4475 39686 4485 39738
rect 4509 39686 4539 39738
rect 4539 39686 4551 39738
rect 4551 39686 4565 39738
rect 4589 39686 4603 39738
rect 4603 39686 4615 39738
rect 4615 39686 4645 39738
rect 4669 39686 4679 39738
rect 4679 39686 4725 39738
rect 4429 39684 4485 39686
rect 4509 39684 4565 39686
rect 4589 39684 4645 39686
rect 4669 39684 4725 39686
rect 4429 38650 4485 38652
rect 4509 38650 4565 38652
rect 4589 38650 4645 38652
rect 4669 38650 4725 38652
rect 4429 38598 4475 38650
rect 4475 38598 4485 38650
rect 4509 38598 4539 38650
rect 4539 38598 4551 38650
rect 4551 38598 4565 38650
rect 4589 38598 4603 38650
rect 4603 38598 4615 38650
rect 4615 38598 4645 38650
rect 4669 38598 4679 38650
rect 4679 38598 4725 38650
rect 4429 38596 4485 38598
rect 4509 38596 4565 38598
rect 4589 38596 4645 38598
rect 4669 38596 4725 38598
rect 4429 37562 4485 37564
rect 4509 37562 4565 37564
rect 4589 37562 4645 37564
rect 4669 37562 4725 37564
rect 4429 37510 4475 37562
rect 4475 37510 4485 37562
rect 4509 37510 4539 37562
rect 4539 37510 4551 37562
rect 4551 37510 4565 37562
rect 4589 37510 4603 37562
rect 4603 37510 4615 37562
rect 4615 37510 4645 37562
rect 4669 37510 4679 37562
rect 4679 37510 4725 37562
rect 4429 37508 4485 37510
rect 4509 37508 4565 37510
rect 4589 37508 4645 37510
rect 4669 37508 4725 37510
rect 2778 34720 2834 34776
rect 4429 36474 4485 36476
rect 4509 36474 4565 36476
rect 4589 36474 4645 36476
rect 4669 36474 4725 36476
rect 4429 36422 4475 36474
rect 4475 36422 4485 36474
rect 4509 36422 4539 36474
rect 4539 36422 4551 36474
rect 4551 36422 4565 36474
rect 4589 36422 4603 36474
rect 4603 36422 4615 36474
rect 4615 36422 4645 36474
rect 4669 36422 4679 36474
rect 4679 36422 4725 36474
rect 4429 36420 4485 36422
rect 4509 36420 4565 36422
rect 4589 36420 4645 36422
rect 4669 36420 4725 36422
rect 4429 35386 4485 35388
rect 4509 35386 4565 35388
rect 4589 35386 4645 35388
rect 4669 35386 4725 35388
rect 4429 35334 4475 35386
rect 4475 35334 4485 35386
rect 4509 35334 4539 35386
rect 4539 35334 4551 35386
rect 4551 35334 4565 35386
rect 4589 35334 4603 35386
rect 4603 35334 4615 35386
rect 4615 35334 4645 35386
rect 4669 35334 4679 35386
rect 4679 35334 4725 35386
rect 4429 35332 4485 35334
rect 4509 35332 4565 35334
rect 4589 35332 4645 35334
rect 4669 35332 4725 35334
rect 3514 33360 3570 33416
rect 2962 32000 3018 32056
rect 2778 25880 2834 25936
rect 2778 19760 2834 19816
rect 3330 19080 3386 19136
rect 2778 17740 2834 17776
rect 2778 17720 2780 17740
rect 2780 17720 2832 17740
rect 2832 17720 2834 17740
rect 2778 15680 2834 15736
rect 2778 14320 2834 14376
rect 3606 12280 3662 12336
rect 2778 11636 2780 11656
rect 2780 11636 2832 11656
rect 2832 11636 2834 11656
rect 2778 11600 2834 11636
rect 2778 8880 2834 8936
rect 2778 7520 2834 7576
rect 4429 34298 4485 34300
rect 4509 34298 4565 34300
rect 4589 34298 4645 34300
rect 4669 34298 4725 34300
rect 4429 34246 4475 34298
rect 4475 34246 4485 34298
rect 4509 34246 4539 34298
rect 4539 34246 4551 34298
rect 4551 34246 4565 34298
rect 4589 34246 4603 34298
rect 4603 34246 4615 34298
rect 4615 34246 4645 34298
rect 4669 34246 4679 34298
rect 4679 34246 4725 34298
rect 4429 34244 4485 34246
rect 4509 34244 4565 34246
rect 4589 34244 4645 34246
rect 4669 34244 4725 34246
rect 4429 33210 4485 33212
rect 4509 33210 4565 33212
rect 4589 33210 4645 33212
rect 4669 33210 4725 33212
rect 4429 33158 4475 33210
rect 4475 33158 4485 33210
rect 4509 33158 4539 33210
rect 4539 33158 4551 33210
rect 4551 33158 4565 33210
rect 4589 33158 4603 33210
rect 4603 33158 4615 33210
rect 4615 33158 4645 33210
rect 4669 33158 4679 33210
rect 4679 33158 4725 33210
rect 4429 33156 4485 33158
rect 4509 33156 4565 33158
rect 4589 33156 4645 33158
rect 4669 33156 4725 33158
rect 4429 32122 4485 32124
rect 4509 32122 4565 32124
rect 4589 32122 4645 32124
rect 4669 32122 4725 32124
rect 4429 32070 4475 32122
rect 4475 32070 4485 32122
rect 4509 32070 4539 32122
rect 4539 32070 4551 32122
rect 4551 32070 4565 32122
rect 4589 32070 4603 32122
rect 4603 32070 4615 32122
rect 4615 32070 4645 32122
rect 4669 32070 4679 32122
rect 4679 32070 4725 32122
rect 4429 32068 4485 32070
rect 4509 32068 4565 32070
rect 4589 32068 4645 32070
rect 4669 32068 4725 32070
rect 4429 31034 4485 31036
rect 4509 31034 4565 31036
rect 4589 31034 4645 31036
rect 4669 31034 4725 31036
rect 4429 30982 4475 31034
rect 4475 30982 4485 31034
rect 4509 30982 4539 31034
rect 4539 30982 4551 31034
rect 4551 30982 4565 31034
rect 4589 30982 4603 31034
rect 4603 30982 4615 31034
rect 4615 30982 4645 31034
rect 4669 30982 4679 31034
rect 4679 30982 4725 31034
rect 4429 30980 4485 30982
rect 4509 30980 4565 30982
rect 4589 30980 4645 30982
rect 4669 30980 4725 30982
rect 4429 29946 4485 29948
rect 4509 29946 4565 29948
rect 4589 29946 4645 29948
rect 4669 29946 4725 29948
rect 4429 29894 4475 29946
rect 4475 29894 4485 29946
rect 4509 29894 4539 29946
rect 4539 29894 4551 29946
rect 4551 29894 4565 29946
rect 4589 29894 4603 29946
rect 4603 29894 4615 29946
rect 4615 29894 4645 29946
rect 4669 29894 4679 29946
rect 4679 29894 4725 29946
rect 4429 29892 4485 29894
rect 4509 29892 4565 29894
rect 4589 29892 4645 29894
rect 4669 29892 4725 29894
rect 4429 28858 4485 28860
rect 4509 28858 4565 28860
rect 4589 28858 4645 28860
rect 4669 28858 4725 28860
rect 4429 28806 4475 28858
rect 4475 28806 4485 28858
rect 4509 28806 4539 28858
rect 4539 28806 4551 28858
rect 4551 28806 4565 28858
rect 4589 28806 4603 28858
rect 4603 28806 4615 28858
rect 4615 28806 4645 28858
rect 4669 28806 4679 28858
rect 4679 28806 4725 28858
rect 4429 28804 4485 28806
rect 4509 28804 4565 28806
rect 4589 28804 4645 28806
rect 4669 28804 4725 28806
rect 4429 27770 4485 27772
rect 4509 27770 4565 27772
rect 4589 27770 4645 27772
rect 4669 27770 4725 27772
rect 4429 27718 4475 27770
rect 4475 27718 4485 27770
rect 4509 27718 4539 27770
rect 4539 27718 4551 27770
rect 4551 27718 4565 27770
rect 4589 27718 4603 27770
rect 4603 27718 4615 27770
rect 4615 27718 4645 27770
rect 4669 27718 4679 27770
rect 4679 27718 4725 27770
rect 4429 27716 4485 27718
rect 4509 27716 4565 27718
rect 4589 27716 4645 27718
rect 4669 27716 4725 27718
rect 7902 46810 7958 46812
rect 7982 46810 8038 46812
rect 8062 46810 8118 46812
rect 8142 46810 8198 46812
rect 7902 46758 7948 46810
rect 7948 46758 7958 46810
rect 7982 46758 8012 46810
rect 8012 46758 8024 46810
rect 8024 46758 8038 46810
rect 8062 46758 8076 46810
rect 8076 46758 8088 46810
rect 8088 46758 8118 46810
rect 8142 46758 8152 46810
rect 8152 46758 8198 46810
rect 7902 46756 7958 46758
rect 7982 46756 8038 46758
rect 8062 46756 8118 46758
rect 8142 46756 8198 46758
rect 7902 45722 7958 45724
rect 7982 45722 8038 45724
rect 8062 45722 8118 45724
rect 8142 45722 8198 45724
rect 7902 45670 7948 45722
rect 7948 45670 7958 45722
rect 7982 45670 8012 45722
rect 8012 45670 8024 45722
rect 8024 45670 8038 45722
rect 8062 45670 8076 45722
rect 8076 45670 8088 45722
rect 8088 45670 8118 45722
rect 8142 45670 8152 45722
rect 8152 45670 8198 45722
rect 7902 45668 7958 45670
rect 7982 45668 8038 45670
rect 8062 45668 8118 45670
rect 8142 45668 8198 45670
rect 11375 47354 11431 47356
rect 11455 47354 11511 47356
rect 11535 47354 11591 47356
rect 11615 47354 11671 47356
rect 11375 47302 11421 47354
rect 11421 47302 11431 47354
rect 11455 47302 11485 47354
rect 11485 47302 11497 47354
rect 11497 47302 11511 47354
rect 11535 47302 11549 47354
rect 11549 47302 11561 47354
rect 11561 47302 11591 47354
rect 11615 47302 11625 47354
rect 11625 47302 11671 47354
rect 11375 47300 11431 47302
rect 11455 47300 11511 47302
rect 11535 47300 11591 47302
rect 11615 47300 11671 47302
rect 11375 46266 11431 46268
rect 11455 46266 11511 46268
rect 11535 46266 11591 46268
rect 11615 46266 11671 46268
rect 11375 46214 11421 46266
rect 11421 46214 11431 46266
rect 11455 46214 11485 46266
rect 11485 46214 11497 46266
rect 11497 46214 11511 46266
rect 11535 46214 11549 46266
rect 11549 46214 11561 46266
rect 11561 46214 11591 46266
rect 11615 46214 11625 46266
rect 11625 46214 11671 46266
rect 11375 46212 11431 46214
rect 11455 46212 11511 46214
rect 11535 46212 11591 46214
rect 11615 46212 11671 46214
rect 14848 46810 14904 46812
rect 14928 46810 14984 46812
rect 15008 46810 15064 46812
rect 15088 46810 15144 46812
rect 14848 46758 14894 46810
rect 14894 46758 14904 46810
rect 14928 46758 14958 46810
rect 14958 46758 14970 46810
rect 14970 46758 14984 46810
rect 15008 46758 15022 46810
rect 15022 46758 15034 46810
rect 15034 46758 15064 46810
rect 15088 46758 15098 46810
rect 15098 46758 15144 46810
rect 14848 46756 14904 46758
rect 14928 46756 14984 46758
rect 15008 46756 15064 46758
rect 15088 46756 15144 46758
rect 7902 44634 7958 44636
rect 7982 44634 8038 44636
rect 8062 44634 8118 44636
rect 8142 44634 8198 44636
rect 7902 44582 7948 44634
rect 7948 44582 7958 44634
rect 7982 44582 8012 44634
rect 8012 44582 8024 44634
rect 8024 44582 8038 44634
rect 8062 44582 8076 44634
rect 8076 44582 8088 44634
rect 8088 44582 8118 44634
rect 8142 44582 8152 44634
rect 8152 44582 8198 44634
rect 7902 44580 7958 44582
rect 7982 44580 8038 44582
rect 8062 44580 8118 44582
rect 8142 44580 8198 44582
rect 11375 45178 11431 45180
rect 11455 45178 11511 45180
rect 11535 45178 11591 45180
rect 11615 45178 11671 45180
rect 11375 45126 11421 45178
rect 11421 45126 11431 45178
rect 11455 45126 11485 45178
rect 11485 45126 11497 45178
rect 11497 45126 11511 45178
rect 11535 45126 11549 45178
rect 11549 45126 11561 45178
rect 11561 45126 11591 45178
rect 11615 45126 11625 45178
rect 11625 45126 11671 45178
rect 11375 45124 11431 45126
rect 11455 45124 11511 45126
rect 11535 45124 11591 45126
rect 11615 45124 11671 45126
rect 11375 44090 11431 44092
rect 11455 44090 11511 44092
rect 11535 44090 11591 44092
rect 11615 44090 11671 44092
rect 11375 44038 11421 44090
rect 11421 44038 11431 44090
rect 11455 44038 11485 44090
rect 11485 44038 11497 44090
rect 11497 44038 11511 44090
rect 11535 44038 11549 44090
rect 11549 44038 11561 44090
rect 11561 44038 11591 44090
rect 11615 44038 11625 44090
rect 11625 44038 11671 44090
rect 11375 44036 11431 44038
rect 11455 44036 11511 44038
rect 11535 44036 11591 44038
rect 11615 44036 11671 44038
rect 7902 43546 7958 43548
rect 7982 43546 8038 43548
rect 8062 43546 8118 43548
rect 8142 43546 8198 43548
rect 7902 43494 7948 43546
rect 7948 43494 7958 43546
rect 7982 43494 8012 43546
rect 8012 43494 8024 43546
rect 8024 43494 8038 43546
rect 8062 43494 8076 43546
rect 8076 43494 8088 43546
rect 8088 43494 8118 43546
rect 8142 43494 8152 43546
rect 8152 43494 8198 43546
rect 7902 43492 7958 43494
rect 7982 43492 8038 43494
rect 8062 43492 8118 43494
rect 8142 43492 8198 43494
rect 11375 43002 11431 43004
rect 11455 43002 11511 43004
rect 11535 43002 11591 43004
rect 11615 43002 11671 43004
rect 11375 42950 11421 43002
rect 11421 42950 11431 43002
rect 11455 42950 11485 43002
rect 11485 42950 11497 43002
rect 11497 42950 11511 43002
rect 11535 42950 11549 43002
rect 11549 42950 11561 43002
rect 11561 42950 11591 43002
rect 11615 42950 11625 43002
rect 11625 42950 11671 43002
rect 11375 42948 11431 42950
rect 11455 42948 11511 42950
rect 11535 42948 11591 42950
rect 11615 42948 11671 42950
rect 7902 42458 7958 42460
rect 7982 42458 8038 42460
rect 8062 42458 8118 42460
rect 8142 42458 8198 42460
rect 7902 42406 7948 42458
rect 7948 42406 7958 42458
rect 7982 42406 8012 42458
rect 8012 42406 8024 42458
rect 8024 42406 8038 42458
rect 8062 42406 8076 42458
rect 8076 42406 8088 42458
rect 8088 42406 8118 42458
rect 8142 42406 8152 42458
rect 8152 42406 8198 42458
rect 7902 42404 7958 42406
rect 7982 42404 8038 42406
rect 8062 42404 8118 42406
rect 8142 42404 8198 42406
rect 11375 41914 11431 41916
rect 11455 41914 11511 41916
rect 11535 41914 11591 41916
rect 11615 41914 11671 41916
rect 11375 41862 11421 41914
rect 11421 41862 11431 41914
rect 11455 41862 11485 41914
rect 11485 41862 11497 41914
rect 11497 41862 11511 41914
rect 11535 41862 11549 41914
rect 11549 41862 11561 41914
rect 11561 41862 11591 41914
rect 11615 41862 11625 41914
rect 11625 41862 11671 41914
rect 11375 41860 11431 41862
rect 11455 41860 11511 41862
rect 11535 41860 11591 41862
rect 11615 41860 11671 41862
rect 7902 41370 7958 41372
rect 7982 41370 8038 41372
rect 8062 41370 8118 41372
rect 8142 41370 8198 41372
rect 7902 41318 7948 41370
rect 7948 41318 7958 41370
rect 7982 41318 8012 41370
rect 8012 41318 8024 41370
rect 8024 41318 8038 41370
rect 8062 41318 8076 41370
rect 8076 41318 8088 41370
rect 8088 41318 8118 41370
rect 8142 41318 8152 41370
rect 8152 41318 8198 41370
rect 7902 41316 7958 41318
rect 7982 41316 8038 41318
rect 8062 41316 8118 41318
rect 8142 41316 8198 41318
rect 11375 40826 11431 40828
rect 11455 40826 11511 40828
rect 11535 40826 11591 40828
rect 11615 40826 11671 40828
rect 11375 40774 11421 40826
rect 11421 40774 11431 40826
rect 11455 40774 11485 40826
rect 11485 40774 11497 40826
rect 11497 40774 11511 40826
rect 11535 40774 11549 40826
rect 11549 40774 11561 40826
rect 11561 40774 11591 40826
rect 11615 40774 11625 40826
rect 11625 40774 11671 40826
rect 11375 40772 11431 40774
rect 11455 40772 11511 40774
rect 11535 40772 11591 40774
rect 11615 40772 11671 40774
rect 7902 40282 7958 40284
rect 7982 40282 8038 40284
rect 8062 40282 8118 40284
rect 8142 40282 8198 40284
rect 7902 40230 7948 40282
rect 7948 40230 7958 40282
rect 7982 40230 8012 40282
rect 8012 40230 8024 40282
rect 8024 40230 8038 40282
rect 8062 40230 8076 40282
rect 8076 40230 8088 40282
rect 8088 40230 8118 40282
rect 8142 40230 8152 40282
rect 8152 40230 8198 40282
rect 7902 40228 7958 40230
rect 7982 40228 8038 40230
rect 8062 40228 8118 40230
rect 8142 40228 8198 40230
rect 11375 39738 11431 39740
rect 11455 39738 11511 39740
rect 11535 39738 11591 39740
rect 11615 39738 11671 39740
rect 11375 39686 11421 39738
rect 11421 39686 11431 39738
rect 11455 39686 11485 39738
rect 11485 39686 11497 39738
rect 11497 39686 11511 39738
rect 11535 39686 11549 39738
rect 11549 39686 11561 39738
rect 11561 39686 11591 39738
rect 11615 39686 11625 39738
rect 11625 39686 11671 39738
rect 11375 39684 11431 39686
rect 11455 39684 11511 39686
rect 11535 39684 11591 39686
rect 11615 39684 11671 39686
rect 7902 39194 7958 39196
rect 7982 39194 8038 39196
rect 8062 39194 8118 39196
rect 8142 39194 8198 39196
rect 7902 39142 7948 39194
rect 7948 39142 7958 39194
rect 7982 39142 8012 39194
rect 8012 39142 8024 39194
rect 8024 39142 8038 39194
rect 8062 39142 8076 39194
rect 8076 39142 8088 39194
rect 8088 39142 8118 39194
rect 8142 39142 8152 39194
rect 8152 39142 8198 39194
rect 7902 39140 7958 39142
rect 7982 39140 8038 39142
rect 8062 39140 8118 39142
rect 8142 39140 8198 39142
rect 11375 38650 11431 38652
rect 11455 38650 11511 38652
rect 11535 38650 11591 38652
rect 11615 38650 11671 38652
rect 11375 38598 11421 38650
rect 11421 38598 11431 38650
rect 11455 38598 11485 38650
rect 11485 38598 11497 38650
rect 11497 38598 11511 38650
rect 11535 38598 11549 38650
rect 11549 38598 11561 38650
rect 11561 38598 11591 38650
rect 11615 38598 11625 38650
rect 11625 38598 11671 38650
rect 11375 38596 11431 38598
rect 11455 38596 11511 38598
rect 11535 38596 11591 38598
rect 11615 38596 11671 38598
rect 7902 38106 7958 38108
rect 7982 38106 8038 38108
rect 8062 38106 8118 38108
rect 8142 38106 8198 38108
rect 7902 38054 7948 38106
rect 7948 38054 7958 38106
rect 7982 38054 8012 38106
rect 8012 38054 8024 38106
rect 8024 38054 8038 38106
rect 8062 38054 8076 38106
rect 8076 38054 8088 38106
rect 8088 38054 8118 38106
rect 8142 38054 8152 38106
rect 8152 38054 8198 38106
rect 7902 38052 7958 38054
rect 7982 38052 8038 38054
rect 8062 38052 8118 38054
rect 8142 38052 8198 38054
rect 11375 37562 11431 37564
rect 11455 37562 11511 37564
rect 11535 37562 11591 37564
rect 11615 37562 11671 37564
rect 11375 37510 11421 37562
rect 11421 37510 11431 37562
rect 11455 37510 11485 37562
rect 11485 37510 11497 37562
rect 11497 37510 11511 37562
rect 11535 37510 11549 37562
rect 11549 37510 11561 37562
rect 11561 37510 11591 37562
rect 11615 37510 11625 37562
rect 11625 37510 11671 37562
rect 11375 37508 11431 37510
rect 11455 37508 11511 37510
rect 11535 37508 11591 37510
rect 11615 37508 11671 37510
rect 7902 37018 7958 37020
rect 7982 37018 8038 37020
rect 8062 37018 8118 37020
rect 8142 37018 8198 37020
rect 7902 36966 7948 37018
rect 7948 36966 7958 37018
rect 7982 36966 8012 37018
rect 8012 36966 8024 37018
rect 8024 36966 8038 37018
rect 8062 36966 8076 37018
rect 8076 36966 8088 37018
rect 8088 36966 8118 37018
rect 8142 36966 8152 37018
rect 8152 36966 8198 37018
rect 7902 36964 7958 36966
rect 7982 36964 8038 36966
rect 8062 36964 8118 36966
rect 8142 36964 8198 36966
rect 11375 36474 11431 36476
rect 11455 36474 11511 36476
rect 11535 36474 11591 36476
rect 11615 36474 11671 36476
rect 11375 36422 11421 36474
rect 11421 36422 11431 36474
rect 11455 36422 11485 36474
rect 11485 36422 11497 36474
rect 11497 36422 11511 36474
rect 11535 36422 11549 36474
rect 11549 36422 11561 36474
rect 11561 36422 11591 36474
rect 11615 36422 11625 36474
rect 11625 36422 11671 36474
rect 11375 36420 11431 36422
rect 11455 36420 11511 36422
rect 11535 36420 11591 36422
rect 11615 36420 11671 36422
rect 7902 35930 7958 35932
rect 7982 35930 8038 35932
rect 8062 35930 8118 35932
rect 8142 35930 8198 35932
rect 7902 35878 7948 35930
rect 7948 35878 7958 35930
rect 7982 35878 8012 35930
rect 8012 35878 8024 35930
rect 8024 35878 8038 35930
rect 8062 35878 8076 35930
rect 8076 35878 8088 35930
rect 8088 35878 8118 35930
rect 8142 35878 8152 35930
rect 8152 35878 8198 35930
rect 7902 35876 7958 35878
rect 7982 35876 8038 35878
rect 8062 35876 8118 35878
rect 8142 35876 8198 35878
rect 14848 45722 14904 45724
rect 14928 45722 14984 45724
rect 15008 45722 15064 45724
rect 15088 45722 15144 45724
rect 14848 45670 14894 45722
rect 14894 45670 14904 45722
rect 14928 45670 14958 45722
rect 14958 45670 14970 45722
rect 14970 45670 14984 45722
rect 15008 45670 15022 45722
rect 15022 45670 15034 45722
rect 15034 45670 15064 45722
rect 15088 45670 15098 45722
rect 15098 45670 15144 45722
rect 14848 45668 14904 45670
rect 14928 45668 14984 45670
rect 15008 45668 15064 45670
rect 15088 45668 15144 45670
rect 18321 47354 18377 47356
rect 18401 47354 18457 47356
rect 18481 47354 18537 47356
rect 18561 47354 18617 47356
rect 18321 47302 18367 47354
rect 18367 47302 18377 47354
rect 18401 47302 18431 47354
rect 18431 47302 18443 47354
rect 18443 47302 18457 47354
rect 18481 47302 18495 47354
rect 18495 47302 18507 47354
rect 18507 47302 18537 47354
rect 18561 47302 18571 47354
rect 18571 47302 18617 47354
rect 18321 47300 18377 47302
rect 18401 47300 18457 47302
rect 18481 47300 18537 47302
rect 18561 47300 18617 47302
rect 18321 46266 18377 46268
rect 18401 46266 18457 46268
rect 18481 46266 18537 46268
rect 18561 46266 18617 46268
rect 18321 46214 18367 46266
rect 18367 46214 18377 46266
rect 18401 46214 18431 46266
rect 18431 46214 18443 46266
rect 18443 46214 18457 46266
rect 18481 46214 18495 46266
rect 18495 46214 18507 46266
rect 18507 46214 18537 46266
rect 18561 46214 18571 46266
rect 18571 46214 18617 46266
rect 18321 46212 18377 46214
rect 18401 46212 18457 46214
rect 18481 46212 18537 46214
rect 18561 46212 18617 46214
rect 21794 46810 21850 46812
rect 21874 46810 21930 46812
rect 21954 46810 22010 46812
rect 22034 46810 22090 46812
rect 21794 46758 21840 46810
rect 21840 46758 21850 46810
rect 21874 46758 21904 46810
rect 21904 46758 21916 46810
rect 21916 46758 21930 46810
rect 21954 46758 21968 46810
rect 21968 46758 21980 46810
rect 21980 46758 22010 46810
rect 22034 46758 22044 46810
rect 22044 46758 22090 46810
rect 21794 46756 21850 46758
rect 21874 46756 21930 46758
rect 21954 46756 22010 46758
rect 22034 46756 22090 46758
rect 14848 44634 14904 44636
rect 14928 44634 14984 44636
rect 15008 44634 15064 44636
rect 15088 44634 15144 44636
rect 14848 44582 14894 44634
rect 14894 44582 14904 44634
rect 14928 44582 14958 44634
rect 14958 44582 14970 44634
rect 14970 44582 14984 44634
rect 15008 44582 15022 44634
rect 15022 44582 15034 44634
rect 15034 44582 15064 44634
rect 15088 44582 15098 44634
rect 15098 44582 15144 44634
rect 14848 44580 14904 44582
rect 14928 44580 14984 44582
rect 15008 44580 15064 44582
rect 15088 44580 15144 44582
rect 11375 35386 11431 35388
rect 11455 35386 11511 35388
rect 11535 35386 11591 35388
rect 11615 35386 11671 35388
rect 11375 35334 11421 35386
rect 11421 35334 11431 35386
rect 11455 35334 11485 35386
rect 11485 35334 11497 35386
rect 11497 35334 11511 35386
rect 11535 35334 11549 35386
rect 11549 35334 11561 35386
rect 11561 35334 11591 35386
rect 11615 35334 11625 35386
rect 11625 35334 11671 35386
rect 11375 35332 11431 35334
rect 11455 35332 11511 35334
rect 11535 35332 11591 35334
rect 11615 35332 11671 35334
rect 7902 34842 7958 34844
rect 7982 34842 8038 34844
rect 8062 34842 8118 34844
rect 8142 34842 8198 34844
rect 7902 34790 7948 34842
rect 7948 34790 7958 34842
rect 7982 34790 8012 34842
rect 8012 34790 8024 34842
rect 8024 34790 8038 34842
rect 8062 34790 8076 34842
rect 8076 34790 8088 34842
rect 8088 34790 8118 34842
rect 8142 34790 8152 34842
rect 8152 34790 8198 34842
rect 7902 34788 7958 34790
rect 7982 34788 8038 34790
rect 8062 34788 8118 34790
rect 8142 34788 8198 34790
rect 4429 26682 4485 26684
rect 4509 26682 4565 26684
rect 4589 26682 4645 26684
rect 4669 26682 4725 26684
rect 4429 26630 4475 26682
rect 4475 26630 4485 26682
rect 4509 26630 4539 26682
rect 4539 26630 4551 26682
rect 4551 26630 4565 26682
rect 4589 26630 4603 26682
rect 4603 26630 4615 26682
rect 4615 26630 4645 26682
rect 4669 26630 4679 26682
rect 4679 26630 4725 26682
rect 4429 26628 4485 26630
rect 4509 26628 4565 26630
rect 4589 26628 4645 26630
rect 4669 26628 4725 26630
rect 4429 25594 4485 25596
rect 4509 25594 4565 25596
rect 4589 25594 4645 25596
rect 4669 25594 4725 25596
rect 4429 25542 4475 25594
rect 4475 25542 4485 25594
rect 4509 25542 4539 25594
rect 4539 25542 4551 25594
rect 4551 25542 4565 25594
rect 4589 25542 4603 25594
rect 4603 25542 4615 25594
rect 4615 25542 4645 25594
rect 4669 25542 4679 25594
rect 4679 25542 4725 25594
rect 4429 25540 4485 25542
rect 4509 25540 4565 25542
rect 4589 25540 4645 25542
rect 4669 25540 4725 25542
rect 4429 24506 4485 24508
rect 4509 24506 4565 24508
rect 4589 24506 4645 24508
rect 4669 24506 4725 24508
rect 4429 24454 4475 24506
rect 4475 24454 4485 24506
rect 4509 24454 4539 24506
rect 4539 24454 4551 24506
rect 4551 24454 4565 24506
rect 4589 24454 4603 24506
rect 4603 24454 4615 24506
rect 4615 24454 4645 24506
rect 4669 24454 4679 24506
rect 4679 24454 4725 24506
rect 4429 24452 4485 24454
rect 4509 24452 4565 24454
rect 4589 24452 4645 24454
rect 4669 24452 4725 24454
rect 4429 23418 4485 23420
rect 4509 23418 4565 23420
rect 4589 23418 4645 23420
rect 4669 23418 4725 23420
rect 4429 23366 4475 23418
rect 4475 23366 4485 23418
rect 4509 23366 4539 23418
rect 4539 23366 4551 23418
rect 4551 23366 4565 23418
rect 4589 23366 4603 23418
rect 4603 23366 4615 23418
rect 4615 23366 4645 23418
rect 4669 23366 4679 23418
rect 4679 23366 4725 23418
rect 4429 23364 4485 23366
rect 4509 23364 4565 23366
rect 4589 23364 4645 23366
rect 4669 23364 4725 23366
rect 4429 22330 4485 22332
rect 4509 22330 4565 22332
rect 4589 22330 4645 22332
rect 4669 22330 4725 22332
rect 4429 22278 4475 22330
rect 4475 22278 4485 22330
rect 4509 22278 4539 22330
rect 4539 22278 4551 22330
rect 4551 22278 4565 22330
rect 4589 22278 4603 22330
rect 4603 22278 4615 22330
rect 4615 22278 4645 22330
rect 4669 22278 4679 22330
rect 4679 22278 4725 22330
rect 4429 22276 4485 22278
rect 4509 22276 4565 22278
rect 4589 22276 4645 22278
rect 4669 22276 4725 22278
rect 4429 21242 4485 21244
rect 4509 21242 4565 21244
rect 4589 21242 4645 21244
rect 4669 21242 4725 21244
rect 4429 21190 4475 21242
rect 4475 21190 4485 21242
rect 4509 21190 4539 21242
rect 4539 21190 4551 21242
rect 4551 21190 4565 21242
rect 4589 21190 4603 21242
rect 4603 21190 4615 21242
rect 4615 21190 4645 21242
rect 4669 21190 4679 21242
rect 4679 21190 4725 21242
rect 4429 21188 4485 21190
rect 4509 21188 4565 21190
rect 4589 21188 4645 21190
rect 4669 21188 4725 21190
rect 4429 20154 4485 20156
rect 4509 20154 4565 20156
rect 4589 20154 4645 20156
rect 4669 20154 4725 20156
rect 4429 20102 4475 20154
rect 4475 20102 4485 20154
rect 4509 20102 4539 20154
rect 4539 20102 4551 20154
rect 4551 20102 4565 20154
rect 4589 20102 4603 20154
rect 4603 20102 4615 20154
rect 4615 20102 4645 20154
rect 4669 20102 4679 20154
rect 4679 20102 4725 20154
rect 4429 20100 4485 20102
rect 4509 20100 4565 20102
rect 4589 20100 4645 20102
rect 4669 20100 4725 20102
rect 4429 19066 4485 19068
rect 4509 19066 4565 19068
rect 4589 19066 4645 19068
rect 4669 19066 4725 19068
rect 4429 19014 4475 19066
rect 4475 19014 4485 19066
rect 4509 19014 4539 19066
rect 4539 19014 4551 19066
rect 4551 19014 4565 19066
rect 4589 19014 4603 19066
rect 4603 19014 4615 19066
rect 4615 19014 4645 19066
rect 4669 19014 4679 19066
rect 4679 19014 4725 19066
rect 4429 19012 4485 19014
rect 4509 19012 4565 19014
rect 4589 19012 4645 19014
rect 4669 19012 4725 19014
rect 4429 17978 4485 17980
rect 4509 17978 4565 17980
rect 4589 17978 4645 17980
rect 4669 17978 4725 17980
rect 4429 17926 4475 17978
rect 4475 17926 4485 17978
rect 4509 17926 4539 17978
rect 4539 17926 4551 17978
rect 4551 17926 4565 17978
rect 4589 17926 4603 17978
rect 4603 17926 4615 17978
rect 4615 17926 4645 17978
rect 4669 17926 4679 17978
rect 4679 17926 4725 17978
rect 4429 17924 4485 17926
rect 4509 17924 4565 17926
rect 4589 17924 4645 17926
rect 4669 17924 4725 17926
rect 7902 33754 7958 33756
rect 7982 33754 8038 33756
rect 8062 33754 8118 33756
rect 8142 33754 8198 33756
rect 7902 33702 7948 33754
rect 7948 33702 7958 33754
rect 7982 33702 8012 33754
rect 8012 33702 8024 33754
rect 8024 33702 8038 33754
rect 8062 33702 8076 33754
rect 8076 33702 8088 33754
rect 8088 33702 8118 33754
rect 8142 33702 8152 33754
rect 8152 33702 8198 33754
rect 7902 33700 7958 33702
rect 7982 33700 8038 33702
rect 8062 33700 8118 33702
rect 8142 33700 8198 33702
rect 7902 32666 7958 32668
rect 7982 32666 8038 32668
rect 8062 32666 8118 32668
rect 8142 32666 8198 32668
rect 7902 32614 7948 32666
rect 7948 32614 7958 32666
rect 7982 32614 8012 32666
rect 8012 32614 8024 32666
rect 8024 32614 8038 32666
rect 8062 32614 8076 32666
rect 8076 32614 8088 32666
rect 8088 32614 8118 32666
rect 8142 32614 8152 32666
rect 8152 32614 8198 32666
rect 7902 32612 7958 32614
rect 7982 32612 8038 32614
rect 8062 32612 8118 32614
rect 8142 32612 8198 32614
rect 7902 31578 7958 31580
rect 7982 31578 8038 31580
rect 8062 31578 8118 31580
rect 8142 31578 8198 31580
rect 7902 31526 7948 31578
rect 7948 31526 7958 31578
rect 7982 31526 8012 31578
rect 8012 31526 8024 31578
rect 8024 31526 8038 31578
rect 8062 31526 8076 31578
rect 8076 31526 8088 31578
rect 8088 31526 8118 31578
rect 8142 31526 8152 31578
rect 8152 31526 8198 31578
rect 7902 31524 7958 31526
rect 7982 31524 8038 31526
rect 8062 31524 8118 31526
rect 8142 31524 8198 31526
rect 7902 30490 7958 30492
rect 7982 30490 8038 30492
rect 8062 30490 8118 30492
rect 8142 30490 8198 30492
rect 7902 30438 7948 30490
rect 7948 30438 7958 30490
rect 7982 30438 8012 30490
rect 8012 30438 8024 30490
rect 8024 30438 8038 30490
rect 8062 30438 8076 30490
rect 8076 30438 8088 30490
rect 8088 30438 8118 30490
rect 8142 30438 8152 30490
rect 8152 30438 8198 30490
rect 7902 30436 7958 30438
rect 7982 30436 8038 30438
rect 8062 30436 8118 30438
rect 8142 30436 8198 30438
rect 7902 29402 7958 29404
rect 7982 29402 8038 29404
rect 8062 29402 8118 29404
rect 8142 29402 8198 29404
rect 7902 29350 7948 29402
rect 7948 29350 7958 29402
rect 7982 29350 8012 29402
rect 8012 29350 8024 29402
rect 8024 29350 8038 29402
rect 8062 29350 8076 29402
rect 8076 29350 8088 29402
rect 8088 29350 8118 29402
rect 8142 29350 8152 29402
rect 8152 29350 8198 29402
rect 7902 29348 7958 29350
rect 7982 29348 8038 29350
rect 8062 29348 8118 29350
rect 8142 29348 8198 29350
rect 7902 28314 7958 28316
rect 7982 28314 8038 28316
rect 8062 28314 8118 28316
rect 8142 28314 8198 28316
rect 7902 28262 7948 28314
rect 7948 28262 7958 28314
rect 7982 28262 8012 28314
rect 8012 28262 8024 28314
rect 8024 28262 8038 28314
rect 8062 28262 8076 28314
rect 8076 28262 8088 28314
rect 8088 28262 8118 28314
rect 8142 28262 8152 28314
rect 8152 28262 8198 28314
rect 7902 28260 7958 28262
rect 7982 28260 8038 28262
rect 8062 28260 8118 28262
rect 8142 28260 8198 28262
rect 7902 27226 7958 27228
rect 7982 27226 8038 27228
rect 8062 27226 8118 27228
rect 8142 27226 8198 27228
rect 7902 27174 7948 27226
rect 7948 27174 7958 27226
rect 7982 27174 8012 27226
rect 8012 27174 8024 27226
rect 8024 27174 8038 27226
rect 8062 27174 8076 27226
rect 8076 27174 8088 27226
rect 8088 27174 8118 27226
rect 8142 27174 8152 27226
rect 8152 27174 8198 27226
rect 7902 27172 7958 27174
rect 7982 27172 8038 27174
rect 8062 27172 8118 27174
rect 8142 27172 8198 27174
rect 7902 26138 7958 26140
rect 7982 26138 8038 26140
rect 8062 26138 8118 26140
rect 8142 26138 8198 26140
rect 7902 26086 7948 26138
rect 7948 26086 7958 26138
rect 7982 26086 8012 26138
rect 8012 26086 8024 26138
rect 8024 26086 8038 26138
rect 8062 26086 8076 26138
rect 8076 26086 8088 26138
rect 8088 26086 8118 26138
rect 8142 26086 8152 26138
rect 8152 26086 8198 26138
rect 7902 26084 7958 26086
rect 7982 26084 8038 26086
rect 8062 26084 8118 26086
rect 8142 26084 8198 26086
rect 7902 25050 7958 25052
rect 7982 25050 8038 25052
rect 8062 25050 8118 25052
rect 8142 25050 8198 25052
rect 7902 24998 7948 25050
rect 7948 24998 7958 25050
rect 7982 24998 8012 25050
rect 8012 24998 8024 25050
rect 8024 24998 8038 25050
rect 8062 24998 8076 25050
rect 8076 24998 8088 25050
rect 8088 24998 8118 25050
rect 8142 24998 8152 25050
rect 8152 24998 8198 25050
rect 7902 24996 7958 24998
rect 7982 24996 8038 24998
rect 8062 24996 8118 24998
rect 8142 24996 8198 24998
rect 7902 23962 7958 23964
rect 7982 23962 8038 23964
rect 8062 23962 8118 23964
rect 8142 23962 8198 23964
rect 7902 23910 7948 23962
rect 7948 23910 7958 23962
rect 7982 23910 8012 23962
rect 8012 23910 8024 23962
rect 8024 23910 8038 23962
rect 8062 23910 8076 23962
rect 8076 23910 8088 23962
rect 8088 23910 8118 23962
rect 8142 23910 8152 23962
rect 8152 23910 8198 23962
rect 7902 23908 7958 23910
rect 7982 23908 8038 23910
rect 8062 23908 8118 23910
rect 8142 23908 8198 23910
rect 7902 22874 7958 22876
rect 7982 22874 8038 22876
rect 8062 22874 8118 22876
rect 8142 22874 8198 22876
rect 7902 22822 7948 22874
rect 7948 22822 7958 22874
rect 7982 22822 8012 22874
rect 8012 22822 8024 22874
rect 8024 22822 8038 22874
rect 8062 22822 8076 22874
rect 8076 22822 8088 22874
rect 8088 22822 8118 22874
rect 8142 22822 8152 22874
rect 8152 22822 8198 22874
rect 7902 22820 7958 22822
rect 7982 22820 8038 22822
rect 8062 22820 8118 22822
rect 8142 22820 8198 22822
rect 7902 21786 7958 21788
rect 7982 21786 8038 21788
rect 8062 21786 8118 21788
rect 8142 21786 8198 21788
rect 7902 21734 7948 21786
rect 7948 21734 7958 21786
rect 7982 21734 8012 21786
rect 8012 21734 8024 21786
rect 8024 21734 8038 21786
rect 8062 21734 8076 21786
rect 8076 21734 8088 21786
rect 8088 21734 8118 21786
rect 8142 21734 8152 21786
rect 8152 21734 8198 21786
rect 7902 21732 7958 21734
rect 7982 21732 8038 21734
rect 8062 21732 8118 21734
rect 8142 21732 8198 21734
rect 7902 20698 7958 20700
rect 7982 20698 8038 20700
rect 8062 20698 8118 20700
rect 8142 20698 8198 20700
rect 7902 20646 7948 20698
rect 7948 20646 7958 20698
rect 7982 20646 8012 20698
rect 8012 20646 8024 20698
rect 8024 20646 8038 20698
rect 8062 20646 8076 20698
rect 8076 20646 8088 20698
rect 8088 20646 8118 20698
rect 8142 20646 8152 20698
rect 8152 20646 8198 20698
rect 7902 20644 7958 20646
rect 7982 20644 8038 20646
rect 8062 20644 8118 20646
rect 8142 20644 8198 20646
rect 7902 19610 7958 19612
rect 7982 19610 8038 19612
rect 8062 19610 8118 19612
rect 8142 19610 8198 19612
rect 7902 19558 7948 19610
rect 7948 19558 7958 19610
rect 7982 19558 8012 19610
rect 8012 19558 8024 19610
rect 8024 19558 8038 19610
rect 8062 19558 8076 19610
rect 8076 19558 8088 19610
rect 8088 19558 8118 19610
rect 8142 19558 8152 19610
rect 8152 19558 8198 19610
rect 7902 19556 7958 19558
rect 7982 19556 8038 19558
rect 8062 19556 8118 19558
rect 8142 19556 8198 19558
rect 7902 18522 7958 18524
rect 7982 18522 8038 18524
rect 8062 18522 8118 18524
rect 8142 18522 8198 18524
rect 7902 18470 7948 18522
rect 7948 18470 7958 18522
rect 7982 18470 8012 18522
rect 8012 18470 8024 18522
rect 8024 18470 8038 18522
rect 8062 18470 8076 18522
rect 8076 18470 8088 18522
rect 8088 18470 8118 18522
rect 8142 18470 8152 18522
rect 8152 18470 8198 18522
rect 7902 18468 7958 18470
rect 7982 18468 8038 18470
rect 8062 18468 8118 18470
rect 8142 18468 8198 18470
rect 7902 17434 7958 17436
rect 7982 17434 8038 17436
rect 8062 17434 8118 17436
rect 8142 17434 8198 17436
rect 7902 17382 7948 17434
rect 7948 17382 7958 17434
rect 7982 17382 8012 17434
rect 8012 17382 8024 17434
rect 8024 17382 8038 17434
rect 8062 17382 8076 17434
rect 8076 17382 8088 17434
rect 8088 17382 8118 17434
rect 8142 17382 8152 17434
rect 8152 17382 8198 17434
rect 7902 17380 7958 17382
rect 7982 17380 8038 17382
rect 8062 17380 8118 17382
rect 8142 17380 8198 17382
rect 4429 16890 4485 16892
rect 4509 16890 4565 16892
rect 4589 16890 4645 16892
rect 4669 16890 4725 16892
rect 4429 16838 4475 16890
rect 4475 16838 4485 16890
rect 4509 16838 4539 16890
rect 4539 16838 4551 16890
rect 4551 16838 4565 16890
rect 4589 16838 4603 16890
rect 4603 16838 4615 16890
rect 4615 16838 4645 16890
rect 4669 16838 4679 16890
rect 4679 16838 4725 16890
rect 4429 16836 4485 16838
rect 4509 16836 4565 16838
rect 4589 16836 4645 16838
rect 4669 16836 4725 16838
rect 4066 8200 4122 8256
rect 7902 16346 7958 16348
rect 7982 16346 8038 16348
rect 8062 16346 8118 16348
rect 8142 16346 8198 16348
rect 7902 16294 7948 16346
rect 7948 16294 7958 16346
rect 7982 16294 8012 16346
rect 8012 16294 8024 16346
rect 8024 16294 8038 16346
rect 8062 16294 8076 16346
rect 8076 16294 8088 16346
rect 8088 16294 8118 16346
rect 8142 16294 8152 16346
rect 8152 16294 8198 16346
rect 7902 16292 7958 16294
rect 7982 16292 8038 16294
rect 8062 16292 8118 16294
rect 8142 16292 8198 16294
rect 4429 15802 4485 15804
rect 4509 15802 4565 15804
rect 4589 15802 4645 15804
rect 4669 15802 4725 15804
rect 4429 15750 4475 15802
rect 4475 15750 4485 15802
rect 4509 15750 4539 15802
rect 4539 15750 4551 15802
rect 4551 15750 4565 15802
rect 4589 15750 4603 15802
rect 4603 15750 4615 15802
rect 4615 15750 4645 15802
rect 4669 15750 4679 15802
rect 4679 15750 4725 15802
rect 4429 15748 4485 15750
rect 4509 15748 4565 15750
rect 4589 15748 4645 15750
rect 4669 15748 4725 15750
rect 7902 15258 7958 15260
rect 7982 15258 8038 15260
rect 8062 15258 8118 15260
rect 8142 15258 8198 15260
rect 7902 15206 7948 15258
rect 7948 15206 7958 15258
rect 7982 15206 8012 15258
rect 8012 15206 8024 15258
rect 8024 15206 8038 15258
rect 8062 15206 8076 15258
rect 8076 15206 8088 15258
rect 8088 15206 8118 15258
rect 8142 15206 8152 15258
rect 8152 15206 8198 15258
rect 7902 15204 7958 15206
rect 7982 15204 8038 15206
rect 8062 15204 8118 15206
rect 8142 15204 8198 15206
rect 4429 14714 4485 14716
rect 4509 14714 4565 14716
rect 4589 14714 4645 14716
rect 4669 14714 4725 14716
rect 4429 14662 4475 14714
rect 4475 14662 4485 14714
rect 4509 14662 4539 14714
rect 4539 14662 4551 14714
rect 4551 14662 4565 14714
rect 4589 14662 4603 14714
rect 4603 14662 4615 14714
rect 4615 14662 4645 14714
rect 4669 14662 4679 14714
rect 4679 14662 4725 14714
rect 4429 14660 4485 14662
rect 4509 14660 4565 14662
rect 4589 14660 4645 14662
rect 4669 14660 4725 14662
rect 11375 34298 11431 34300
rect 11455 34298 11511 34300
rect 11535 34298 11591 34300
rect 11615 34298 11671 34300
rect 11375 34246 11421 34298
rect 11421 34246 11431 34298
rect 11455 34246 11485 34298
rect 11485 34246 11497 34298
rect 11497 34246 11511 34298
rect 11535 34246 11549 34298
rect 11549 34246 11561 34298
rect 11561 34246 11591 34298
rect 11615 34246 11625 34298
rect 11625 34246 11671 34298
rect 11375 34244 11431 34246
rect 11455 34244 11511 34246
rect 11535 34244 11591 34246
rect 11615 34244 11671 34246
rect 11375 33210 11431 33212
rect 11455 33210 11511 33212
rect 11535 33210 11591 33212
rect 11615 33210 11671 33212
rect 11375 33158 11421 33210
rect 11421 33158 11431 33210
rect 11455 33158 11485 33210
rect 11485 33158 11497 33210
rect 11497 33158 11511 33210
rect 11535 33158 11549 33210
rect 11549 33158 11561 33210
rect 11561 33158 11591 33210
rect 11615 33158 11625 33210
rect 11625 33158 11671 33210
rect 11375 33156 11431 33158
rect 11455 33156 11511 33158
rect 11535 33156 11591 33158
rect 11615 33156 11671 33158
rect 11375 32122 11431 32124
rect 11455 32122 11511 32124
rect 11535 32122 11591 32124
rect 11615 32122 11671 32124
rect 11375 32070 11421 32122
rect 11421 32070 11431 32122
rect 11455 32070 11485 32122
rect 11485 32070 11497 32122
rect 11497 32070 11511 32122
rect 11535 32070 11549 32122
rect 11549 32070 11561 32122
rect 11561 32070 11591 32122
rect 11615 32070 11625 32122
rect 11625 32070 11671 32122
rect 11375 32068 11431 32070
rect 11455 32068 11511 32070
rect 11535 32068 11591 32070
rect 11615 32068 11671 32070
rect 11375 31034 11431 31036
rect 11455 31034 11511 31036
rect 11535 31034 11591 31036
rect 11615 31034 11671 31036
rect 11375 30982 11421 31034
rect 11421 30982 11431 31034
rect 11455 30982 11485 31034
rect 11485 30982 11497 31034
rect 11497 30982 11511 31034
rect 11535 30982 11549 31034
rect 11549 30982 11561 31034
rect 11561 30982 11591 31034
rect 11615 30982 11625 31034
rect 11625 30982 11671 31034
rect 11375 30980 11431 30982
rect 11455 30980 11511 30982
rect 11535 30980 11591 30982
rect 11615 30980 11671 30982
rect 11375 29946 11431 29948
rect 11455 29946 11511 29948
rect 11535 29946 11591 29948
rect 11615 29946 11671 29948
rect 11375 29894 11421 29946
rect 11421 29894 11431 29946
rect 11455 29894 11485 29946
rect 11485 29894 11497 29946
rect 11497 29894 11511 29946
rect 11535 29894 11549 29946
rect 11549 29894 11561 29946
rect 11561 29894 11591 29946
rect 11615 29894 11625 29946
rect 11625 29894 11671 29946
rect 11375 29892 11431 29894
rect 11455 29892 11511 29894
rect 11535 29892 11591 29894
rect 11615 29892 11671 29894
rect 11375 28858 11431 28860
rect 11455 28858 11511 28860
rect 11535 28858 11591 28860
rect 11615 28858 11671 28860
rect 11375 28806 11421 28858
rect 11421 28806 11431 28858
rect 11455 28806 11485 28858
rect 11485 28806 11497 28858
rect 11497 28806 11511 28858
rect 11535 28806 11549 28858
rect 11549 28806 11561 28858
rect 11561 28806 11591 28858
rect 11615 28806 11625 28858
rect 11625 28806 11671 28858
rect 11375 28804 11431 28806
rect 11455 28804 11511 28806
rect 11535 28804 11591 28806
rect 11615 28804 11671 28806
rect 11375 27770 11431 27772
rect 11455 27770 11511 27772
rect 11535 27770 11591 27772
rect 11615 27770 11671 27772
rect 11375 27718 11421 27770
rect 11421 27718 11431 27770
rect 11455 27718 11485 27770
rect 11485 27718 11497 27770
rect 11497 27718 11511 27770
rect 11535 27718 11549 27770
rect 11549 27718 11561 27770
rect 11561 27718 11591 27770
rect 11615 27718 11625 27770
rect 11625 27718 11671 27770
rect 11375 27716 11431 27718
rect 11455 27716 11511 27718
rect 11535 27716 11591 27718
rect 11615 27716 11671 27718
rect 11375 26682 11431 26684
rect 11455 26682 11511 26684
rect 11535 26682 11591 26684
rect 11615 26682 11671 26684
rect 11375 26630 11421 26682
rect 11421 26630 11431 26682
rect 11455 26630 11485 26682
rect 11485 26630 11497 26682
rect 11497 26630 11511 26682
rect 11535 26630 11549 26682
rect 11549 26630 11561 26682
rect 11561 26630 11591 26682
rect 11615 26630 11625 26682
rect 11625 26630 11671 26682
rect 11375 26628 11431 26630
rect 11455 26628 11511 26630
rect 11535 26628 11591 26630
rect 11615 26628 11671 26630
rect 11375 25594 11431 25596
rect 11455 25594 11511 25596
rect 11535 25594 11591 25596
rect 11615 25594 11671 25596
rect 11375 25542 11421 25594
rect 11421 25542 11431 25594
rect 11455 25542 11485 25594
rect 11485 25542 11497 25594
rect 11497 25542 11511 25594
rect 11535 25542 11549 25594
rect 11549 25542 11561 25594
rect 11561 25542 11591 25594
rect 11615 25542 11625 25594
rect 11625 25542 11671 25594
rect 11375 25540 11431 25542
rect 11455 25540 11511 25542
rect 11535 25540 11591 25542
rect 11615 25540 11671 25542
rect 7902 14170 7958 14172
rect 7982 14170 8038 14172
rect 8062 14170 8118 14172
rect 8142 14170 8198 14172
rect 7902 14118 7948 14170
rect 7948 14118 7958 14170
rect 7982 14118 8012 14170
rect 8012 14118 8024 14170
rect 8024 14118 8038 14170
rect 8062 14118 8076 14170
rect 8076 14118 8088 14170
rect 8088 14118 8118 14170
rect 8142 14118 8152 14170
rect 8152 14118 8198 14170
rect 7902 14116 7958 14118
rect 7982 14116 8038 14118
rect 8062 14116 8118 14118
rect 8142 14116 8198 14118
rect 4429 13626 4485 13628
rect 4509 13626 4565 13628
rect 4589 13626 4645 13628
rect 4669 13626 4725 13628
rect 4429 13574 4475 13626
rect 4475 13574 4485 13626
rect 4509 13574 4539 13626
rect 4539 13574 4551 13626
rect 4551 13574 4565 13626
rect 4589 13574 4603 13626
rect 4603 13574 4615 13626
rect 4615 13574 4645 13626
rect 4669 13574 4679 13626
rect 4679 13574 4725 13626
rect 4429 13572 4485 13574
rect 4509 13572 4565 13574
rect 4589 13572 4645 13574
rect 4669 13572 4725 13574
rect 7902 13082 7958 13084
rect 7982 13082 8038 13084
rect 8062 13082 8118 13084
rect 8142 13082 8198 13084
rect 7902 13030 7948 13082
rect 7948 13030 7958 13082
rect 7982 13030 8012 13082
rect 8012 13030 8024 13082
rect 8024 13030 8038 13082
rect 8062 13030 8076 13082
rect 8076 13030 8088 13082
rect 8088 13030 8118 13082
rect 8142 13030 8152 13082
rect 8152 13030 8198 13082
rect 7902 13028 7958 13030
rect 7982 13028 8038 13030
rect 8062 13028 8118 13030
rect 8142 13028 8198 13030
rect 4429 12538 4485 12540
rect 4509 12538 4565 12540
rect 4589 12538 4645 12540
rect 4669 12538 4725 12540
rect 4429 12486 4475 12538
rect 4475 12486 4485 12538
rect 4509 12486 4539 12538
rect 4539 12486 4551 12538
rect 4551 12486 4565 12538
rect 4589 12486 4603 12538
rect 4603 12486 4615 12538
rect 4615 12486 4645 12538
rect 4669 12486 4679 12538
rect 4679 12486 4725 12538
rect 4429 12484 4485 12486
rect 4509 12484 4565 12486
rect 4589 12484 4645 12486
rect 4669 12484 4725 12486
rect 7902 11994 7958 11996
rect 7982 11994 8038 11996
rect 8062 11994 8118 11996
rect 8142 11994 8198 11996
rect 7902 11942 7948 11994
rect 7948 11942 7958 11994
rect 7982 11942 8012 11994
rect 8012 11942 8024 11994
rect 8024 11942 8038 11994
rect 8062 11942 8076 11994
rect 8076 11942 8088 11994
rect 8088 11942 8118 11994
rect 8142 11942 8152 11994
rect 8152 11942 8198 11994
rect 7902 11940 7958 11942
rect 7982 11940 8038 11942
rect 8062 11940 8118 11942
rect 8142 11940 8198 11942
rect 4429 11450 4485 11452
rect 4509 11450 4565 11452
rect 4589 11450 4645 11452
rect 4669 11450 4725 11452
rect 4429 11398 4475 11450
rect 4475 11398 4485 11450
rect 4509 11398 4539 11450
rect 4539 11398 4551 11450
rect 4551 11398 4565 11450
rect 4589 11398 4603 11450
rect 4603 11398 4615 11450
rect 4615 11398 4645 11450
rect 4669 11398 4679 11450
rect 4679 11398 4725 11450
rect 4429 11396 4485 11398
rect 4509 11396 4565 11398
rect 4589 11396 4645 11398
rect 4669 11396 4725 11398
rect 7902 10906 7958 10908
rect 7982 10906 8038 10908
rect 8062 10906 8118 10908
rect 8142 10906 8198 10908
rect 7902 10854 7948 10906
rect 7948 10854 7958 10906
rect 7982 10854 8012 10906
rect 8012 10854 8024 10906
rect 8024 10854 8038 10906
rect 8062 10854 8076 10906
rect 8076 10854 8088 10906
rect 8088 10854 8118 10906
rect 8142 10854 8152 10906
rect 8152 10854 8198 10906
rect 7902 10852 7958 10854
rect 7982 10852 8038 10854
rect 8062 10852 8118 10854
rect 8142 10852 8198 10854
rect 4429 10362 4485 10364
rect 4509 10362 4565 10364
rect 4589 10362 4645 10364
rect 4669 10362 4725 10364
rect 4429 10310 4475 10362
rect 4475 10310 4485 10362
rect 4509 10310 4539 10362
rect 4539 10310 4551 10362
rect 4551 10310 4565 10362
rect 4589 10310 4603 10362
rect 4603 10310 4615 10362
rect 4615 10310 4645 10362
rect 4669 10310 4679 10362
rect 4679 10310 4725 10362
rect 4429 10308 4485 10310
rect 4509 10308 4565 10310
rect 4589 10308 4645 10310
rect 4669 10308 4725 10310
rect 7902 9818 7958 9820
rect 7982 9818 8038 9820
rect 8062 9818 8118 9820
rect 8142 9818 8198 9820
rect 7902 9766 7948 9818
rect 7948 9766 7958 9818
rect 7982 9766 8012 9818
rect 8012 9766 8024 9818
rect 8024 9766 8038 9818
rect 8062 9766 8076 9818
rect 8076 9766 8088 9818
rect 8088 9766 8118 9818
rect 8142 9766 8152 9818
rect 8152 9766 8198 9818
rect 7902 9764 7958 9766
rect 7982 9764 8038 9766
rect 8062 9764 8118 9766
rect 8142 9764 8198 9766
rect 4429 9274 4485 9276
rect 4509 9274 4565 9276
rect 4589 9274 4645 9276
rect 4669 9274 4725 9276
rect 4429 9222 4475 9274
rect 4475 9222 4485 9274
rect 4509 9222 4539 9274
rect 4539 9222 4551 9274
rect 4551 9222 4565 9274
rect 4589 9222 4603 9274
rect 4603 9222 4615 9274
rect 4615 9222 4645 9274
rect 4669 9222 4679 9274
rect 4679 9222 4725 9274
rect 4429 9220 4485 9222
rect 4509 9220 4565 9222
rect 4589 9220 4645 9222
rect 4669 9220 4725 9222
rect 7902 8730 7958 8732
rect 7982 8730 8038 8732
rect 8062 8730 8118 8732
rect 8142 8730 8198 8732
rect 7902 8678 7948 8730
rect 7948 8678 7958 8730
rect 7982 8678 8012 8730
rect 8012 8678 8024 8730
rect 8024 8678 8038 8730
rect 8062 8678 8076 8730
rect 8076 8678 8088 8730
rect 8088 8678 8118 8730
rect 8142 8678 8152 8730
rect 8152 8678 8198 8730
rect 7902 8676 7958 8678
rect 7982 8676 8038 8678
rect 8062 8676 8118 8678
rect 8142 8676 8198 8678
rect 4429 8186 4485 8188
rect 4509 8186 4565 8188
rect 4589 8186 4645 8188
rect 4669 8186 4725 8188
rect 4429 8134 4475 8186
rect 4475 8134 4485 8186
rect 4509 8134 4539 8186
rect 4539 8134 4551 8186
rect 4551 8134 4565 8186
rect 4589 8134 4603 8186
rect 4603 8134 4615 8186
rect 4615 8134 4645 8186
rect 4669 8134 4679 8186
rect 4679 8134 4725 8186
rect 4429 8132 4485 8134
rect 4509 8132 4565 8134
rect 4589 8132 4645 8134
rect 4669 8132 4725 8134
rect 4429 7098 4485 7100
rect 4509 7098 4565 7100
rect 4589 7098 4645 7100
rect 4669 7098 4725 7100
rect 4429 7046 4475 7098
rect 4475 7046 4485 7098
rect 4509 7046 4539 7098
rect 4539 7046 4551 7098
rect 4551 7046 4565 7098
rect 4589 7046 4603 7098
rect 4603 7046 4615 7098
rect 4615 7046 4645 7098
rect 4669 7046 4679 7098
rect 4679 7046 4725 7098
rect 4429 7044 4485 7046
rect 4509 7044 4565 7046
rect 4589 7044 4645 7046
rect 4669 7044 4725 7046
rect 3606 6160 3662 6216
rect 2778 4800 2834 4856
rect 4066 4120 4122 4176
rect 3054 3440 3110 3496
rect 2870 2760 2926 2816
rect 2778 1400 2834 1456
rect 3514 2080 3570 2136
rect 4429 6010 4485 6012
rect 4509 6010 4565 6012
rect 4589 6010 4645 6012
rect 4669 6010 4725 6012
rect 4429 5958 4475 6010
rect 4475 5958 4485 6010
rect 4509 5958 4539 6010
rect 4539 5958 4551 6010
rect 4551 5958 4565 6010
rect 4589 5958 4603 6010
rect 4603 5958 4615 6010
rect 4615 5958 4645 6010
rect 4669 5958 4679 6010
rect 4679 5958 4725 6010
rect 4429 5956 4485 5958
rect 4509 5956 4565 5958
rect 4589 5956 4645 5958
rect 4669 5956 4725 5958
rect 4429 4922 4485 4924
rect 4509 4922 4565 4924
rect 4589 4922 4645 4924
rect 4669 4922 4725 4924
rect 4429 4870 4475 4922
rect 4475 4870 4485 4922
rect 4509 4870 4539 4922
rect 4539 4870 4551 4922
rect 4551 4870 4565 4922
rect 4589 4870 4603 4922
rect 4603 4870 4615 4922
rect 4615 4870 4645 4922
rect 4669 4870 4679 4922
rect 4679 4870 4725 4922
rect 4429 4868 4485 4870
rect 4509 4868 4565 4870
rect 4589 4868 4645 4870
rect 4669 4868 4725 4870
rect 4429 3834 4485 3836
rect 4509 3834 4565 3836
rect 4589 3834 4645 3836
rect 4669 3834 4725 3836
rect 4429 3782 4475 3834
rect 4475 3782 4485 3834
rect 4509 3782 4539 3834
rect 4539 3782 4551 3834
rect 4551 3782 4565 3834
rect 4589 3782 4603 3834
rect 4603 3782 4615 3834
rect 4615 3782 4645 3834
rect 4669 3782 4679 3834
rect 4679 3782 4725 3834
rect 4429 3780 4485 3782
rect 4509 3780 4565 3782
rect 4589 3780 4645 3782
rect 4669 3780 4725 3782
rect 7902 7642 7958 7644
rect 7982 7642 8038 7644
rect 8062 7642 8118 7644
rect 8142 7642 8198 7644
rect 7902 7590 7948 7642
rect 7948 7590 7958 7642
rect 7982 7590 8012 7642
rect 8012 7590 8024 7642
rect 8024 7590 8038 7642
rect 8062 7590 8076 7642
rect 8076 7590 8088 7642
rect 8088 7590 8118 7642
rect 8142 7590 8152 7642
rect 8152 7590 8198 7642
rect 7902 7588 7958 7590
rect 7982 7588 8038 7590
rect 8062 7588 8118 7590
rect 8142 7588 8198 7590
rect 7902 6554 7958 6556
rect 7982 6554 8038 6556
rect 8062 6554 8118 6556
rect 8142 6554 8198 6556
rect 7902 6502 7948 6554
rect 7948 6502 7958 6554
rect 7982 6502 8012 6554
rect 8012 6502 8024 6554
rect 8024 6502 8038 6554
rect 8062 6502 8076 6554
rect 8076 6502 8088 6554
rect 8088 6502 8118 6554
rect 8142 6502 8152 6554
rect 8152 6502 8198 6554
rect 7902 6500 7958 6502
rect 7982 6500 8038 6502
rect 8062 6500 8118 6502
rect 8142 6500 8198 6502
rect 7902 5466 7958 5468
rect 7982 5466 8038 5468
rect 8062 5466 8118 5468
rect 8142 5466 8198 5468
rect 7902 5414 7948 5466
rect 7948 5414 7958 5466
rect 7982 5414 8012 5466
rect 8012 5414 8024 5466
rect 8024 5414 8038 5466
rect 8062 5414 8076 5466
rect 8076 5414 8088 5466
rect 8088 5414 8118 5466
rect 8142 5414 8152 5466
rect 8152 5414 8198 5466
rect 7902 5412 7958 5414
rect 7982 5412 8038 5414
rect 8062 5412 8118 5414
rect 8142 5412 8198 5414
rect 4429 2746 4485 2748
rect 4509 2746 4565 2748
rect 4589 2746 4645 2748
rect 4669 2746 4725 2748
rect 4429 2694 4475 2746
rect 4475 2694 4485 2746
rect 4509 2694 4539 2746
rect 4539 2694 4551 2746
rect 4551 2694 4565 2746
rect 4589 2694 4603 2746
rect 4603 2694 4615 2746
rect 4615 2694 4645 2746
rect 4669 2694 4679 2746
rect 4679 2694 4725 2746
rect 4429 2692 4485 2694
rect 4509 2692 4565 2694
rect 4589 2692 4645 2694
rect 4669 2692 4725 2694
rect 7902 4378 7958 4380
rect 7982 4378 8038 4380
rect 8062 4378 8118 4380
rect 8142 4378 8198 4380
rect 7902 4326 7948 4378
rect 7948 4326 7958 4378
rect 7982 4326 8012 4378
rect 8012 4326 8024 4378
rect 8024 4326 8038 4378
rect 8062 4326 8076 4378
rect 8076 4326 8088 4378
rect 8088 4326 8118 4378
rect 8142 4326 8152 4378
rect 8152 4326 8198 4378
rect 7902 4324 7958 4326
rect 7982 4324 8038 4326
rect 8062 4324 8118 4326
rect 8142 4324 8198 4326
rect 7902 3290 7958 3292
rect 7982 3290 8038 3292
rect 8062 3290 8118 3292
rect 8142 3290 8198 3292
rect 7902 3238 7948 3290
rect 7948 3238 7958 3290
rect 7982 3238 8012 3290
rect 8012 3238 8024 3290
rect 8024 3238 8038 3290
rect 8062 3238 8076 3290
rect 8076 3238 8088 3290
rect 8088 3238 8118 3290
rect 8142 3238 8152 3290
rect 8152 3238 8198 3290
rect 7902 3236 7958 3238
rect 7982 3236 8038 3238
rect 8062 3236 8118 3238
rect 8142 3236 8198 3238
rect 7902 2202 7958 2204
rect 7982 2202 8038 2204
rect 8062 2202 8118 2204
rect 8142 2202 8198 2204
rect 7902 2150 7948 2202
rect 7948 2150 7958 2202
rect 7982 2150 8012 2202
rect 8012 2150 8024 2202
rect 8024 2150 8038 2202
rect 8062 2150 8076 2202
rect 8076 2150 8088 2202
rect 8088 2150 8118 2202
rect 8142 2150 8152 2202
rect 8152 2150 8198 2202
rect 7902 2148 7958 2150
rect 7982 2148 8038 2150
rect 8062 2148 8118 2150
rect 8142 2148 8198 2150
rect 11375 24506 11431 24508
rect 11455 24506 11511 24508
rect 11535 24506 11591 24508
rect 11615 24506 11671 24508
rect 11375 24454 11421 24506
rect 11421 24454 11431 24506
rect 11455 24454 11485 24506
rect 11485 24454 11497 24506
rect 11497 24454 11511 24506
rect 11535 24454 11549 24506
rect 11549 24454 11561 24506
rect 11561 24454 11591 24506
rect 11615 24454 11625 24506
rect 11625 24454 11671 24506
rect 11375 24452 11431 24454
rect 11455 24452 11511 24454
rect 11535 24452 11591 24454
rect 11615 24452 11671 24454
rect 11375 23418 11431 23420
rect 11455 23418 11511 23420
rect 11535 23418 11591 23420
rect 11615 23418 11671 23420
rect 11375 23366 11421 23418
rect 11421 23366 11431 23418
rect 11455 23366 11485 23418
rect 11485 23366 11497 23418
rect 11497 23366 11511 23418
rect 11535 23366 11549 23418
rect 11549 23366 11561 23418
rect 11561 23366 11591 23418
rect 11615 23366 11625 23418
rect 11625 23366 11671 23418
rect 11375 23364 11431 23366
rect 11455 23364 11511 23366
rect 11535 23364 11591 23366
rect 11615 23364 11671 23366
rect 11375 22330 11431 22332
rect 11455 22330 11511 22332
rect 11535 22330 11591 22332
rect 11615 22330 11671 22332
rect 11375 22278 11421 22330
rect 11421 22278 11431 22330
rect 11455 22278 11485 22330
rect 11485 22278 11497 22330
rect 11497 22278 11511 22330
rect 11535 22278 11549 22330
rect 11549 22278 11561 22330
rect 11561 22278 11591 22330
rect 11615 22278 11625 22330
rect 11625 22278 11671 22330
rect 11375 22276 11431 22278
rect 11455 22276 11511 22278
rect 11535 22276 11591 22278
rect 11615 22276 11671 22278
rect 11375 21242 11431 21244
rect 11455 21242 11511 21244
rect 11535 21242 11591 21244
rect 11615 21242 11671 21244
rect 11375 21190 11421 21242
rect 11421 21190 11431 21242
rect 11455 21190 11485 21242
rect 11485 21190 11497 21242
rect 11497 21190 11511 21242
rect 11535 21190 11549 21242
rect 11549 21190 11561 21242
rect 11561 21190 11591 21242
rect 11615 21190 11625 21242
rect 11625 21190 11671 21242
rect 11375 21188 11431 21190
rect 11455 21188 11511 21190
rect 11535 21188 11591 21190
rect 11615 21188 11671 21190
rect 11375 20154 11431 20156
rect 11455 20154 11511 20156
rect 11535 20154 11591 20156
rect 11615 20154 11671 20156
rect 11375 20102 11421 20154
rect 11421 20102 11431 20154
rect 11455 20102 11485 20154
rect 11485 20102 11497 20154
rect 11497 20102 11511 20154
rect 11535 20102 11549 20154
rect 11549 20102 11561 20154
rect 11561 20102 11591 20154
rect 11615 20102 11625 20154
rect 11625 20102 11671 20154
rect 11375 20100 11431 20102
rect 11455 20100 11511 20102
rect 11535 20100 11591 20102
rect 11615 20100 11671 20102
rect 11375 19066 11431 19068
rect 11455 19066 11511 19068
rect 11535 19066 11591 19068
rect 11615 19066 11671 19068
rect 11375 19014 11421 19066
rect 11421 19014 11431 19066
rect 11455 19014 11485 19066
rect 11485 19014 11497 19066
rect 11497 19014 11511 19066
rect 11535 19014 11549 19066
rect 11549 19014 11561 19066
rect 11561 19014 11591 19066
rect 11615 19014 11625 19066
rect 11625 19014 11671 19066
rect 11375 19012 11431 19014
rect 11455 19012 11511 19014
rect 11535 19012 11591 19014
rect 11615 19012 11671 19014
rect 11375 17978 11431 17980
rect 11455 17978 11511 17980
rect 11535 17978 11591 17980
rect 11615 17978 11671 17980
rect 11375 17926 11421 17978
rect 11421 17926 11431 17978
rect 11455 17926 11485 17978
rect 11485 17926 11497 17978
rect 11497 17926 11511 17978
rect 11535 17926 11549 17978
rect 11549 17926 11561 17978
rect 11561 17926 11591 17978
rect 11615 17926 11625 17978
rect 11625 17926 11671 17978
rect 11375 17924 11431 17926
rect 11455 17924 11511 17926
rect 11535 17924 11591 17926
rect 11615 17924 11671 17926
rect 11375 16890 11431 16892
rect 11455 16890 11511 16892
rect 11535 16890 11591 16892
rect 11615 16890 11671 16892
rect 11375 16838 11421 16890
rect 11421 16838 11431 16890
rect 11455 16838 11485 16890
rect 11485 16838 11497 16890
rect 11497 16838 11511 16890
rect 11535 16838 11549 16890
rect 11549 16838 11561 16890
rect 11561 16838 11591 16890
rect 11615 16838 11625 16890
rect 11625 16838 11671 16890
rect 11375 16836 11431 16838
rect 11455 16836 11511 16838
rect 11535 16836 11591 16838
rect 11615 16836 11671 16838
rect 11375 15802 11431 15804
rect 11455 15802 11511 15804
rect 11535 15802 11591 15804
rect 11615 15802 11671 15804
rect 11375 15750 11421 15802
rect 11421 15750 11431 15802
rect 11455 15750 11485 15802
rect 11485 15750 11497 15802
rect 11497 15750 11511 15802
rect 11535 15750 11549 15802
rect 11549 15750 11561 15802
rect 11561 15750 11591 15802
rect 11615 15750 11625 15802
rect 11625 15750 11671 15802
rect 11375 15748 11431 15750
rect 11455 15748 11511 15750
rect 11535 15748 11591 15750
rect 11615 15748 11671 15750
rect 11375 14714 11431 14716
rect 11455 14714 11511 14716
rect 11535 14714 11591 14716
rect 11615 14714 11671 14716
rect 11375 14662 11421 14714
rect 11421 14662 11431 14714
rect 11455 14662 11485 14714
rect 11485 14662 11497 14714
rect 11497 14662 11511 14714
rect 11535 14662 11549 14714
rect 11549 14662 11561 14714
rect 11561 14662 11591 14714
rect 11615 14662 11625 14714
rect 11625 14662 11671 14714
rect 11375 14660 11431 14662
rect 11455 14660 11511 14662
rect 11535 14660 11591 14662
rect 11615 14660 11671 14662
rect 11375 13626 11431 13628
rect 11455 13626 11511 13628
rect 11535 13626 11591 13628
rect 11615 13626 11671 13628
rect 11375 13574 11421 13626
rect 11421 13574 11431 13626
rect 11455 13574 11485 13626
rect 11485 13574 11497 13626
rect 11497 13574 11511 13626
rect 11535 13574 11549 13626
rect 11549 13574 11561 13626
rect 11561 13574 11591 13626
rect 11615 13574 11625 13626
rect 11625 13574 11671 13626
rect 11375 13572 11431 13574
rect 11455 13572 11511 13574
rect 11535 13572 11591 13574
rect 11615 13572 11671 13574
rect 11375 12538 11431 12540
rect 11455 12538 11511 12540
rect 11535 12538 11591 12540
rect 11615 12538 11671 12540
rect 11375 12486 11421 12538
rect 11421 12486 11431 12538
rect 11455 12486 11485 12538
rect 11485 12486 11497 12538
rect 11497 12486 11511 12538
rect 11535 12486 11549 12538
rect 11549 12486 11561 12538
rect 11561 12486 11591 12538
rect 11615 12486 11625 12538
rect 11625 12486 11671 12538
rect 11375 12484 11431 12486
rect 11455 12484 11511 12486
rect 11535 12484 11591 12486
rect 11615 12484 11671 12486
rect 11375 11450 11431 11452
rect 11455 11450 11511 11452
rect 11535 11450 11591 11452
rect 11615 11450 11671 11452
rect 11375 11398 11421 11450
rect 11421 11398 11431 11450
rect 11455 11398 11485 11450
rect 11485 11398 11497 11450
rect 11497 11398 11511 11450
rect 11535 11398 11549 11450
rect 11549 11398 11561 11450
rect 11561 11398 11591 11450
rect 11615 11398 11625 11450
rect 11625 11398 11671 11450
rect 11375 11396 11431 11398
rect 11455 11396 11511 11398
rect 11535 11396 11591 11398
rect 11615 11396 11671 11398
rect 11375 10362 11431 10364
rect 11455 10362 11511 10364
rect 11535 10362 11591 10364
rect 11615 10362 11671 10364
rect 11375 10310 11421 10362
rect 11421 10310 11431 10362
rect 11455 10310 11485 10362
rect 11485 10310 11497 10362
rect 11497 10310 11511 10362
rect 11535 10310 11549 10362
rect 11549 10310 11561 10362
rect 11561 10310 11591 10362
rect 11615 10310 11625 10362
rect 11625 10310 11671 10362
rect 11375 10308 11431 10310
rect 11455 10308 11511 10310
rect 11535 10308 11591 10310
rect 11615 10308 11671 10310
rect 11375 9274 11431 9276
rect 11455 9274 11511 9276
rect 11535 9274 11591 9276
rect 11615 9274 11671 9276
rect 11375 9222 11421 9274
rect 11421 9222 11431 9274
rect 11455 9222 11485 9274
rect 11485 9222 11497 9274
rect 11497 9222 11511 9274
rect 11535 9222 11549 9274
rect 11549 9222 11561 9274
rect 11561 9222 11591 9274
rect 11615 9222 11625 9274
rect 11625 9222 11671 9274
rect 11375 9220 11431 9222
rect 11455 9220 11511 9222
rect 11535 9220 11591 9222
rect 11615 9220 11671 9222
rect 14848 43546 14904 43548
rect 14928 43546 14984 43548
rect 15008 43546 15064 43548
rect 15088 43546 15144 43548
rect 14848 43494 14894 43546
rect 14894 43494 14904 43546
rect 14928 43494 14958 43546
rect 14958 43494 14970 43546
rect 14970 43494 14984 43546
rect 15008 43494 15022 43546
rect 15022 43494 15034 43546
rect 15034 43494 15064 43546
rect 15088 43494 15098 43546
rect 15098 43494 15144 43546
rect 14848 43492 14904 43494
rect 14928 43492 14984 43494
rect 15008 43492 15064 43494
rect 15088 43492 15144 43494
rect 18321 45178 18377 45180
rect 18401 45178 18457 45180
rect 18481 45178 18537 45180
rect 18561 45178 18617 45180
rect 18321 45126 18367 45178
rect 18367 45126 18377 45178
rect 18401 45126 18431 45178
rect 18431 45126 18443 45178
rect 18443 45126 18457 45178
rect 18481 45126 18495 45178
rect 18495 45126 18507 45178
rect 18507 45126 18537 45178
rect 18561 45126 18571 45178
rect 18571 45126 18617 45178
rect 18321 45124 18377 45126
rect 18401 45124 18457 45126
rect 18481 45124 18537 45126
rect 18561 45124 18617 45126
rect 18321 44090 18377 44092
rect 18401 44090 18457 44092
rect 18481 44090 18537 44092
rect 18561 44090 18617 44092
rect 18321 44038 18367 44090
rect 18367 44038 18377 44090
rect 18401 44038 18431 44090
rect 18431 44038 18443 44090
rect 18443 44038 18457 44090
rect 18481 44038 18495 44090
rect 18495 44038 18507 44090
rect 18507 44038 18537 44090
rect 18561 44038 18571 44090
rect 18571 44038 18617 44090
rect 18321 44036 18377 44038
rect 18401 44036 18457 44038
rect 18481 44036 18537 44038
rect 18561 44036 18617 44038
rect 21794 45722 21850 45724
rect 21874 45722 21930 45724
rect 21954 45722 22010 45724
rect 22034 45722 22090 45724
rect 21794 45670 21840 45722
rect 21840 45670 21850 45722
rect 21874 45670 21904 45722
rect 21904 45670 21916 45722
rect 21916 45670 21930 45722
rect 21954 45670 21968 45722
rect 21968 45670 21980 45722
rect 21980 45670 22010 45722
rect 22034 45670 22044 45722
rect 22044 45670 22090 45722
rect 21794 45668 21850 45670
rect 21874 45668 21930 45670
rect 21954 45668 22010 45670
rect 22034 45668 22090 45670
rect 18321 43002 18377 43004
rect 18401 43002 18457 43004
rect 18481 43002 18537 43004
rect 18561 43002 18617 43004
rect 18321 42950 18367 43002
rect 18367 42950 18377 43002
rect 18401 42950 18431 43002
rect 18431 42950 18443 43002
rect 18443 42950 18457 43002
rect 18481 42950 18495 43002
rect 18495 42950 18507 43002
rect 18507 42950 18537 43002
rect 18561 42950 18571 43002
rect 18571 42950 18617 43002
rect 18321 42948 18377 42950
rect 18401 42948 18457 42950
rect 18481 42948 18537 42950
rect 18561 42948 18617 42950
rect 19430 42880 19486 42936
rect 14848 42458 14904 42460
rect 14928 42458 14984 42460
rect 15008 42458 15064 42460
rect 15088 42458 15144 42460
rect 14848 42406 14894 42458
rect 14894 42406 14904 42458
rect 14928 42406 14958 42458
rect 14958 42406 14970 42458
rect 14970 42406 14984 42458
rect 15008 42406 15022 42458
rect 15022 42406 15034 42458
rect 15034 42406 15064 42458
rect 15088 42406 15098 42458
rect 15098 42406 15144 42458
rect 14848 42404 14904 42406
rect 14928 42404 14984 42406
rect 15008 42404 15064 42406
rect 15088 42404 15144 42406
rect 18321 41914 18377 41916
rect 18401 41914 18457 41916
rect 18481 41914 18537 41916
rect 18561 41914 18617 41916
rect 18321 41862 18367 41914
rect 18367 41862 18377 41914
rect 18401 41862 18431 41914
rect 18431 41862 18443 41914
rect 18443 41862 18457 41914
rect 18481 41862 18495 41914
rect 18495 41862 18507 41914
rect 18507 41862 18537 41914
rect 18561 41862 18571 41914
rect 18571 41862 18617 41914
rect 18321 41860 18377 41862
rect 18401 41860 18457 41862
rect 18481 41860 18537 41862
rect 18561 41860 18617 41862
rect 14848 41370 14904 41372
rect 14928 41370 14984 41372
rect 15008 41370 15064 41372
rect 15088 41370 15144 41372
rect 14848 41318 14894 41370
rect 14894 41318 14904 41370
rect 14928 41318 14958 41370
rect 14958 41318 14970 41370
rect 14970 41318 14984 41370
rect 15008 41318 15022 41370
rect 15022 41318 15034 41370
rect 15034 41318 15064 41370
rect 15088 41318 15098 41370
rect 15098 41318 15144 41370
rect 14848 41316 14904 41318
rect 14928 41316 14984 41318
rect 15008 41316 15064 41318
rect 15088 41316 15144 41318
rect 18321 40826 18377 40828
rect 18401 40826 18457 40828
rect 18481 40826 18537 40828
rect 18561 40826 18617 40828
rect 18321 40774 18367 40826
rect 18367 40774 18377 40826
rect 18401 40774 18431 40826
rect 18431 40774 18443 40826
rect 18443 40774 18457 40826
rect 18481 40774 18495 40826
rect 18495 40774 18507 40826
rect 18507 40774 18537 40826
rect 18561 40774 18571 40826
rect 18571 40774 18617 40826
rect 18321 40772 18377 40774
rect 18401 40772 18457 40774
rect 18481 40772 18537 40774
rect 18561 40772 18617 40774
rect 14848 40282 14904 40284
rect 14928 40282 14984 40284
rect 15008 40282 15064 40284
rect 15088 40282 15144 40284
rect 14848 40230 14894 40282
rect 14894 40230 14904 40282
rect 14928 40230 14958 40282
rect 14958 40230 14970 40282
rect 14970 40230 14984 40282
rect 15008 40230 15022 40282
rect 15022 40230 15034 40282
rect 15034 40230 15064 40282
rect 15088 40230 15098 40282
rect 15098 40230 15144 40282
rect 14848 40228 14904 40230
rect 14928 40228 14984 40230
rect 15008 40228 15064 40230
rect 15088 40228 15144 40230
rect 14848 39194 14904 39196
rect 14928 39194 14984 39196
rect 15008 39194 15064 39196
rect 15088 39194 15144 39196
rect 14848 39142 14894 39194
rect 14894 39142 14904 39194
rect 14928 39142 14958 39194
rect 14958 39142 14970 39194
rect 14970 39142 14984 39194
rect 15008 39142 15022 39194
rect 15022 39142 15034 39194
rect 15034 39142 15064 39194
rect 15088 39142 15098 39194
rect 15098 39142 15144 39194
rect 14848 39140 14904 39142
rect 14928 39140 14984 39142
rect 15008 39140 15064 39142
rect 15088 39140 15144 39142
rect 14848 38106 14904 38108
rect 14928 38106 14984 38108
rect 15008 38106 15064 38108
rect 15088 38106 15144 38108
rect 14848 38054 14894 38106
rect 14894 38054 14904 38106
rect 14928 38054 14958 38106
rect 14958 38054 14970 38106
rect 14970 38054 14984 38106
rect 15008 38054 15022 38106
rect 15022 38054 15034 38106
rect 15034 38054 15064 38106
rect 15088 38054 15098 38106
rect 15098 38054 15144 38106
rect 14848 38052 14904 38054
rect 14928 38052 14984 38054
rect 15008 38052 15064 38054
rect 15088 38052 15144 38054
rect 14848 37018 14904 37020
rect 14928 37018 14984 37020
rect 15008 37018 15064 37020
rect 15088 37018 15144 37020
rect 14848 36966 14894 37018
rect 14894 36966 14904 37018
rect 14928 36966 14958 37018
rect 14958 36966 14970 37018
rect 14970 36966 14984 37018
rect 15008 36966 15022 37018
rect 15022 36966 15034 37018
rect 15034 36966 15064 37018
rect 15088 36966 15098 37018
rect 15098 36966 15144 37018
rect 14848 36964 14904 36966
rect 14928 36964 14984 36966
rect 15008 36964 15064 36966
rect 15088 36964 15144 36966
rect 14848 35930 14904 35932
rect 14928 35930 14984 35932
rect 15008 35930 15064 35932
rect 15088 35930 15144 35932
rect 14848 35878 14894 35930
rect 14894 35878 14904 35930
rect 14928 35878 14958 35930
rect 14958 35878 14970 35930
rect 14970 35878 14984 35930
rect 15008 35878 15022 35930
rect 15022 35878 15034 35930
rect 15034 35878 15064 35930
rect 15088 35878 15098 35930
rect 15098 35878 15144 35930
rect 14848 35876 14904 35878
rect 14928 35876 14984 35878
rect 15008 35876 15064 35878
rect 15088 35876 15144 35878
rect 14848 34842 14904 34844
rect 14928 34842 14984 34844
rect 15008 34842 15064 34844
rect 15088 34842 15144 34844
rect 14848 34790 14894 34842
rect 14894 34790 14904 34842
rect 14928 34790 14958 34842
rect 14958 34790 14970 34842
rect 14970 34790 14984 34842
rect 15008 34790 15022 34842
rect 15022 34790 15034 34842
rect 15034 34790 15064 34842
rect 15088 34790 15098 34842
rect 15098 34790 15144 34842
rect 14848 34788 14904 34790
rect 14928 34788 14984 34790
rect 15008 34788 15064 34790
rect 15088 34788 15144 34790
rect 14848 33754 14904 33756
rect 14928 33754 14984 33756
rect 15008 33754 15064 33756
rect 15088 33754 15144 33756
rect 14848 33702 14894 33754
rect 14894 33702 14904 33754
rect 14928 33702 14958 33754
rect 14958 33702 14970 33754
rect 14970 33702 14984 33754
rect 15008 33702 15022 33754
rect 15022 33702 15034 33754
rect 15034 33702 15064 33754
rect 15088 33702 15098 33754
rect 15098 33702 15144 33754
rect 14848 33700 14904 33702
rect 14928 33700 14984 33702
rect 15008 33700 15064 33702
rect 15088 33700 15144 33702
rect 14848 32666 14904 32668
rect 14928 32666 14984 32668
rect 15008 32666 15064 32668
rect 15088 32666 15144 32668
rect 14848 32614 14894 32666
rect 14894 32614 14904 32666
rect 14928 32614 14958 32666
rect 14958 32614 14970 32666
rect 14970 32614 14984 32666
rect 15008 32614 15022 32666
rect 15022 32614 15034 32666
rect 15034 32614 15064 32666
rect 15088 32614 15098 32666
rect 15098 32614 15144 32666
rect 14848 32612 14904 32614
rect 14928 32612 14984 32614
rect 15008 32612 15064 32614
rect 15088 32612 15144 32614
rect 14848 31578 14904 31580
rect 14928 31578 14984 31580
rect 15008 31578 15064 31580
rect 15088 31578 15144 31580
rect 14848 31526 14894 31578
rect 14894 31526 14904 31578
rect 14928 31526 14958 31578
rect 14958 31526 14970 31578
rect 14970 31526 14984 31578
rect 15008 31526 15022 31578
rect 15022 31526 15034 31578
rect 15034 31526 15064 31578
rect 15088 31526 15098 31578
rect 15098 31526 15144 31578
rect 14848 31524 14904 31526
rect 14928 31524 14984 31526
rect 15008 31524 15064 31526
rect 15088 31524 15144 31526
rect 14848 30490 14904 30492
rect 14928 30490 14984 30492
rect 15008 30490 15064 30492
rect 15088 30490 15144 30492
rect 14848 30438 14894 30490
rect 14894 30438 14904 30490
rect 14928 30438 14958 30490
rect 14958 30438 14970 30490
rect 14970 30438 14984 30490
rect 15008 30438 15022 30490
rect 15022 30438 15034 30490
rect 15034 30438 15064 30490
rect 15088 30438 15098 30490
rect 15098 30438 15144 30490
rect 14848 30436 14904 30438
rect 14928 30436 14984 30438
rect 15008 30436 15064 30438
rect 15088 30436 15144 30438
rect 14848 29402 14904 29404
rect 14928 29402 14984 29404
rect 15008 29402 15064 29404
rect 15088 29402 15144 29404
rect 14848 29350 14894 29402
rect 14894 29350 14904 29402
rect 14928 29350 14958 29402
rect 14958 29350 14970 29402
rect 14970 29350 14984 29402
rect 15008 29350 15022 29402
rect 15022 29350 15034 29402
rect 15034 29350 15064 29402
rect 15088 29350 15098 29402
rect 15098 29350 15144 29402
rect 14848 29348 14904 29350
rect 14928 29348 14984 29350
rect 15008 29348 15064 29350
rect 15088 29348 15144 29350
rect 14848 28314 14904 28316
rect 14928 28314 14984 28316
rect 15008 28314 15064 28316
rect 15088 28314 15144 28316
rect 14848 28262 14894 28314
rect 14894 28262 14904 28314
rect 14928 28262 14958 28314
rect 14958 28262 14970 28314
rect 14970 28262 14984 28314
rect 15008 28262 15022 28314
rect 15022 28262 15034 28314
rect 15034 28262 15064 28314
rect 15088 28262 15098 28314
rect 15098 28262 15144 28314
rect 14848 28260 14904 28262
rect 14928 28260 14984 28262
rect 15008 28260 15064 28262
rect 15088 28260 15144 28262
rect 14848 27226 14904 27228
rect 14928 27226 14984 27228
rect 15008 27226 15064 27228
rect 15088 27226 15144 27228
rect 14848 27174 14894 27226
rect 14894 27174 14904 27226
rect 14928 27174 14958 27226
rect 14958 27174 14970 27226
rect 14970 27174 14984 27226
rect 15008 27174 15022 27226
rect 15022 27174 15034 27226
rect 15034 27174 15064 27226
rect 15088 27174 15098 27226
rect 15098 27174 15144 27226
rect 14848 27172 14904 27174
rect 14928 27172 14984 27174
rect 15008 27172 15064 27174
rect 15088 27172 15144 27174
rect 14848 26138 14904 26140
rect 14928 26138 14984 26140
rect 15008 26138 15064 26140
rect 15088 26138 15144 26140
rect 14848 26086 14894 26138
rect 14894 26086 14904 26138
rect 14928 26086 14958 26138
rect 14958 26086 14970 26138
rect 14970 26086 14984 26138
rect 15008 26086 15022 26138
rect 15022 26086 15034 26138
rect 15034 26086 15064 26138
rect 15088 26086 15098 26138
rect 15098 26086 15144 26138
rect 14848 26084 14904 26086
rect 14928 26084 14984 26086
rect 15008 26084 15064 26086
rect 15088 26084 15144 26086
rect 14848 25050 14904 25052
rect 14928 25050 14984 25052
rect 15008 25050 15064 25052
rect 15088 25050 15144 25052
rect 14848 24998 14894 25050
rect 14894 24998 14904 25050
rect 14928 24998 14958 25050
rect 14958 24998 14970 25050
rect 14970 24998 14984 25050
rect 15008 24998 15022 25050
rect 15022 24998 15034 25050
rect 15034 24998 15064 25050
rect 15088 24998 15098 25050
rect 15098 24998 15144 25050
rect 14848 24996 14904 24998
rect 14928 24996 14984 24998
rect 15008 24996 15064 24998
rect 15088 24996 15144 24998
rect 14848 23962 14904 23964
rect 14928 23962 14984 23964
rect 15008 23962 15064 23964
rect 15088 23962 15144 23964
rect 14848 23910 14894 23962
rect 14894 23910 14904 23962
rect 14928 23910 14958 23962
rect 14958 23910 14970 23962
rect 14970 23910 14984 23962
rect 15008 23910 15022 23962
rect 15022 23910 15034 23962
rect 15034 23910 15064 23962
rect 15088 23910 15098 23962
rect 15098 23910 15144 23962
rect 14848 23908 14904 23910
rect 14928 23908 14984 23910
rect 15008 23908 15064 23910
rect 15088 23908 15144 23910
rect 14848 22874 14904 22876
rect 14928 22874 14984 22876
rect 15008 22874 15064 22876
rect 15088 22874 15144 22876
rect 14848 22822 14894 22874
rect 14894 22822 14904 22874
rect 14928 22822 14958 22874
rect 14958 22822 14970 22874
rect 14970 22822 14984 22874
rect 15008 22822 15022 22874
rect 15022 22822 15034 22874
rect 15034 22822 15064 22874
rect 15088 22822 15098 22874
rect 15098 22822 15144 22874
rect 14848 22820 14904 22822
rect 14928 22820 14984 22822
rect 15008 22820 15064 22822
rect 15088 22820 15144 22822
rect 14848 21786 14904 21788
rect 14928 21786 14984 21788
rect 15008 21786 15064 21788
rect 15088 21786 15144 21788
rect 14848 21734 14894 21786
rect 14894 21734 14904 21786
rect 14928 21734 14958 21786
rect 14958 21734 14970 21786
rect 14970 21734 14984 21786
rect 15008 21734 15022 21786
rect 15022 21734 15034 21786
rect 15034 21734 15064 21786
rect 15088 21734 15098 21786
rect 15098 21734 15144 21786
rect 14848 21732 14904 21734
rect 14928 21732 14984 21734
rect 15008 21732 15064 21734
rect 15088 21732 15144 21734
rect 14848 20698 14904 20700
rect 14928 20698 14984 20700
rect 15008 20698 15064 20700
rect 15088 20698 15144 20700
rect 14848 20646 14894 20698
rect 14894 20646 14904 20698
rect 14928 20646 14958 20698
rect 14958 20646 14970 20698
rect 14970 20646 14984 20698
rect 15008 20646 15022 20698
rect 15022 20646 15034 20698
rect 15034 20646 15064 20698
rect 15088 20646 15098 20698
rect 15098 20646 15144 20698
rect 14848 20644 14904 20646
rect 14928 20644 14984 20646
rect 15008 20644 15064 20646
rect 15088 20644 15144 20646
rect 18321 39738 18377 39740
rect 18401 39738 18457 39740
rect 18481 39738 18537 39740
rect 18561 39738 18617 39740
rect 18321 39686 18367 39738
rect 18367 39686 18377 39738
rect 18401 39686 18431 39738
rect 18431 39686 18443 39738
rect 18443 39686 18457 39738
rect 18481 39686 18495 39738
rect 18495 39686 18507 39738
rect 18507 39686 18537 39738
rect 18561 39686 18571 39738
rect 18571 39686 18617 39738
rect 18321 39684 18377 39686
rect 18401 39684 18457 39686
rect 18481 39684 18537 39686
rect 18561 39684 18617 39686
rect 18321 38650 18377 38652
rect 18401 38650 18457 38652
rect 18481 38650 18537 38652
rect 18561 38650 18617 38652
rect 18321 38598 18367 38650
rect 18367 38598 18377 38650
rect 18401 38598 18431 38650
rect 18431 38598 18443 38650
rect 18443 38598 18457 38650
rect 18481 38598 18495 38650
rect 18495 38598 18507 38650
rect 18507 38598 18537 38650
rect 18561 38598 18571 38650
rect 18571 38598 18617 38650
rect 18321 38596 18377 38598
rect 18401 38596 18457 38598
rect 18481 38596 18537 38598
rect 18561 38596 18617 38598
rect 18321 37562 18377 37564
rect 18401 37562 18457 37564
rect 18481 37562 18537 37564
rect 18561 37562 18617 37564
rect 18321 37510 18367 37562
rect 18367 37510 18377 37562
rect 18401 37510 18431 37562
rect 18431 37510 18443 37562
rect 18443 37510 18457 37562
rect 18481 37510 18495 37562
rect 18495 37510 18507 37562
rect 18507 37510 18537 37562
rect 18561 37510 18571 37562
rect 18571 37510 18617 37562
rect 18321 37508 18377 37510
rect 18401 37508 18457 37510
rect 18481 37508 18537 37510
rect 18561 37508 18617 37510
rect 18321 36474 18377 36476
rect 18401 36474 18457 36476
rect 18481 36474 18537 36476
rect 18561 36474 18617 36476
rect 18321 36422 18367 36474
rect 18367 36422 18377 36474
rect 18401 36422 18431 36474
rect 18431 36422 18443 36474
rect 18443 36422 18457 36474
rect 18481 36422 18495 36474
rect 18495 36422 18507 36474
rect 18507 36422 18537 36474
rect 18561 36422 18571 36474
rect 18571 36422 18617 36474
rect 18321 36420 18377 36422
rect 18401 36420 18457 36422
rect 18481 36420 18537 36422
rect 18561 36420 18617 36422
rect 18321 35386 18377 35388
rect 18401 35386 18457 35388
rect 18481 35386 18537 35388
rect 18561 35386 18617 35388
rect 18321 35334 18367 35386
rect 18367 35334 18377 35386
rect 18401 35334 18431 35386
rect 18431 35334 18443 35386
rect 18443 35334 18457 35386
rect 18481 35334 18495 35386
rect 18495 35334 18507 35386
rect 18507 35334 18537 35386
rect 18561 35334 18571 35386
rect 18571 35334 18617 35386
rect 18321 35332 18377 35334
rect 18401 35332 18457 35334
rect 18481 35332 18537 35334
rect 18561 35332 18617 35334
rect 18321 34298 18377 34300
rect 18401 34298 18457 34300
rect 18481 34298 18537 34300
rect 18561 34298 18617 34300
rect 18321 34246 18367 34298
rect 18367 34246 18377 34298
rect 18401 34246 18431 34298
rect 18431 34246 18443 34298
rect 18443 34246 18457 34298
rect 18481 34246 18495 34298
rect 18495 34246 18507 34298
rect 18507 34246 18537 34298
rect 18561 34246 18571 34298
rect 18571 34246 18617 34298
rect 18321 34244 18377 34246
rect 18401 34244 18457 34246
rect 18481 34244 18537 34246
rect 18561 34244 18617 34246
rect 18321 33210 18377 33212
rect 18401 33210 18457 33212
rect 18481 33210 18537 33212
rect 18561 33210 18617 33212
rect 18321 33158 18367 33210
rect 18367 33158 18377 33210
rect 18401 33158 18431 33210
rect 18431 33158 18443 33210
rect 18443 33158 18457 33210
rect 18481 33158 18495 33210
rect 18495 33158 18507 33210
rect 18507 33158 18537 33210
rect 18561 33158 18571 33210
rect 18571 33158 18617 33210
rect 18321 33156 18377 33158
rect 18401 33156 18457 33158
rect 18481 33156 18537 33158
rect 18561 33156 18617 33158
rect 18321 32122 18377 32124
rect 18401 32122 18457 32124
rect 18481 32122 18537 32124
rect 18561 32122 18617 32124
rect 18321 32070 18367 32122
rect 18367 32070 18377 32122
rect 18401 32070 18431 32122
rect 18431 32070 18443 32122
rect 18443 32070 18457 32122
rect 18481 32070 18495 32122
rect 18495 32070 18507 32122
rect 18507 32070 18537 32122
rect 18561 32070 18571 32122
rect 18571 32070 18617 32122
rect 18321 32068 18377 32070
rect 18401 32068 18457 32070
rect 18481 32068 18537 32070
rect 18561 32068 18617 32070
rect 18321 31034 18377 31036
rect 18401 31034 18457 31036
rect 18481 31034 18537 31036
rect 18561 31034 18617 31036
rect 18321 30982 18367 31034
rect 18367 30982 18377 31034
rect 18401 30982 18431 31034
rect 18431 30982 18443 31034
rect 18443 30982 18457 31034
rect 18481 30982 18495 31034
rect 18495 30982 18507 31034
rect 18507 30982 18537 31034
rect 18561 30982 18571 31034
rect 18571 30982 18617 31034
rect 18321 30980 18377 30982
rect 18401 30980 18457 30982
rect 18481 30980 18537 30982
rect 18561 30980 18617 30982
rect 18321 29946 18377 29948
rect 18401 29946 18457 29948
rect 18481 29946 18537 29948
rect 18561 29946 18617 29948
rect 18321 29894 18367 29946
rect 18367 29894 18377 29946
rect 18401 29894 18431 29946
rect 18431 29894 18443 29946
rect 18443 29894 18457 29946
rect 18481 29894 18495 29946
rect 18495 29894 18507 29946
rect 18507 29894 18537 29946
rect 18561 29894 18571 29946
rect 18571 29894 18617 29946
rect 18321 29892 18377 29894
rect 18401 29892 18457 29894
rect 18481 29892 18537 29894
rect 18561 29892 18617 29894
rect 14848 19610 14904 19612
rect 14928 19610 14984 19612
rect 15008 19610 15064 19612
rect 15088 19610 15144 19612
rect 14848 19558 14894 19610
rect 14894 19558 14904 19610
rect 14928 19558 14958 19610
rect 14958 19558 14970 19610
rect 14970 19558 14984 19610
rect 15008 19558 15022 19610
rect 15022 19558 15034 19610
rect 15034 19558 15064 19610
rect 15088 19558 15098 19610
rect 15098 19558 15144 19610
rect 14848 19556 14904 19558
rect 14928 19556 14984 19558
rect 15008 19556 15064 19558
rect 15088 19556 15144 19558
rect 14848 18522 14904 18524
rect 14928 18522 14984 18524
rect 15008 18522 15064 18524
rect 15088 18522 15144 18524
rect 14848 18470 14894 18522
rect 14894 18470 14904 18522
rect 14928 18470 14958 18522
rect 14958 18470 14970 18522
rect 14970 18470 14984 18522
rect 15008 18470 15022 18522
rect 15022 18470 15034 18522
rect 15034 18470 15064 18522
rect 15088 18470 15098 18522
rect 15098 18470 15144 18522
rect 14848 18468 14904 18470
rect 14928 18468 14984 18470
rect 15008 18468 15064 18470
rect 15088 18468 15144 18470
rect 14848 17434 14904 17436
rect 14928 17434 14984 17436
rect 15008 17434 15064 17436
rect 15088 17434 15144 17436
rect 14848 17382 14894 17434
rect 14894 17382 14904 17434
rect 14928 17382 14958 17434
rect 14958 17382 14970 17434
rect 14970 17382 14984 17434
rect 15008 17382 15022 17434
rect 15022 17382 15034 17434
rect 15034 17382 15064 17434
rect 15088 17382 15098 17434
rect 15098 17382 15144 17434
rect 14848 17380 14904 17382
rect 14928 17380 14984 17382
rect 15008 17380 15064 17382
rect 15088 17380 15144 17382
rect 18321 28858 18377 28860
rect 18401 28858 18457 28860
rect 18481 28858 18537 28860
rect 18561 28858 18617 28860
rect 18321 28806 18367 28858
rect 18367 28806 18377 28858
rect 18401 28806 18431 28858
rect 18431 28806 18443 28858
rect 18443 28806 18457 28858
rect 18481 28806 18495 28858
rect 18495 28806 18507 28858
rect 18507 28806 18537 28858
rect 18561 28806 18571 28858
rect 18571 28806 18617 28858
rect 18321 28804 18377 28806
rect 18401 28804 18457 28806
rect 18481 28804 18537 28806
rect 18561 28804 18617 28806
rect 18321 27770 18377 27772
rect 18401 27770 18457 27772
rect 18481 27770 18537 27772
rect 18561 27770 18617 27772
rect 18321 27718 18367 27770
rect 18367 27718 18377 27770
rect 18401 27718 18431 27770
rect 18431 27718 18443 27770
rect 18443 27718 18457 27770
rect 18481 27718 18495 27770
rect 18495 27718 18507 27770
rect 18507 27718 18537 27770
rect 18561 27718 18571 27770
rect 18571 27718 18617 27770
rect 18321 27716 18377 27718
rect 18401 27716 18457 27718
rect 18481 27716 18537 27718
rect 18561 27716 18617 27718
rect 18321 26682 18377 26684
rect 18401 26682 18457 26684
rect 18481 26682 18537 26684
rect 18561 26682 18617 26684
rect 18321 26630 18367 26682
rect 18367 26630 18377 26682
rect 18401 26630 18431 26682
rect 18431 26630 18443 26682
rect 18443 26630 18457 26682
rect 18481 26630 18495 26682
rect 18495 26630 18507 26682
rect 18507 26630 18537 26682
rect 18561 26630 18571 26682
rect 18571 26630 18617 26682
rect 18321 26628 18377 26630
rect 18401 26628 18457 26630
rect 18481 26628 18537 26630
rect 18561 26628 18617 26630
rect 18321 25594 18377 25596
rect 18401 25594 18457 25596
rect 18481 25594 18537 25596
rect 18561 25594 18617 25596
rect 18321 25542 18367 25594
rect 18367 25542 18377 25594
rect 18401 25542 18431 25594
rect 18431 25542 18443 25594
rect 18443 25542 18457 25594
rect 18481 25542 18495 25594
rect 18495 25542 18507 25594
rect 18507 25542 18537 25594
rect 18561 25542 18571 25594
rect 18571 25542 18617 25594
rect 18321 25540 18377 25542
rect 18401 25540 18457 25542
rect 18481 25540 18537 25542
rect 18561 25540 18617 25542
rect 18786 24676 18842 24712
rect 18786 24656 18788 24676
rect 18788 24656 18840 24676
rect 18840 24656 18842 24676
rect 18321 24506 18377 24508
rect 18401 24506 18457 24508
rect 18481 24506 18537 24508
rect 18561 24506 18617 24508
rect 18321 24454 18367 24506
rect 18367 24454 18377 24506
rect 18401 24454 18431 24506
rect 18431 24454 18443 24506
rect 18443 24454 18457 24506
rect 18481 24454 18495 24506
rect 18495 24454 18507 24506
rect 18507 24454 18537 24506
rect 18561 24454 18571 24506
rect 18571 24454 18617 24506
rect 18321 24452 18377 24454
rect 18401 24452 18457 24454
rect 18481 24452 18537 24454
rect 18561 24452 18617 24454
rect 18321 23418 18377 23420
rect 18401 23418 18457 23420
rect 18481 23418 18537 23420
rect 18561 23418 18617 23420
rect 18321 23366 18367 23418
rect 18367 23366 18377 23418
rect 18401 23366 18431 23418
rect 18431 23366 18443 23418
rect 18443 23366 18457 23418
rect 18481 23366 18495 23418
rect 18495 23366 18507 23418
rect 18507 23366 18537 23418
rect 18561 23366 18571 23418
rect 18571 23366 18617 23418
rect 18321 23364 18377 23366
rect 18401 23364 18457 23366
rect 18481 23364 18537 23366
rect 18561 23364 18617 23366
rect 18321 22330 18377 22332
rect 18401 22330 18457 22332
rect 18481 22330 18537 22332
rect 18561 22330 18617 22332
rect 18321 22278 18367 22330
rect 18367 22278 18377 22330
rect 18401 22278 18431 22330
rect 18431 22278 18443 22330
rect 18443 22278 18457 22330
rect 18481 22278 18495 22330
rect 18495 22278 18507 22330
rect 18507 22278 18537 22330
rect 18561 22278 18571 22330
rect 18571 22278 18617 22330
rect 18321 22276 18377 22278
rect 18401 22276 18457 22278
rect 18481 22276 18537 22278
rect 18561 22276 18617 22278
rect 18321 21242 18377 21244
rect 18401 21242 18457 21244
rect 18481 21242 18537 21244
rect 18561 21242 18617 21244
rect 18321 21190 18367 21242
rect 18367 21190 18377 21242
rect 18401 21190 18431 21242
rect 18431 21190 18443 21242
rect 18443 21190 18457 21242
rect 18481 21190 18495 21242
rect 18495 21190 18507 21242
rect 18507 21190 18537 21242
rect 18561 21190 18571 21242
rect 18571 21190 18617 21242
rect 18321 21188 18377 21190
rect 18401 21188 18457 21190
rect 18481 21188 18537 21190
rect 18561 21188 18617 21190
rect 14848 16346 14904 16348
rect 14928 16346 14984 16348
rect 15008 16346 15064 16348
rect 15088 16346 15144 16348
rect 14848 16294 14894 16346
rect 14894 16294 14904 16346
rect 14928 16294 14958 16346
rect 14958 16294 14970 16346
rect 14970 16294 14984 16346
rect 15008 16294 15022 16346
rect 15022 16294 15034 16346
rect 15034 16294 15064 16346
rect 15088 16294 15098 16346
rect 15098 16294 15144 16346
rect 14848 16292 14904 16294
rect 14928 16292 14984 16294
rect 15008 16292 15064 16294
rect 15088 16292 15144 16294
rect 14848 15258 14904 15260
rect 14928 15258 14984 15260
rect 15008 15258 15064 15260
rect 15088 15258 15144 15260
rect 14848 15206 14894 15258
rect 14894 15206 14904 15258
rect 14928 15206 14958 15258
rect 14958 15206 14970 15258
rect 14970 15206 14984 15258
rect 15008 15206 15022 15258
rect 15022 15206 15034 15258
rect 15034 15206 15064 15258
rect 15088 15206 15098 15258
rect 15098 15206 15144 15258
rect 14848 15204 14904 15206
rect 14928 15204 14984 15206
rect 15008 15204 15064 15206
rect 15088 15204 15144 15206
rect 14848 14170 14904 14172
rect 14928 14170 14984 14172
rect 15008 14170 15064 14172
rect 15088 14170 15144 14172
rect 14848 14118 14894 14170
rect 14894 14118 14904 14170
rect 14928 14118 14958 14170
rect 14958 14118 14970 14170
rect 14970 14118 14984 14170
rect 15008 14118 15022 14170
rect 15022 14118 15034 14170
rect 15034 14118 15064 14170
rect 15088 14118 15098 14170
rect 15098 14118 15144 14170
rect 14848 14116 14904 14118
rect 14928 14116 14984 14118
rect 15008 14116 15064 14118
rect 15088 14116 15144 14118
rect 14848 13082 14904 13084
rect 14928 13082 14984 13084
rect 15008 13082 15064 13084
rect 15088 13082 15144 13084
rect 14848 13030 14894 13082
rect 14894 13030 14904 13082
rect 14928 13030 14958 13082
rect 14958 13030 14970 13082
rect 14970 13030 14984 13082
rect 15008 13030 15022 13082
rect 15022 13030 15034 13082
rect 15034 13030 15064 13082
rect 15088 13030 15098 13082
rect 15098 13030 15144 13082
rect 14848 13028 14904 13030
rect 14928 13028 14984 13030
rect 15008 13028 15064 13030
rect 15088 13028 15144 13030
rect 14848 11994 14904 11996
rect 14928 11994 14984 11996
rect 15008 11994 15064 11996
rect 15088 11994 15144 11996
rect 14848 11942 14894 11994
rect 14894 11942 14904 11994
rect 14928 11942 14958 11994
rect 14958 11942 14970 11994
rect 14970 11942 14984 11994
rect 15008 11942 15022 11994
rect 15022 11942 15034 11994
rect 15034 11942 15064 11994
rect 15088 11942 15098 11994
rect 15098 11942 15144 11994
rect 14848 11940 14904 11942
rect 14928 11940 14984 11942
rect 15008 11940 15064 11942
rect 15088 11940 15144 11942
rect 14848 10906 14904 10908
rect 14928 10906 14984 10908
rect 15008 10906 15064 10908
rect 15088 10906 15144 10908
rect 14848 10854 14894 10906
rect 14894 10854 14904 10906
rect 14928 10854 14958 10906
rect 14958 10854 14970 10906
rect 14970 10854 14984 10906
rect 15008 10854 15022 10906
rect 15022 10854 15034 10906
rect 15034 10854 15064 10906
rect 15088 10854 15098 10906
rect 15098 10854 15144 10906
rect 14848 10852 14904 10854
rect 14928 10852 14984 10854
rect 15008 10852 15064 10854
rect 15088 10852 15144 10854
rect 11375 8186 11431 8188
rect 11455 8186 11511 8188
rect 11535 8186 11591 8188
rect 11615 8186 11671 8188
rect 11375 8134 11421 8186
rect 11421 8134 11431 8186
rect 11455 8134 11485 8186
rect 11485 8134 11497 8186
rect 11497 8134 11511 8186
rect 11535 8134 11549 8186
rect 11549 8134 11561 8186
rect 11561 8134 11591 8186
rect 11615 8134 11625 8186
rect 11625 8134 11671 8186
rect 11375 8132 11431 8134
rect 11455 8132 11511 8134
rect 11535 8132 11591 8134
rect 11615 8132 11671 8134
rect 11375 7098 11431 7100
rect 11455 7098 11511 7100
rect 11535 7098 11591 7100
rect 11615 7098 11671 7100
rect 11375 7046 11421 7098
rect 11421 7046 11431 7098
rect 11455 7046 11485 7098
rect 11485 7046 11497 7098
rect 11497 7046 11511 7098
rect 11535 7046 11549 7098
rect 11549 7046 11561 7098
rect 11561 7046 11591 7098
rect 11615 7046 11625 7098
rect 11625 7046 11671 7098
rect 11375 7044 11431 7046
rect 11455 7044 11511 7046
rect 11535 7044 11591 7046
rect 11615 7044 11671 7046
rect 11375 6010 11431 6012
rect 11455 6010 11511 6012
rect 11535 6010 11591 6012
rect 11615 6010 11671 6012
rect 11375 5958 11421 6010
rect 11421 5958 11431 6010
rect 11455 5958 11485 6010
rect 11485 5958 11497 6010
rect 11497 5958 11511 6010
rect 11535 5958 11549 6010
rect 11549 5958 11561 6010
rect 11561 5958 11591 6010
rect 11615 5958 11625 6010
rect 11625 5958 11671 6010
rect 11375 5956 11431 5958
rect 11455 5956 11511 5958
rect 11535 5956 11591 5958
rect 11615 5956 11671 5958
rect 11375 4922 11431 4924
rect 11455 4922 11511 4924
rect 11535 4922 11591 4924
rect 11615 4922 11671 4924
rect 11375 4870 11421 4922
rect 11421 4870 11431 4922
rect 11455 4870 11485 4922
rect 11485 4870 11497 4922
rect 11497 4870 11511 4922
rect 11535 4870 11549 4922
rect 11549 4870 11561 4922
rect 11561 4870 11591 4922
rect 11615 4870 11625 4922
rect 11625 4870 11671 4922
rect 11375 4868 11431 4870
rect 11455 4868 11511 4870
rect 11535 4868 11591 4870
rect 11615 4868 11671 4870
rect 11375 3834 11431 3836
rect 11455 3834 11511 3836
rect 11535 3834 11591 3836
rect 11615 3834 11671 3836
rect 11375 3782 11421 3834
rect 11421 3782 11431 3834
rect 11455 3782 11485 3834
rect 11485 3782 11497 3834
rect 11497 3782 11511 3834
rect 11535 3782 11549 3834
rect 11549 3782 11561 3834
rect 11561 3782 11591 3834
rect 11615 3782 11625 3834
rect 11625 3782 11671 3834
rect 11375 3780 11431 3782
rect 11455 3780 11511 3782
rect 11535 3780 11591 3782
rect 11615 3780 11671 3782
rect 14848 9818 14904 9820
rect 14928 9818 14984 9820
rect 15008 9818 15064 9820
rect 15088 9818 15144 9820
rect 14848 9766 14894 9818
rect 14894 9766 14904 9818
rect 14928 9766 14958 9818
rect 14958 9766 14970 9818
rect 14970 9766 14984 9818
rect 15008 9766 15022 9818
rect 15022 9766 15034 9818
rect 15034 9766 15064 9818
rect 15088 9766 15098 9818
rect 15098 9766 15144 9818
rect 14848 9764 14904 9766
rect 14928 9764 14984 9766
rect 15008 9764 15064 9766
rect 15088 9764 15144 9766
rect 14848 8730 14904 8732
rect 14928 8730 14984 8732
rect 15008 8730 15064 8732
rect 15088 8730 15144 8732
rect 14848 8678 14894 8730
rect 14894 8678 14904 8730
rect 14928 8678 14958 8730
rect 14958 8678 14970 8730
rect 14970 8678 14984 8730
rect 15008 8678 15022 8730
rect 15022 8678 15034 8730
rect 15034 8678 15064 8730
rect 15088 8678 15098 8730
rect 15098 8678 15144 8730
rect 14848 8676 14904 8678
rect 14928 8676 14984 8678
rect 15008 8676 15064 8678
rect 15088 8676 15144 8678
rect 14848 7642 14904 7644
rect 14928 7642 14984 7644
rect 15008 7642 15064 7644
rect 15088 7642 15144 7644
rect 14848 7590 14894 7642
rect 14894 7590 14904 7642
rect 14928 7590 14958 7642
rect 14958 7590 14970 7642
rect 14970 7590 14984 7642
rect 15008 7590 15022 7642
rect 15022 7590 15034 7642
rect 15034 7590 15064 7642
rect 15088 7590 15098 7642
rect 15098 7590 15144 7642
rect 14848 7588 14904 7590
rect 14928 7588 14984 7590
rect 15008 7588 15064 7590
rect 15088 7588 15144 7590
rect 18321 20154 18377 20156
rect 18401 20154 18457 20156
rect 18481 20154 18537 20156
rect 18561 20154 18617 20156
rect 18321 20102 18367 20154
rect 18367 20102 18377 20154
rect 18401 20102 18431 20154
rect 18431 20102 18443 20154
rect 18443 20102 18457 20154
rect 18481 20102 18495 20154
rect 18495 20102 18507 20154
rect 18507 20102 18537 20154
rect 18561 20102 18571 20154
rect 18571 20102 18617 20154
rect 18321 20100 18377 20102
rect 18401 20100 18457 20102
rect 18481 20100 18537 20102
rect 18561 20100 18617 20102
rect 18694 19080 18750 19136
rect 18321 19066 18377 19068
rect 18401 19066 18457 19068
rect 18481 19066 18537 19068
rect 18561 19066 18617 19068
rect 18321 19014 18367 19066
rect 18367 19014 18377 19066
rect 18401 19014 18431 19066
rect 18431 19014 18443 19066
rect 18443 19014 18457 19066
rect 18481 19014 18495 19066
rect 18495 19014 18507 19066
rect 18507 19014 18537 19066
rect 18561 19014 18571 19066
rect 18571 19014 18617 19066
rect 18321 19012 18377 19014
rect 18401 19012 18457 19014
rect 18481 19012 18537 19014
rect 18561 19012 18617 19014
rect 18321 17978 18377 17980
rect 18401 17978 18457 17980
rect 18481 17978 18537 17980
rect 18561 17978 18617 17980
rect 18321 17926 18367 17978
rect 18367 17926 18377 17978
rect 18401 17926 18431 17978
rect 18431 17926 18443 17978
rect 18443 17926 18457 17978
rect 18481 17926 18495 17978
rect 18495 17926 18507 17978
rect 18507 17926 18537 17978
rect 18561 17926 18571 17978
rect 18571 17926 18617 17978
rect 18321 17924 18377 17926
rect 18401 17924 18457 17926
rect 18481 17924 18537 17926
rect 18561 17924 18617 17926
rect 18321 16890 18377 16892
rect 18401 16890 18457 16892
rect 18481 16890 18537 16892
rect 18561 16890 18617 16892
rect 18321 16838 18367 16890
rect 18367 16838 18377 16890
rect 18401 16838 18431 16890
rect 18431 16838 18443 16890
rect 18443 16838 18457 16890
rect 18481 16838 18495 16890
rect 18495 16838 18507 16890
rect 18507 16838 18537 16890
rect 18561 16838 18571 16890
rect 18571 16838 18617 16890
rect 18321 16836 18377 16838
rect 18401 16836 18457 16838
rect 18481 16836 18537 16838
rect 18561 16836 18617 16838
rect 19154 19116 19156 19136
rect 19156 19116 19208 19136
rect 19208 19116 19210 19136
rect 19154 19080 19210 19116
rect 21794 44634 21850 44636
rect 21874 44634 21930 44636
rect 21954 44634 22010 44636
rect 22034 44634 22090 44636
rect 21794 44582 21840 44634
rect 21840 44582 21850 44634
rect 21874 44582 21904 44634
rect 21904 44582 21916 44634
rect 21916 44582 21930 44634
rect 21954 44582 21968 44634
rect 21968 44582 21980 44634
rect 21980 44582 22010 44634
rect 22034 44582 22044 44634
rect 22044 44582 22090 44634
rect 21794 44580 21850 44582
rect 21874 44580 21930 44582
rect 21954 44580 22010 44582
rect 22034 44580 22090 44582
rect 21794 43546 21850 43548
rect 21874 43546 21930 43548
rect 21954 43546 22010 43548
rect 22034 43546 22090 43548
rect 21794 43494 21840 43546
rect 21840 43494 21850 43546
rect 21874 43494 21904 43546
rect 21904 43494 21916 43546
rect 21916 43494 21930 43546
rect 21954 43494 21968 43546
rect 21968 43494 21980 43546
rect 21980 43494 22010 43546
rect 22034 43494 22044 43546
rect 22044 43494 22090 43546
rect 21794 43492 21850 43494
rect 21874 43492 21930 43494
rect 21954 43492 22010 43494
rect 22034 43492 22090 43494
rect 21794 42458 21850 42460
rect 21874 42458 21930 42460
rect 21954 42458 22010 42460
rect 22034 42458 22090 42460
rect 21794 42406 21840 42458
rect 21840 42406 21850 42458
rect 21874 42406 21904 42458
rect 21904 42406 21916 42458
rect 21916 42406 21930 42458
rect 21954 42406 21968 42458
rect 21968 42406 21980 42458
rect 21980 42406 22010 42458
rect 22034 42406 22044 42458
rect 22044 42406 22090 42458
rect 21794 42404 21850 42406
rect 21874 42404 21930 42406
rect 21954 42404 22010 42406
rect 22034 42404 22090 42406
rect 21794 41370 21850 41372
rect 21874 41370 21930 41372
rect 21954 41370 22010 41372
rect 22034 41370 22090 41372
rect 21794 41318 21840 41370
rect 21840 41318 21850 41370
rect 21874 41318 21904 41370
rect 21904 41318 21916 41370
rect 21916 41318 21930 41370
rect 21954 41318 21968 41370
rect 21968 41318 21980 41370
rect 21980 41318 22010 41370
rect 22034 41318 22044 41370
rect 22044 41318 22090 41370
rect 21794 41316 21850 41318
rect 21874 41316 21930 41318
rect 21954 41316 22010 41318
rect 22034 41316 22090 41318
rect 21794 40282 21850 40284
rect 21874 40282 21930 40284
rect 21954 40282 22010 40284
rect 22034 40282 22090 40284
rect 21794 40230 21840 40282
rect 21840 40230 21850 40282
rect 21874 40230 21904 40282
rect 21904 40230 21916 40282
rect 21916 40230 21930 40282
rect 21954 40230 21968 40282
rect 21968 40230 21980 40282
rect 21980 40230 22010 40282
rect 22034 40230 22044 40282
rect 22044 40230 22090 40282
rect 21794 40228 21850 40230
rect 21874 40228 21930 40230
rect 21954 40228 22010 40230
rect 22034 40228 22090 40230
rect 21794 39194 21850 39196
rect 21874 39194 21930 39196
rect 21954 39194 22010 39196
rect 22034 39194 22090 39196
rect 21794 39142 21840 39194
rect 21840 39142 21850 39194
rect 21874 39142 21904 39194
rect 21904 39142 21916 39194
rect 21916 39142 21930 39194
rect 21954 39142 21968 39194
rect 21968 39142 21980 39194
rect 21980 39142 22010 39194
rect 22034 39142 22044 39194
rect 22044 39142 22090 39194
rect 21794 39140 21850 39142
rect 21874 39140 21930 39142
rect 21954 39140 22010 39142
rect 22034 39140 22090 39142
rect 21794 38106 21850 38108
rect 21874 38106 21930 38108
rect 21954 38106 22010 38108
rect 22034 38106 22090 38108
rect 21794 38054 21840 38106
rect 21840 38054 21850 38106
rect 21874 38054 21904 38106
rect 21904 38054 21916 38106
rect 21916 38054 21930 38106
rect 21954 38054 21968 38106
rect 21968 38054 21980 38106
rect 21980 38054 22010 38106
rect 22034 38054 22044 38106
rect 22044 38054 22090 38106
rect 21794 38052 21850 38054
rect 21874 38052 21930 38054
rect 21954 38052 22010 38054
rect 22034 38052 22090 38054
rect 21794 37018 21850 37020
rect 21874 37018 21930 37020
rect 21954 37018 22010 37020
rect 22034 37018 22090 37020
rect 21794 36966 21840 37018
rect 21840 36966 21850 37018
rect 21874 36966 21904 37018
rect 21904 36966 21916 37018
rect 21916 36966 21930 37018
rect 21954 36966 21968 37018
rect 21968 36966 21980 37018
rect 21980 36966 22010 37018
rect 22034 36966 22044 37018
rect 22044 36966 22090 37018
rect 21794 36964 21850 36966
rect 21874 36964 21930 36966
rect 21954 36964 22010 36966
rect 22034 36964 22090 36966
rect 21794 35930 21850 35932
rect 21874 35930 21930 35932
rect 21954 35930 22010 35932
rect 22034 35930 22090 35932
rect 21794 35878 21840 35930
rect 21840 35878 21850 35930
rect 21874 35878 21904 35930
rect 21904 35878 21916 35930
rect 21916 35878 21930 35930
rect 21954 35878 21968 35930
rect 21968 35878 21980 35930
rect 21980 35878 22010 35930
rect 22034 35878 22044 35930
rect 22044 35878 22090 35930
rect 21794 35876 21850 35878
rect 21874 35876 21930 35878
rect 21954 35876 22010 35878
rect 22034 35876 22090 35878
rect 21794 34842 21850 34844
rect 21874 34842 21930 34844
rect 21954 34842 22010 34844
rect 22034 34842 22090 34844
rect 21794 34790 21840 34842
rect 21840 34790 21850 34842
rect 21874 34790 21904 34842
rect 21904 34790 21916 34842
rect 21916 34790 21930 34842
rect 21954 34790 21968 34842
rect 21968 34790 21980 34842
rect 21980 34790 22010 34842
rect 22034 34790 22044 34842
rect 22044 34790 22090 34842
rect 21794 34788 21850 34790
rect 21874 34788 21930 34790
rect 21954 34788 22010 34790
rect 22034 34788 22090 34790
rect 21794 33754 21850 33756
rect 21874 33754 21930 33756
rect 21954 33754 22010 33756
rect 22034 33754 22090 33756
rect 21794 33702 21840 33754
rect 21840 33702 21850 33754
rect 21874 33702 21904 33754
rect 21904 33702 21916 33754
rect 21916 33702 21930 33754
rect 21954 33702 21968 33754
rect 21968 33702 21980 33754
rect 21980 33702 22010 33754
rect 22034 33702 22044 33754
rect 22044 33702 22090 33754
rect 21794 33700 21850 33702
rect 21874 33700 21930 33702
rect 21954 33700 22010 33702
rect 22034 33700 22090 33702
rect 21794 32666 21850 32668
rect 21874 32666 21930 32668
rect 21954 32666 22010 32668
rect 22034 32666 22090 32668
rect 21794 32614 21840 32666
rect 21840 32614 21850 32666
rect 21874 32614 21904 32666
rect 21904 32614 21916 32666
rect 21916 32614 21930 32666
rect 21954 32614 21968 32666
rect 21968 32614 21980 32666
rect 21980 32614 22010 32666
rect 22034 32614 22044 32666
rect 22044 32614 22090 32666
rect 21794 32612 21850 32614
rect 21874 32612 21930 32614
rect 21954 32612 22010 32614
rect 22034 32612 22090 32614
rect 18321 15802 18377 15804
rect 18401 15802 18457 15804
rect 18481 15802 18537 15804
rect 18561 15802 18617 15804
rect 18321 15750 18367 15802
rect 18367 15750 18377 15802
rect 18401 15750 18431 15802
rect 18431 15750 18443 15802
rect 18443 15750 18457 15802
rect 18481 15750 18495 15802
rect 18495 15750 18507 15802
rect 18507 15750 18537 15802
rect 18561 15750 18571 15802
rect 18571 15750 18617 15802
rect 18321 15748 18377 15750
rect 18401 15748 18457 15750
rect 18481 15748 18537 15750
rect 18561 15748 18617 15750
rect 18321 14714 18377 14716
rect 18401 14714 18457 14716
rect 18481 14714 18537 14716
rect 18561 14714 18617 14716
rect 18321 14662 18367 14714
rect 18367 14662 18377 14714
rect 18401 14662 18431 14714
rect 18431 14662 18443 14714
rect 18443 14662 18457 14714
rect 18481 14662 18495 14714
rect 18495 14662 18507 14714
rect 18507 14662 18537 14714
rect 18561 14662 18571 14714
rect 18571 14662 18617 14714
rect 18321 14660 18377 14662
rect 18401 14660 18457 14662
rect 18481 14660 18537 14662
rect 18561 14660 18617 14662
rect 14848 6554 14904 6556
rect 14928 6554 14984 6556
rect 15008 6554 15064 6556
rect 15088 6554 15144 6556
rect 14848 6502 14894 6554
rect 14894 6502 14904 6554
rect 14928 6502 14958 6554
rect 14958 6502 14970 6554
rect 14970 6502 14984 6554
rect 15008 6502 15022 6554
rect 15022 6502 15034 6554
rect 15034 6502 15064 6554
rect 15088 6502 15098 6554
rect 15098 6502 15144 6554
rect 14848 6500 14904 6502
rect 14928 6500 14984 6502
rect 15008 6500 15064 6502
rect 15088 6500 15144 6502
rect 14848 5466 14904 5468
rect 14928 5466 14984 5468
rect 15008 5466 15064 5468
rect 15088 5466 15144 5468
rect 14848 5414 14894 5466
rect 14894 5414 14904 5466
rect 14928 5414 14958 5466
rect 14958 5414 14970 5466
rect 14970 5414 14984 5466
rect 15008 5414 15022 5466
rect 15022 5414 15034 5466
rect 15034 5414 15064 5466
rect 15088 5414 15098 5466
rect 15098 5414 15144 5466
rect 14848 5412 14904 5414
rect 14928 5412 14984 5414
rect 15008 5412 15064 5414
rect 15088 5412 15144 5414
rect 14848 4378 14904 4380
rect 14928 4378 14984 4380
rect 15008 4378 15064 4380
rect 15088 4378 15144 4380
rect 14848 4326 14894 4378
rect 14894 4326 14904 4378
rect 14928 4326 14958 4378
rect 14958 4326 14970 4378
rect 14970 4326 14984 4378
rect 15008 4326 15022 4378
rect 15022 4326 15034 4378
rect 15034 4326 15064 4378
rect 15088 4326 15098 4378
rect 15098 4326 15144 4378
rect 14848 4324 14904 4326
rect 14928 4324 14984 4326
rect 15008 4324 15064 4326
rect 15088 4324 15144 4326
rect 11375 2746 11431 2748
rect 11455 2746 11511 2748
rect 11535 2746 11591 2748
rect 11615 2746 11671 2748
rect 11375 2694 11421 2746
rect 11421 2694 11431 2746
rect 11455 2694 11485 2746
rect 11485 2694 11497 2746
rect 11497 2694 11511 2746
rect 11535 2694 11549 2746
rect 11549 2694 11561 2746
rect 11561 2694 11591 2746
rect 11615 2694 11625 2746
rect 11625 2694 11671 2746
rect 11375 2692 11431 2694
rect 11455 2692 11511 2694
rect 11535 2692 11591 2694
rect 11615 2692 11671 2694
rect 14848 3290 14904 3292
rect 14928 3290 14984 3292
rect 15008 3290 15064 3292
rect 15088 3290 15144 3292
rect 14848 3238 14894 3290
rect 14894 3238 14904 3290
rect 14928 3238 14958 3290
rect 14958 3238 14970 3290
rect 14970 3238 14984 3290
rect 15008 3238 15022 3290
rect 15022 3238 15034 3290
rect 15034 3238 15064 3290
rect 15088 3238 15098 3290
rect 15098 3238 15144 3290
rect 14848 3236 14904 3238
rect 14928 3236 14984 3238
rect 15008 3236 15064 3238
rect 15088 3236 15144 3238
rect 14848 2202 14904 2204
rect 14928 2202 14984 2204
rect 15008 2202 15064 2204
rect 15088 2202 15144 2204
rect 14848 2150 14894 2202
rect 14894 2150 14904 2202
rect 14928 2150 14958 2202
rect 14958 2150 14970 2202
rect 14970 2150 14984 2202
rect 15008 2150 15022 2202
rect 15022 2150 15034 2202
rect 15034 2150 15064 2202
rect 15088 2150 15098 2202
rect 15098 2150 15144 2202
rect 14848 2148 14904 2150
rect 14928 2148 14984 2150
rect 15008 2148 15064 2150
rect 15088 2148 15144 2150
rect 18321 13626 18377 13628
rect 18401 13626 18457 13628
rect 18481 13626 18537 13628
rect 18561 13626 18617 13628
rect 18321 13574 18367 13626
rect 18367 13574 18377 13626
rect 18401 13574 18431 13626
rect 18431 13574 18443 13626
rect 18443 13574 18457 13626
rect 18481 13574 18495 13626
rect 18495 13574 18507 13626
rect 18507 13574 18537 13626
rect 18561 13574 18571 13626
rect 18571 13574 18617 13626
rect 18321 13572 18377 13574
rect 18401 13572 18457 13574
rect 18481 13572 18537 13574
rect 18561 13572 18617 13574
rect 18321 12538 18377 12540
rect 18401 12538 18457 12540
rect 18481 12538 18537 12540
rect 18561 12538 18617 12540
rect 18321 12486 18367 12538
rect 18367 12486 18377 12538
rect 18401 12486 18431 12538
rect 18431 12486 18443 12538
rect 18443 12486 18457 12538
rect 18481 12486 18495 12538
rect 18495 12486 18507 12538
rect 18507 12486 18537 12538
rect 18561 12486 18571 12538
rect 18571 12486 18617 12538
rect 18321 12484 18377 12486
rect 18401 12484 18457 12486
rect 18481 12484 18537 12486
rect 18561 12484 18617 12486
rect 18321 11450 18377 11452
rect 18401 11450 18457 11452
rect 18481 11450 18537 11452
rect 18561 11450 18617 11452
rect 18321 11398 18367 11450
rect 18367 11398 18377 11450
rect 18401 11398 18431 11450
rect 18431 11398 18443 11450
rect 18443 11398 18457 11450
rect 18481 11398 18495 11450
rect 18495 11398 18507 11450
rect 18507 11398 18537 11450
rect 18561 11398 18571 11450
rect 18571 11398 18617 11450
rect 18321 11396 18377 11398
rect 18401 11396 18457 11398
rect 18481 11396 18537 11398
rect 18561 11396 18617 11398
rect 26146 49000 26202 49056
rect 25267 47354 25323 47356
rect 25347 47354 25403 47356
rect 25427 47354 25483 47356
rect 25507 47354 25563 47356
rect 25267 47302 25313 47354
rect 25313 47302 25323 47354
rect 25347 47302 25377 47354
rect 25377 47302 25389 47354
rect 25389 47302 25403 47354
rect 25427 47302 25441 47354
rect 25441 47302 25453 47354
rect 25453 47302 25483 47354
rect 25507 47302 25517 47354
rect 25517 47302 25563 47354
rect 25267 47300 25323 47302
rect 25347 47300 25403 47302
rect 25427 47300 25483 47302
rect 25507 47300 25563 47302
rect 26054 46960 26110 47016
rect 25267 46266 25323 46268
rect 25347 46266 25403 46268
rect 25427 46266 25483 46268
rect 25507 46266 25563 46268
rect 25267 46214 25313 46266
rect 25313 46214 25323 46266
rect 25347 46214 25377 46266
rect 25377 46214 25389 46266
rect 25389 46214 25403 46266
rect 25427 46214 25441 46266
rect 25441 46214 25453 46266
rect 25453 46214 25483 46266
rect 25507 46214 25517 46266
rect 25517 46214 25563 46266
rect 25267 46212 25323 46214
rect 25347 46212 25403 46214
rect 25427 46212 25483 46214
rect 25507 46212 25563 46214
rect 25267 45178 25323 45180
rect 25347 45178 25403 45180
rect 25427 45178 25483 45180
rect 25507 45178 25563 45180
rect 25267 45126 25313 45178
rect 25313 45126 25323 45178
rect 25347 45126 25377 45178
rect 25377 45126 25389 45178
rect 25389 45126 25403 45178
rect 25427 45126 25441 45178
rect 25441 45126 25453 45178
rect 25453 45126 25483 45178
rect 25507 45126 25517 45178
rect 25517 45126 25563 45178
rect 25267 45124 25323 45126
rect 25347 45124 25403 45126
rect 25427 45124 25483 45126
rect 25507 45124 25563 45126
rect 25267 44090 25323 44092
rect 25347 44090 25403 44092
rect 25427 44090 25483 44092
rect 25507 44090 25563 44092
rect 25267 44038 25313 44090
rect 25313 44038 25323 44090
rect 25347 44038 25377 44090
rect 25377 44038 25389 44090
rect 25389 44038 25403 44090
rect 25427 44038 25441 44090
rect 25441 44038 25453 44090
rect 25453 44038 25483 44090
rect 25507 44038 25517 44090
rect 25517 44038 25563 44090
rect 25267 44036 25323 44038
rect 25347 44036 25403 44038
rect 25427 44036 25483 44038
rect 25507 44036 25563 44038
rect 25267 43002 25323 43004
rect 25347 43002 25403 43004
rect 25427 43002 25483 43004
rect 25507 43002 25563 43004
rect 25267 42950 25313 43002
rect 25313 42950 25323 43002
rect 25347 42950 25377 43002
rect 25377 42950 25389 43002
rect 25389 42950 25403 43002
rect 25427 42950 25441 43002
rect 25441 42950 25453 43002
rect 25453 42950 25483 43002
rect 25507 42950 25517 43002
rect 25517 42950 25563 43002
rect 25267 42948 25323 42950
rect 25347 42948 25403 42950
rect 25427 42948 25483 42950
rect 25507 42948 25563 42950
rect 26054 42200 26110 42256
rect 25267 41914 25323 41916
rect 25347 41914 25403 41916
rect 25427 41914 25483 41916
rect 25507 41914 25563 41916
rect 25267 41862 25313 41914
rect 25313 41862 25323 41914
rect 25347 41862 25377 41914
rect 25377 41862 25389 41914
rect 25389 41862 25403 41914
rect 25427 41862 25441 41914
rect 25441 41862 25453 41914
rect 25453 41862 25483 41914
rect 25507 41862 25517 41914
rect 25517 41862 25563 41914
rect 25267 41860 25323 41862
rect 25347 41860 25403 41862
rect 25427 41860 25483 41862
rect 25507 41860 25563 41862
rect 25267 40826 25323 40828
rect 25347 40826 25403 40828
rect 25427 40826 25483 40828
rect 25507 40826 25563 40828
rect 25267 40774 25313 40826
rect 25313 40774 25323 40826
rect 25347 40774 25377 40826
rect 25377 40774 25389 40826
rect 25389 40774 25403 40826
rect 25427 40774 25441 40826
rect 25441 40774 25453 40826
rect 25453 40774 25483 40826
rect 25507 40774 25517 40826
rect 25517 40774 25563 40826
rect 25267 40772 25323 40774
rect 25347 40772 25403 40774
rect 25427 40772 25483 40774
rect 25507 40772 25563 40774
rect 25267 39738 25323 39740
rect 25347 39738 25403 39740
rect 25427 39738 25483 39740
rect 25507 39738 25563 39740
rect 25267 39686 25313 39738
rect 25313 39686 25323 39738
rect 25347 39686 25377 39738
rect 25377 39686 25389 39738
rect 25389 39686 25403 39738
rect 25427 39686 25441 39738
rect 25441 39686 25453 39738
rect 25453 39686 25483 39738
rect 25507 39686 25517 39738
rect 25517 39686 25563 39738
rect 25267 39684 25323 39686
rect 25347 39684 25403 39686
rect 25427 39684 25483 39686
rect 25507 39684 25563 39686
rect 25267 38650 25323 38652
rect 25347 38650 25403 38652
rect 25427 38650 25483 38652
rect 25507 38650 25563 38652
rect 25267 38598 25313 38650
rect 25313 38598 25323 38650
rect 25347 38598 25377 38650
rect 25377 38598 25389 38650
rect 25389 38598 25403 38650
rect 25427 38598 25441 38650
rect 25441 38598 25453 38650
rect 25453 38598 25483 38650
rect 25507 38598 25517 38650
rect 25517 38598 25563 38650
rect 25267 38596 25323 38598
rect 25347 38596 25403 38598
rect 25427 38596 25483 38598
rect 25507 38596 25563 38598
rect 25267 37562 25323 37564
rect 25347 37562 25403 37564
rect 25427 37562 25483 37564
rect 25507 37562 25563 37564
rect 25267 37510 25313 37562
rect 25313 37510 25323 37562
rect 25347 37510 25377 37562
rect 25377 37510 25389 37562
rect 25389 37510 25403 37562
rect 25427 37510 25441 37562
rect 25441 37510 25453 37562
rect 25453 37510 25483 37562
rect 25507 37510 25517 37562
rect 25517 37510 25563 37562
rect 25267 37508 25323 37510
rect 25347 37508 25403 37510
rect 25427 37508 25483 37510
rect 25507 37508 25563 37510
rect 26146 39480 26202 39536
rect 21794 31578 21850 31580
rect 21874 31578 21930 31580
rect 21954 31578 22010 31580
rect 22034 31578 22090 31580
rect 21794 31526 21840 31578
rect 21840 31526 21850 31578
rect 21874 31526 21904 31578
rect 21904 31526 21916 31578
rect 21916 31526 21930 31578
rect 21954 31526 21968 31578
rect 21968 31526 21980 31578
rect 21980 31526 22010 31578
rect 22034 31526 22044 31578
rect 22044 31526 22090 31578
rect 21794 31524 21850 31526
rect 21874 31524 21930 31526
rect 21954 31524 22010 31526
rect 22034 31524 22090 31526
rect 21794 30490 21850 30492
rect 21874 30490 21930 30492
rect 21954 30490 22010 30492
rect 22034 30490 22090 30492
rect 21794 30438 21840 30490
rect 21840 30438 21850 30490
rect 21874 30438 21904 30490
rect 21904 30438 21916 30490
rect 21916 30438 21930 30490
rect 21954 30438 21968 30490
rect 21968 30438 21980 30490
rect 21980 30438 22010 30490
rect 22034 30438 22044 30490
rect 22044 30438 22090 30490
rect 21794 30436 21850 30438
rect 21874 30436 21930 30438
rect 21954 30436 22010 30438
rect 22034 30436 22090 30438
rect 21794 29402 21850 29404
rect 21874 29402 21930 29404
rect 21954 29402 22010 29404
rect 22034 29402 22090 29404
rect 21794 29350 21840 29402
rect 21840 29350 21850 29402
rect 21874 29350 21904 29402
rect 21904 29350 21916 29402
rect 21916 29350 21930 29402
rect 21954 29350 21968 29402
rect 21968 29350 21980 29402
rect 21980 29350 22010 29402
rect 22034 29350 22044 29402
rect 22044 29350 22090 29402
rect 21794 29348 21850 29350
rect 21874 29348 21930 29350
rect 21954 29348 22010 29350
rect 22034 29348 22090 29350
rect 21794 28314 21850 28316
rect 21874 28314 21930 28316
rect 21954 28314 22010 28316
rect 22034 28314 22090 28316
rect 21794 28262 21840 28314
rect 21840 28262 21850 28314
rect 21874 28262 21904 28314
rect 21904 28262 21916 28314
rect 21916 28262 21930 28314
rect 21954 28262 21968 28314
rect 21968 28262 21980 28314
rect 21980 28262 22010 28314
rect 22034 28262 22044 28314
rect 22044 28262 22090 28314
rect 21794 28260 21850 28262
rect 21874 28260 21930 28262
rect 21954 28260 22010 28262
rect 22034 28260 22090 28262
rect 21794 27226 21850 27228
rect 21874 27226 21930 27228
rect 21954 27226 22010 27228
rect 22034 27226 22090 27228
rect 21794 27174 21840 27226
rect 21840 27174 21850 27226
rect 21874 27174 21904 27226
rect 21904 27174 21916 27226
rect 21916 27174 21930 27226
rect 21954 27174 21968 27226
rect 21968 27174 21980 27226
rect 21980 27174 22010 27226
rect 22034 27174 22044 27226
rect 22044 27174 22090 27226
rect 21794 27172 21850 27174
rect 21874 27172 21930 27174
rect 21954 27172 22010 27174
rect 22034 27172 22090 27174
rect 21794 26138 21850 26140
rect 21874 26138 21930 26140
rect 21954 26138 22010 26140
rect 22034 26138 22090 26140
rect 21794 26086 21840 26138
rect 21840 26086 21850 26138
rect 21874 26086 21904 26138
rect 21904 26086 21916 26138
rect 21916 26086 21930 26138
rect 21954 26086 21968 26138
rect 21968 26086 21980 26138
rect 21980 26086 22010 26138
rect 22034 26086 22044 26138
rect 22044 26086 22090 26138
rect 21794 26084 21850 26086
rect 21874 26084 21930 26086
rect 21954 26084 22010 26086
rect 22034 26084 22090 26086
rect 21794 25050 21850 25052
rect 21874 25050 21930 25052
rect 21954 25050 22010 25052
rect 22034 25050 22090 25052
rect 21794 24998 21840 25050
rect 21840 24998 21850 25050
rect 21874 24998 21904 25050
rect 21904 24998 21916 25050
rect 21916 24998 21930 25050
rect 21954 24998 21968 25050
rect 21968 24998 21980 25050
rect 21980 24998 22010 25050
rect 22034 24998 22044 25050
rect 22044 24998 22090 25050
rect 21794 24996 21850 24998
rect 21874 24996 21930 24998
rect 21954 24996 22010 24998
rect 22034 24996 22090 24998
rect 21794 23962 21850 23964
rect 21874 23962 21930 23964
rect 21954 23962 22010 23964
rect 22034 23962 22090 23964
rect 21794 23910 21840 23962
rect 21840 23910 21850 23962
rect 21874 23910 21904 23962
rect 21904 23910 21916 23962
rect 21916 23910 21930 23962
rect 21954 23910 21968 23962
rect 21968 23910 21980 23962
rect 21980 23910 22010 23962
rect 22034 23910 22044 23962
rect 22044 23910 22090 23962
rect 21794 23908 21850 23910
rect 21874 23908 21930 23910
rect 21954 23908 22010 23910
rect 22034 23908 22090 23910
rect 21794 22874 21850 22876
rect 21874 22874 21930 22876
rect 21954 22874 22010 22876
rect 22034 22874 22090 22876
rect 21794 22822 21840 22874
rect 21840 22822 21850 22874
rect 21874 22822 21904 22874
rect 21904 22822 21916 22874
rect 21916 22822 21930 22874
rect 21954 22822 21968 22874
rect 21968 22822 21980 22874
rect 21980 22822 22010 22874
rect 22034 22822 22044 22874
rect 22044 22822 22090 22874
rect 21794 22820 21850 22822
rect 21874 22820 21930 22822
rect 21954 22820 22010 22822
rect 22034 22820 22090 22822
rect 21794 21786 21850 21788
rect 21874 21786 21930 21788
rect 21954 21786 22010 21788
rect 22034 21786 22090 21788
rect 21794 21734 21840 21786
rect 21840 21734 21850 21786
rect 21874 21734 21904 21786
rect 21904 21734 21916 21786
rect 21916 21734 21930 21786
rect 21954 21734 21968 21786
rect 21968 21734 21980 21786
rect 21980 21734 22010 21786
rect 22034 21734 22044 21786
rect 22044 21734 22090 21786
rect 21794 21732 21850 21734
rect 21874 21732 21930 21734
rect 21954 21732 22010 21734
rect 22034 21732 22090 21734
rect 21794 20698 21850 20700
rect 21874 20698 21930 20700
rect 21954 20698 22010 20700
rect 22034 20698 22090 20700
rect 21794 20646 21840 20698
rect 21840 20646 21850 20698
rect 21874 20646 21904 20698
rect 21904 20646 21916 20698
rect 21916 20646 21930 20698
rect 21954 20646 21968 20698
rect 21968 20646 21980 20698
rect 21980 20646 22010 20698
rect 22034 20646 22044 20698
rect 22044 20646 22090 20698
rect 21794 20644 21850 20646
rect 21874 20644 21930 20646
rect 21954 20644 22010 20646
rect 22034 20644 22090 20646
rect 21794 19610 21850 19612
rect 21874 19610 21930 19612
rect 21954 19610 22010 19612
rect 22034 19610 22090 19612
rect 21794 19558 21840 19610
rect 21840 19558 21850 19610
rect 21874 19558 21904 19610
rect 21904 19558 21916 19610
rect 21916 19558 21930 19610
rect 21954 19558 21968 19610
rect 21968 19558 21980 19610
rect 21980 19558 22010 19610
rect 22034 19558 22044 19610
rect 22044 19558 22090 19610
rect 21794 19556 21850 19558
rect 21874 19556 21930 19558
rect 21954 19556 22010 19558
rect 22034 19556 22090 19558
rect 21794 18522 21850 18524
rect 21874 18522 21930 18524
rect 21954 18522 22010 18524
rect 22034 18522 22090 18524
rect 21794 18470 21840 18522
rect 21840 18470 21850 18522
rect 21874 18470 21904 18522
rect 21904 18470 21916 18522
rect 21916 18470 21930 18522
rect 21954 18470 21968 18522
rect 21968 18470 21980 18522
rect 21980 18470 22010 18522
rect 22034 18470 22044 18522
rect 22044 18470 22090 18522
rect 21794 18468 21850 18470
rect 21874 18468 21930 18470
rect 21954 18468 22010 18470
rect 22034 18468 22090 18470
rect 25267 36474 25323 36476
rect 25347 36474 25403 36476
rect 25427 36474 25483 36476
rect 25507 36474 25563 36476
rect 25267 36422 25313 36474
rect 25313 36422 25323 36474
rect 25347 36422 25377 36474
rect 25377 36422 25389 36474
rect 25389 36422 25403 36474
rect 25427 36422 25441 36474
rect 25441 36422 25453 36474
rect 25453 36422 25483 36474
rect 25507 36422 25517 36474
rect 25517 36422 25563 36474
rect 25267 36420 25323 36422
rect 25347 36420 25403 36422
rect 25427 36420 25483 36422
rect 25507 36420 25563 36422
rect 25267 35386 25323 35388
rect 25347 35386 25403 35388
rect 25427 35386 25483 35388
rect 25507 35386 25563 35388
rect 25267 35334 25313 35386
rect 25313 35334 25323 35386
rect 25347 35334 25377 35386
rect 25377 35334 25389 35386
rect 25389 35334 25403 35386
rect 25427 35334 25441 35386
rect 25441 35334 25453 35386
rect 25453 35334 25483 35386
rect 25507 35334 25517 35386
rect 25517 35334 25563 35386
rect 25267 35332 25323 35334
rect 25347 35332 25403 35334
rect 25427 35332 25483 35334
rect 25507 35332 25563 35334
rect 25267 34298 25323 34300
rect 25347 34298 25403 34300
rect 25427 34298 25483 34300
rect 25507 34298 25563 34300
rect 25267 34246 25313 34298
rect 25313 34246 25323 34298
rect 25347 34246 25377 34298
rect 25377 34246 25389 34298
rect 25389 34246 25403 34298
rect 25427 34246 25441 34298
rect 25441 34246 25453 34298
rect 25453 34246 25483 34298
rect 25507 34246 25517 34298
rect 25517 34246 25563 34298
rect 25267 34244 25323 34246
rect 25347 34244 25403 34246
rect 25427 34244 25483 34246
rect 25507 34244 25563 34246
rect 25267 33210 25323 33212
rect 25347 33210 25403 33212
rect 25427 33210 25483 33212
rect 25507 33210 25563 33212
rect 25267 33158 25313 33210
rect 25313 33158 25323 33210
rect 25347 33158 25377 33210
rect 25377 33158 25389 33210
rect 25389 33158 25403 33210
rect 25427 33158 25441 33210
rect 25441 33158 25453 33210
rect 25453 33158 25483 33210
rect 25507 33158 25517 33210
rect 25517 33158 25563 33210
rect 25267 33156 25323 33158
rect 25347 33156 25403 33158
rect 25427 33156 25483 33158
rect 25507 33156 25563 33158
rect 25267 32122 25323 32124
rect 25347 32122 25403 32124
rect 25427 32122 25483 32124
rect 25507 32122 25563 32124
rect 25267 32070 25313 32122
rect 25313 32070 25323 32122
rect 25347 32070 25377 32122
rect 25377 32070 25389 32122
rect 25389 32070 25403 32122
rect 25427 32070 25441 32122
rect 25441 32070 25453 32122
rect 25453 32070 25483 32122
rect 25507 32070 25517 32122
rect 25517 32070 25563 32122
rect 25267 32068 25323 32070
rect 25347 32068 25403 32070
rect 25427 32068 25483 32070
rect 25507 32068 25563 32070
rect 27526 46280 27582 46336
rect 28262 47640 28318 47696
rect 28078 44920 28134 44976
rect 27526 41520 27582 41576
rect 27526 40588 27582 40624
rect 27526 40568 27528 40588
rect 27528 40568 27580 40588
rect 27580 40568 27582 40588
rect 28740 46810 28796 46812
rect 28820 46810 28876 46812
rect 28900 46810 28956 46812
rect 28980 46810 29036 46812
rect 28740 46758 28786 46810
rect 28786 46758 28796 46810
rect 28820 46758 28850 46810
rect 28850 46758 28862 46810
rect 28862 46758 28876 46810
rect 28900 46758 28914 46810
rect 28914 46758 28926 46810
rect 28926 46758 28956 46810
rect 28980 46758 28990 46810
rect 28990 46758 29036 46810
rect 28740 46756 28796 46758
rect 28820 46756 28876 46758
rect 28900 46756 28956 46758
rect 28980 46756 29036 46758
rect 28354 42880 28410 42936
rect 25267 31034 25323 31036
rect 25347 31034 25403 31036
rect 25427 31034 25483 31036
rect 25507 31034 25563 31036
rect 25267 30982 25313 31034
rect 25313 30982 25323 31034
rect 25347 30982 25377 31034
rect 25377 30982 25389 31034
rect 25389 30982 25403 31034
rect 25427 30982 25441 31034
rect 25441 30982 25453 31034
rect 25453 30982 25483 31034
rect 25507 30982 25517 31034
rect 25517 30982 25563 31034
rect 25267 30980 25323 30982
rect 25347 30980 25403 30982
rect 25427 30980 25483 30982
rect 25507 30980 25563 30982
rect 26146 30640 26202 30696
rect 25267 29946 25323 29948
rect 25347 29946 25403 29948
rect 25427 29946 25483 29948
rect 25507 29946 25563 29948
rect 25267 29894 25313 29946
rect 25313 29894 25323 29946
rect 25347 29894 25377 29946
rect 25377 29894 25389 29946
rect 25389 29894 25403 29946
rect 25427 29894 25441 29946
rect 25441 29894 25453 29946
rect 25453 29894 25483 29946
rect 25507 29894 25517 29946
rect 25517 29894 25563 29946
rect 25267 29892 25323 29894
rect 25347 29892 25403 29894
rect 25427 29892 25483 29894
rect 25507 29892 25563 29894
rect 24858 29008 24914 29064
rect 21794 17434 21850 17436
rect 21874 17434 21930 17436
rect 21954 17434 22010 17436
rect 22034 17434 22090 17436
rect 21794 17382 21840 17434
rect 21840 17382 21850 17434
rect 21874 17382 21904 17434
rect 21904 17382 21916 17434
rect 21916 17382 21930 17434
rect 21954 17382 21968 17434
rect 21968 17382 21980 17434
rect 21980 17382 22010 17434
rect 22034 17382 22044 17434
rect 22044 17382 22090 17434
rect 21794 17380 21850 17382
rect 21874 17380 21930 17382
rect 21954 17380 22010 17382
rect 22034 17380 22090 17382
rect 21794 16346 21850 16348
rect 21874 16346 21930 16348
rect 21954 16346 22010 16348
rect 22034 16346 22090 16348
rect 21794 16294 21840 16346
rect 21840 16294 21850 16346
rect 21874 16294 21904 16346
rect 21904 16294 21916 16346
rect 21916 16294 21930 16346
rect 21954 16294 21968 16346
rect 21968 16294 21980 16346
rect 21980 16294 22010 16346
rect 22034 16294 22044 16346
rect 22044 16294 22090 16346
rect 21794 16292 21850 16294
rect 21874 16292 21930 16294
rect 21954 16292 22010 16294
rect 22034 16292 22090 16294
rect 21794 15258 21850 15260
rect 21874 15258 21930 15260
rect 21954 15258 22010 15260
rect 22034 15258 22090 15260
rect 21794 15206 21840 15258
rect 21840 15206 21850 15258
rect 21874 15206 21904 15258
rect 21904 15206 21916 15258
rect 21916 15206 21930 15258
rect 21954 15206 21968 15258
rect 21968 15206 21980 15258
rect 21980 15206 22010 15258
rect 22034 15206 22044 15258
rect 22044 15206 22090 15258
rect 21794 15204 21850 15206
rect 21874 15204 21930 15206
rect 21954 15204 22010 15206
rect 22034 15204 22090 15206
rect 21794 14170 21850 14172
rect 21874 14170 21930 14172
rect 21954 14170 22010 14172
rect 22034 14170 22090 14172
rect 21794 14118 21840 14170
rect 21840 14118 21850 14170
rect 21874 14118 21904 14170
rect 21904 14118 21916 14170
rect 21916 14118 21930 14170
rect 21954 14118 21968 14170
rect 21968 14118 21980 14170
rect 21980 14118 22010 14170
rect 22034 14118 22044 14170
rect 22044 14118 22090 14170
rect 21794 14116 21850 14118
rect 21874 14116 21930 14118
rect 21954 14116 22010 14118
rect 22034 14116 22090 14118
rect 18321 10362 18377 10364
rect 18401 10362 18457 10364
rect 18481 10362 18537 10364
rect 18561 10362 18617 10364
rect 18321 10310 18367 10362
rect 18367 10310 18377 10362
rect 18401 10310 18431 10362
rect 18431 10310 18443 10362
rect 18443 10310 18457 10362
rect 18481 10310 18495 10362
rect 18495 10310 18507 10362
rect 18507 10310 18537 10362
rect 18561 10310 18571 10362
rect 18571 10310 18617 10362
rect 18321 10308 18377 10310
rect 18401 10308 18457 10310
rect 18481 10308 18537 10310
rect 18561 10308 18617 10310
rect 18321 9274 18377 9276
rect 18401 9274 18457 9276
rect 18481 9274 18537 9276
rect 18561 9274 18617 9276
rect 18321 9222 18367 9274
rect 18367 9222 18377 9274
rect 18401 9222 18431 9274
rect 18431 9222 18443 9274
rect 18443 9222 18457 9274
rect 18481 9222 18495 9274
rect 18495 9222 18507 9274
rect 18507 9222 18537 9274
rect 18561 9222 18571 9274
rect 18571 9222 18617 9274
rect 18321 9220 18377 9222
rect 18401 9220 18457 9222
rect 18481 9220 18537 9222
rect 18561 9220 18617 9222
rect 18321 8186 18377 8188
rect 18401 8186 18457 8188
rect 18481 8186 18537 8188
rect 18561 8186 18617 8188
rect 18321 8134 18367 8186
rect 18367 8134 18377 8186
rect 18401 8134 18431 8186
rect 18431 8134 18443 8186
rect 18443 8134 18457 8186
rect 18481 8134 18495 8186
rect 18495 8134 18507 8186
rect 18507 8134 18537 8186
rect 18561 8134 18571 8186
rect 18571 8134 18617 8186
rect 18321 8132 18377 8134
rect 18401 8132 18457 8134
rect 18481 8132 18537 8134
rect 18561 8132 18617 8134
rect 18321 7098 18377 7100
rect 18401 7098 18457 7100
rect 18481 7098 18537 7100
rect 18561 7098 18617 7100
rect 18321 7046 18367 7098
rect 18367 7046 18377 7098
rect 18401 7046 18431 7098
rect 18431 7046 18443 7098
rect 18443 7046 18457 7098
rect 18481 7046 18495 7098
rect 18495 7046 18507 7098
rect 18507 7046 18537 7098
rect 18561 7046 18571 7098
rect 18571 7046 18617 7098
rect 18321 7044 18377 7046
rect 18401 7044 18457 7046
rect 18481 7044 18537 7046
rect 18561 7044 18617 7046
rect 21794 13082 21850 13084
rect 21874 13082 21930 13084
rect 21954 13082 22010 13084
rect 22034 13082 22090 13084
rect 21794 13030 21840 13082
rect 21840 13030 21850 13082
rect 21874 13030 21904 13082
rect 21904 13030 21916 13082
rect 21916 13030 21930 13082
rect 21954 13030 21968 13082
rect 21968 13030 21980 13082
rect 21980 13030 22010 13082
rect 22034 13030 22044 13082
rect 22044 13030 22090 13082
rect 21794 13028 21850 13030
rect 21874 13028 21930 13030
rect 21954 13028 22010 13030
rect 22034 13028 22090 13030
rect 21794 11994 21850 11996
rect 21874 11994 21930 11996
rect 21954 11994 22010 11996
rect 22034 11994 22090 11996
rect 21794 11942 21840 11994
rect 21840 11942 21850 11994
rect 21874 11942 21904 11994
rect 21904 11942 21916 11994
rect 21916 11942 21930 11994
rect 21954 11942 21968 11994
rect 21968 11942 21980 11994
rect 21980 11942 22010 11994
rect 22034 11942 22044 11994
rect 22044 11942 22090 11994
rect 21794 11940 21850 11942
rect 21874 11940 21930 11942
rect 21954 11940 22010 11942
rect 22034 11940 22090 11942
rect 21794 10906 21850 10908
rect 21874 10906 21930 10908
rect 21954 10906 22010 10908
rect 22034 10906 22090 10908
rect 21794 10854 21840 10906
rect 21840 10854 21850 10906
rect 21874 10854 21904 10906
rect 21904 10854 21916 10906
rect 21916 10854 21930 10906
rect 21954 10854 21968 10906
rect 21968 10854 21980 10906
rect 21980 10854 22010 10906
rect 22034 10854 22044 10906
rect 22044 10854 22090 10906
rect 21794 10852 21850 10854
rect 21874 10852 21930 10854
rect 21954 10852 22010 10854
rect 22034 10852 22090 10854
rect 25267 28858 25323 28860
rect 25347 28858 25403 28860
rect 25427 28858 25483 28860
rect 25507 28858 25563 28860
rect 25267 28806 25313 28858
rect 25313 28806 25323 28858
rect 25347 28806 25377 28858
rect 25377 28806 25389 28858
rect 25389 28806 25403 28858
rect 25427 28806 25441 28858
rect 25441 28806 25453 28858
rect 25453 28806 25483 28858
rect 25507 28806 25517 28858
rect 25517 28806 25563 28858
rect 25267 28804 25323 28806
rect 25347 28804 25403 28806
rect 25427 28804 25483 28806
rect 25507 28804 25563 28806
rect 25267 27770 25323 27772
rect 25347 27770 25403 27772
rect 25427 27770 25483 27772
rect 25507 27770 25563 27772
rect 25267 27718 25313 27770
rect 25313 27718 25323 27770
rect 25347 27718 25377 27770
rect 25377 27718 25389 27770
rect 25389 27718 25403 27770
rect 25427 27718 25441 27770
rect 25441 27718 25453 27770
rect 25453 27718 25483 27770
rect 25507 27718 25517 27770
rect 25517 27718 25563 27770
rect 25267 27716 25323 27718
rect 25347 27716 25403 27718
rect 25427 27716 25483 27718
rect 25507 27716 25563 27718
rect 25267 26682 25323 26684
rect 25347 26682 25403 26684
rect 25427 26682 25483 26684
rect 25507 26682 25563 26684
rect 25267 26630 25313 26682
rect 25313 26630 25323 26682
rect 25347 26630 25377 26682
rect 25377 26630 25389 26682
rect 25389 26630 25403 26682
rect 25427 26630 25441 26682
rect 25441 26630 25453 26682
rect 25453 26630 25483 26682
rect 25507 26630 25517 26682
rect 25517 26630 25563 26682
rect 25267 26628 25323 26630
rect 25347 26628 25403 26630
rect 25427 26628 25483 26630
rect 25507 26628 25563 26630
rect 25267 25594 25323 25596
rect 25347 25594 25403 25596
rect 25427 25594 25483 25596
rect 25507 25594 25563 25596
rect 25267 25542 25313 25594
rect 25313 25542 25323 25594
rect 25347 25542 25377 25594
rect 25377 25542 25389 25594
rect 25389 25542 25403 25594
rect 25427 25542 25441 25594
rect 25441 25542 25453 25594
rect 25453 25542 25483 25594
rect 25507 25542 25517 25594
rect 25517 25542 25563 25594
rect 25267 25540 25323 25542
rect 25347 25540 25403 25542
rect 25427 25540 25483 25542
rect 25507 25540 25563 25542
rect 25267 24506 25323 24508
rect 25347 24506 25403 24508
rect 25427 24506 25483 24508
rect 25507 24506 25563 24508
rect 25267 24454 25313 24506
rect 25313 24454 25323 24506
rect 25347 24454 25377 24506
rect 25377 24454 25389 24506
rect 25389 24454 25403 24506
rect 25427 24454 25441 24506
rect 25441 24454 25453 24506
rect 25453 24454 25483 24506
rect 25507 24454 25517 24506
rect 25517 24454 25563 24506
rect 25267 24452 25323 24454
rect 25347 24452 25403 24454
rect 25427 24452 25483 24454
rect 25507 24452 25563 24454
rect 25267 23418 25323 23420
rect 25347 23418 25403 23420
rect 25427 23418 25483 23420
rect 25507 23418 25563 23420
rect 25267 23366 25313 23418
rect 25313 23366 25323 23418
rect 25347 23366 25377 23418
rect 25377 23366 25389 23418
rect 25389 23366 25403 23418
rect 25427 23366 25441 23418
rect 25441 23366 25453 23418
rect 25453 23366 25483 23418
rect 25507 23366 25517 23418
rect 25517 23366 25563 23418
rect 25267 23364 25323 23366
rect 25347 23364 25403 23366
rect 25427 23364 25483 23366
rect 25507 23364 25563 23366
rect 25267 22330 25323 22332
rect 25347 22330 25403 22332
rect 25427 22330 25483 22332
rect 25507 22330 25563 22332
rect 25267 22278 25313 22330
rect 25313 22278 25323 22330
rect 25347 22278 25377 22330
rect 25377 22278 25389 22330
rect 25389 22278 25403 22330
rect 25427 22278 25441 22330
rect 25441 22278 25453 22330
rect 25453 22278 25483 22330
rect 25507 22278 25517 22330
rect 25517 22278 25563 22330
rect 25267 22276 25323 22278
rect 25347 22276 25403 22278
rect 25427 22276 25483 22278
rect 25507 22276 25563 22278
rect 25267 21242 25323 21244
rect 25347 21242 25403 21244
rect 25427 21242 25483 21244
rect 25507 21242 25563 21244
rect 25267 21190 25313 21242
rect 25313 21190 25323 21242
rect 25347 21190 25377 21242
rect 25377 21190 25389 21242
rect 25389 21190 25403 21242
rect 25427 21190 25441 21242
rect 25441 21190 25453 21242
rect 25453 21190 25483 21242
rect 25507 21190 25517 21242
rect 25517 21190 25563 21242
rect 25267 21188 25323 21190
rect 25347 21188 25403 21190
rect 25427 21188 25483 21190
rect 25507 21188 25563 21190
rect 25267 20154 25323 20156
rect 25347 20154 25403 20156
rect 25427 20154 25483 20156
rect 25507 20154 25563 20156
rect 25267 20102 25313 20154
rect 25313 20102 25323 20154
rect 25347 20102 25377 20154
rect 25377 20102 25389 20154
rect 25389 20102 25403 20154
rect 25427 20102 25441 20154
rect 25441 20102 25453 20154
rect 25453 20102 25483 20154
rect 25507 20102 25517 20154
rect 25517 20102 25563 20154
rect 25267 20100 25323 20102
rect 25347 20100 25403 20102
rect 25427 20100 25483 20102
rect 25507 20100 25563 20102
rect 26146 19760 26202 19816
rect 25267 19066 25323 19068
rect 25347 19066 25403 19068
rect 25427 19066 25483 19068
rect 25507 19066 25563 19068
rect 25267 19014 25313 19066
rect 25313 19014 25323 19066
rect 25347 19014 25377 19066
rect 25377 19014 25389 19066
rect 25389 19014 25403 19066
rect 25427 19014 25441 19066
rect 25441 19014 25453 19066
rect 25453 19014 25483 19066
rect 25507 19014 25517 19066
rect 25517 19014 25563 19066
rect 25267 19012 25323 19014
rect 25347 19012 25403 19014
rect 25427 19012 25483 19014
rect 25507 19012 25563 19014
rect 25267 17978 25323 17980
rect 25347 17978 25403 17980
rect 25427 17978 25483 17980
rect 25507 17978 25563 17980
rect 25267 17926 25313 17978
rect 25313 17926 25323 17978
rect 25347 17926 25377 17978
rect 25377 17926 25389 17978
rect 25389 17926 25403 17978
rect 25427 17926 25441 17978
rect 25441 17926 25453 17978
rect 25453 17926 25483 17978
rect 25507 17926 25517 17978
rect 25517 17926 25563 17978
rect 25267 17924 25323 17926
rect 25347 17924 25403 17926
rect 25427 17924 25483 17926
rect 25507 17924 25563 17926
rect 21794 9818 21850 9820
rect 21874 9818 21930 9820
rect 21954 9818 22010 9820
rect 22034 9818 22090 9820
rect 21794 9766 21840 9818
rect 21840 9766 21850 9818
rect 21874 9766 21904 9818
rect 21904 9766 21916 9818
rect 21916 9766 21930 9818
rect 21954 9766 21968 9818
rect 21968 9766 21980 9818
rect 21980 9766 22010 9818
rect 22034 9766 22044 9818
rect 22044 9766 22090 9818
rect 21794 9764 21850 9766
rect 21874 9764 21930 9766
rect 21954 9764 22010 9766
rect 22034 9764 22090 9766
rect 21794 8730 21850 8732
rect 21874 8730 21930 8732
rect 21954 8730 22010 8732
rect 22034 8730 22090 8732
rect 21794 8678 21840 8730
rect 21840 8678 21850 8730
rect 21874 8678 21904 8730
rect 21904 8678 21916 8730
rect 21916 8678 21930 8730
rect 21954 8678 21968 8730
rect 21968 8678 21980 8730
rect 21980 8678 22010 8730
rect 22034 8678 22044 8730
rect 22044 8678 22090 8730
rect 21794 8676 21850 8678
rect 21874 8676 21930 8678
rect 21954 8676 22010 8678
rect 22034 8676 22090 8678
rect 21794 7642 21850 7644
rect 21874 7642 21930 7644
rect 21954 7642 22010 7644
rect 22034 7642 22090 7644
rect 21794 7590 21840 7642
rect 21840 7590 21850 7642
rect 21874 7590 21904 7642
rect 21904 7590 21916 7642
rect 21916 7590 21930 7642
rect 21954 7590 21968 7642
rect 21968 7590 21980 7642
rect 21980 7590 22010 7642
rect 22034 7590 22044 7642
rect 22044 7590 22090 7642
rect 21794 7588 21850 7590
rect 21874 7588 21930 7590
rect 21954 7588 22010 7590
rect 22034 7588 22090 7590
rect 21794 6554 21850 6556
rect 21874 6554 21930 6556
rect 21954 6554 22010 6556
rect 22034 6554 22090 6556
rect 21794 6502 21840 6554
rect 21840 6502 21850 6554
rect 21874 6502 21904 6554
rect 21904 6502 21916 6554
rect 21916 6502 21930 6554
rect 21954 6502 21968 6554
rect 21968 6502 21980 6554
rect 21980 6502 22010 6554
rect 22034 6502 22044 6554
rect 22044 6502 22090 6554
rect 21794 6500 21850 6502
rect 21874 6500 21930 6502
rect 21954 6500 22010 6502
rect 22034 6500 22090 6502
rect 18321 6010 18377 6012
rect 18401 6010 18457 6012
rect 18481 6010 18537 6012
rect 18561 6010 18617 6012
rect 18321 5958 18367 6010
rect 18367 5958 18377 6010
rect 18401 5958 18431 6010
rect 18431 5958 18443 6010
rect 18443 5958 18457 6010
rect 18481 5958 18495 6010
rect 18495 5958 18507 6010
rect 18507 5958 18537 6010
rect 18561 5958 18571 6010
rect 18571 5958 18617 6010
rect 18321 5956 18377 5958
rect 18401 5956 18457 5958
rect 18481 5956 18537 5958
rect 18561 5956 18617 5958
rect 21794 5466 21850 5468
rect 21874 5466 21930 5468
rect 21954 5466 22010 5468
rect 22034 5466 22090 5468
rect 21794 5414 21840 5466
rect 21840 5414 21850 5466
rect 21874 5414 21904 5466
rect 21904 5414 21916 5466
rect 21916 5414 21930 5466
rect 21954 5414 21968 5466
rect 21968 5414 21980 5466
rect 21980 5414 22010 5466
rect 22034 5414 22044 5466
rect 22044 5414 22090 5466
rect 21794 5412 21850 5414
rect 21874 5412 21930 5414
rect 21954 5412 22010 5414
rect 22034 5412 22090 5414
rect 18321 4922 18377 4924
rect 18401 4922 18457 4924
rect 18481 4922 18537 4924
rect 18561 4922 18617 4924
rect 18321 4870 18367 4922
rect 18367 4870 18377 4922
rect 18401 4870 18431 4922
rect 18431 4870 18443 4922
rect 18443 4870 18457 4922
rect 18481 4870 18495 4922
rect 18495 4870 18507 4922
rect 18507 4870 18537 4922
rect 18561 4870 18571 4922
rect 18571 4870 18617 4922
rect 18321 4868 18377 4870
rect 18401 4868 18457 4870
rect 18481 4868 18537 4870
rect 18561 4868 18617 4870
rect 21794 4378 21850 4380
rect 21874 4378 21930 4380
rect 21954 4378 22010 4380
rect 22034 4378 22090 4380
rect 21794 4326 21840 4378
rect 21840 4326 21850 4378
rect 21874 4326 21904 4378
rect 21904 4326 21916 4378
rect 21916 4326 21930 4378
rect 21954 4326 21968 4378
rect 21968 4326 21980 4378
rect 21980 4326 22010 4378
rect 22034 4326 22044 4378
rect 22044 4326 22090 4378
rect 21794 4324 21850 4326
rect 21874 4324 21930 4326
rect 21954 4324 22010 4326
rect 22034 4324 22090 4326
rect 18321 3834 18377 3836
rect 18401 3834 18457 3836
rect 18481 3834 18537 3836
rect 18561 3834 18617 3836
rect 18321 3782 18367 3834
rect 18367 3782 18377 3834
rect 18401 3782 18431 3834
rect 18431 3782 18443 3834
rect 18443 3782 18457 3834
rect 18481 3782 18495 3834
rect 18495 3782 18507 3834
rect 18507 3782 18537 3834
rect 18561 3782 18571 3834
rect 18571 3782 18617 3834
rect 18321 3780 18377 3782
rect 18401 3780 18457 3782
rect 18481 3780 18537 3782
rect 18561 3780 18617 3782
rect 18321 2746 18377 2748
rect 18401 2746 18457 2748
rect 18481 2746 18537 2748
rect 18561 2746 18617 2748
rect 18321 2694 18367 2746
rect 18367 2694 18377 2746
rect 18401 2694 18431 2746
rect 18431 2694 18443 2746
rect 18443 2694 18457 2746
rect 18481 2694 18495 2746
rect 18495 2694 18507 2746
rect 18507 2694 18537 2746
rect 18561 2694 18571 2746
rect 18571 2694 18617 2746
rect 18321 2692 18377 2694
rect 18401 2692 18457 2694
rect 18481 2692 18537 2694
rect 18561 2692 18617 2694
rect 21794 3290 21850 3292
rect 21874 3290 21930 3292
rect 21954 3290 22010 3292
rect 22034 3290 22090 3292
rect 21794 3238 21840 3290
rect 21840 3238 21850 3290
rect 21874 3238 21904 3290
rect 21904 3238 21916 3290
rect 21916 3238 21930 3290
rect 21954 3238 21968 3290
rect 21968 3238 21980 3290
rect 21980 3238 22010 3290
rect 22034 3238 22044 3290
rect 22044 3238 22090 3290
rect 21794 3236 21850 3238
rect 21874 3236 21930 3238
rect 21954 3236 22010 3238
rect 22034 3236 22090 3238
rect 21794 2202 21850 2204
rect 21874 2202 21930 2204
rect 21954 2202 22010 2204
rect 22034 2202 22090 2204
rect 21794 2150 21840 2202
rect 21840 2150 21850 2202
rect 21874 2150 21904 2202
rect 21904 2150 21916 2202
rect 21916 2150 21930 2202
rect 21954 2150 21968 2202
rect 21968 2150 21980 2202
rect 21980 2150 22010 2202
rect 22034 2150 22044 2202
rect 22044 2150 22090 2202
rect 21794 2148 21850 2150
rect 21874 2148 21930 2150
rect 21954 2148 22010 2150
rect 22034 2148 22090 2150
rect 25267 16890 25323 16892
rect 25347 16890 25403 16892
rect 25427 16890 25483 16892
rect 25507 16890 25563 16892
rect 25267 16838 25313 16890
rect 25313 16838 25323 16890
rect 25347 16838 25377 16890
rect 25377 16838 25389 16890
rect 25389 16838 25403 16890
rect 25427 16838 25441 16890
rect 25441 16838 25453 16890
rect 25453 16838 25483 16890
rect 25507 16838 25517 16890
rect 25517 16838 25563 16890
rect 25267 16836 25323 16838
rect 25347 16836 25403 16838
rect 25427 16836 25483 16838
rect 25507 16836 25563 16838
rect 25267 15802 25323 15804
rect 25347 15802 25403 15804
rect 25427 15802 25483 15804
rect 25507 15802 25563 15804
rect 25267 15750 25313 15802
rect 25313 15750 25323 15802
rect 25347 15750 25377 15802
rect 25377 15750 25389 15802
rect 25389 15750 25403 15802
rect 25427 15750 25441 15802
rect 25441 15750 25453 15802
rect 25453 15750 25483 15802
rect 25507 15750 25517 15802
rect 25517 15750 25563 15802
rect 25267 15748 25323 15750
rect 25347 15748 25403 15750
rect 25427 15748 25483 15750
rect 25507 15748 25563 15750
rect 25267 14714 25323 14716
rect 25347 14714 25403 14716
rect 25427 14714 25483 14716
rect 25507 14714 25563 14716
rect 25267 14662 25313 14714
rect 25313 14662 25323 14714
rect 25347 14662 25377 14714
rect 25377 14662 25389 14714
rect 25389 14662 25403 14714
rect 25427 14662 25441 14714
rect 25441 14662 25453 14714
rect 25453 14662 25483 14714
rect 25507 14662 25517 14714
rect 25517 14662 25563 14714
rect 25267 14660 25323 14662
rect 25347 14660 25403 14662
rect 25427 14660 25483 14662
rect 25507 14660 25563 14662
rect 25267 13626 25323 13628
rect 25347 13626 25403 13628
rect 25427 13626 25483 13628
rect 25507 13626 25563 13628
rect 25267 13574 25313 13626
rect 25313 13574 25323 13626
rect 25347 13574 25377 13626
rect 25377 13574 25389 13626
rect 25389 13574 25403 13626
rect 25427 13574 25441 13626
rect 25441 13574 25453 13626
rect 25453 13574 25483 13626
rect 25507 13574 25517 13626
rect 25517 13574 25563 13626
rect 25267 13572 25323 13574
rect 25347 13572 25403 13574
rect 25427 13572 25483 13574
rect 25507 13572 25563 13574
rect 25267 12538 25323 12540
rect 25347 12538 25403 12540
rect 25427 12538 25483 12540
rect 25507 12538 25563 12540
rect 25267 12486 25313 12538
rect 25313 12486 25323 12538
rect 25347 12486 25377 12538
rect 25377 12486 25389 12538
rect 25389 12486 25403 12538
rect 25427 12486 25441 12538
rect 25441 12486 25453 12538
rect 25453 12486 25483 12538
rect 25507 12486 25517 12538
rect 25517 12486 25563 12538
rect 25267 12484 25323 12486
rect 25347 12484 25403 12486
rect 25427 12484 25483 12486
rect 25507 12484 25563 12486
rect 25267 11450 25323 11452
rect 25347 11450 25403 11452
rect 25427 11450 25483 11452
rect 25507 11450 25563 11452
rect 25267 11398 25313 11450
rect 25313 11398 25323 11450
rect 25347 11398 25377 11450
rect 25377 11398 25389 11450
rect 25389 11398 25403 11450
rect 25427 11398 25441 11450
rect 25441 11398 25453 11450
rect 25453 11398 25483 11450
rect 25507 11398 25517 11450
rect 25517 11398 25563 11450
rect 25267 11396 25323 11398
rect 25347 11396 25403 11398
rect 25427 11396 25483 11398
rect 25507 11396 25563 11398
rect 25267 10362 25323 10364
rect 25347 10362 25403 10364
rect 25427 10362 25483 10364
rect 25507 10362 25563 10364
rect 25267 10310 25313 10362
rect 25313 10310 25323 10362
rect 25347 10310 25377 10362
rect 25377 10310 25389 10362
rect 25389 10310 25403 10362
rect 25427 10310 25441 10362
rect 25441 10310 25453 10362
rect 25453 10310 25483 10362
rect 25507 10310 25517 10362
rect 25517 10310 25563 10362
rect 25267 10308 25323 10310
rect 25347 10308 25403 10310
rect 25427 10308 25483 10310
rect 25507 10308 25563 10310
rect 25267 9274 25323 9276
rect 25347 9274 25403 9276
rect 25427 9274 25483 9276
rect 25507 9274 25563 9276
rect 25267 9222 25313 9274
rect 25313 9222 25323 9274
rect 25347 9222 25377 9274
rect 25377 9222 25389 9274
rect 25389 9222 25403 9274
rect 25427 9222 25441 9274
rect 25441 9222 25453 9274
rect 25453 9222 25483 9274
rect 25507 9222 25517 9274
rect 25517 9222 25563 9274
rect 25267 9220 25323 9222
rect 25347 9220 25403 9222
rect 25427 9220 25483 9222
rect 25507 9220 25563 9222
rect 25267 8186 25323 8188
rect 25347 8186 25403 8188
rect 25427 8186 25483 8188
rect 25507 8186 25563 8188
rect 25267 8134 25313 8186
rect 25313 8134 25323 8186
rect 25347 8134 25377 8186
rect 25377 8134 25389 8186
rect 25389 8134 25403 8186
rect 25427 8134 25441 8186
rect 25441 8134 25453 8186
rect 25453 8134 25483 8186
rect 25507 8134 25517 8186
rect 25517 8134 25563 8186
rect 25267 8132 25323 8134
rect 25347 8132 25403 8134
rect 25427 8132 25483 8134
rect 25507 8132 25563 8134
rect 25267 7098 25323 7100
rect 25347 7098 25403 7100
rect 25427 7098 25483 7100
rect 25507 7098 25563 7100
rect 25267 7046 25313 7098
rect 25313 7046 25323 7098
rect 25347 7046 25377 7098
rect 25377 7046 25389 7098
rect 25389 7046 25403 7098
rect 25427 7046 25441 7098
rect 25441 7046 25453 7098
rect 25453 7046 25483 7098
rect 25507 7046 25517 7098
rect 25517 7046 25563 7098
rect 25267 7044 25323 7046
rect 25347 7044 25403 7046
rect 25427 7044 25483 7046
rect 25507 7044 25563 7046
rect 25267 6010 25323 6012
rect 25347 6010 25403 6012
rect 25427 6010 25483 6012
rect 25507 6010 25563 6012
rect 25267 5958 25313 6010
rect 25313 5958 25323 6010
rect 25347 5958 25377 6010
rect 25377 5958 25389 6010
rect 25389 5958 25403 6010
rect 25427 5958 25441 6010
rect 25441 5958 25453 6010
rect 25453 5958 25483 6010
rect 25507 5958 25517 6010
rect 25517 5958 25563 6010
rect 25267 5956 25323 5958
rect 25347 5956 25403 5958
rect 25427 5956 25483 5958
rect 25507 5956 25563 5958
rect 25267 4922 25323 4924
rect 25347 4922 25403 4924
rect 25427 4922 25483 4924
rect 25507 4922 25563 4924
rect 25267 4870 25313 4922
rect 25313 4870 25323 4922
rect 25347 4870 25377 4922
rect 25377 4870 25389 4922
rect 25389 4870 25403 4922
rect 25427 4870 25441 4922
rect 25441 4870 25453 4922
rect 25453 4870 25483 4922
rect 25507 4870 25517 4922
rect 25517 4870 25563 4922
rect 25267 4868 25323 4870
rect 25347 4868 25403 4870
rect 25427 4868 25483 4870
rect 25507 4868 25563 4870
rect 25267 3834 25323 3836
rect 25347 3834 25403 3836
rect 25427 3834 25483 3836
rect 25507 3834 25563 3836
rect 25267 3782 25313 3834
rect 25313 3782 25323 3834
rect 25347 3782 25377 3834
rect 25377 3782 25389 3834
rect 25389 3782 25403 3834
rect 25427 3782 25441 3834
rect 25441 3782 25453 3834
rect 25453 3782 25483 3834
rect 25507 3782 25517 3834
rect 25517 3782 25563 3834
rect 25267 3780 25323 3782
rect 25347 3780 25403 3782
rect 25427 3780 25483 3782
rect 25507 3780 25563 3782
rect 25267 2746 25323 2748
rect 25347 2746 25403 2748
rect 25427 2746 25483 2748
rect 25507 2746 25563 2748
rect 25267 2694 25313 2746
rect 25313 2694 25323 2746
rect 25347 2694 25377 2746
rect 25377 2694 25389 2746
rect 25389 2694 25403 2746
rect 25427 2694 25441 2746
rect 25441 2694 25453 2746
rect 25453 2694 25483 2746
rect 25507 2694 25517 2746
rect 25517 2694 25563 2746
rect 25267 2692 25323 2694
rect 25347 2692 25403 2694
rect 25427 2692 25483 2694
rect 25507 2692 25563 2694
rect 27526 34060 27582 34096
rect 27526 34040 27528 34060
rect 27528 34040 27580 34060
rect 27580 34040 27582 34060
rect 27526 32972 27582 33008
rect 27526 32952 27528 32972
rect 27528 32952 27580 32972
rect 27580 32952 27582 32972
rect 26146 8200 26202 8256
rect 26146 6840 26202 6896
rect 27526 31320 27582 31376
rect 28354 36760 28410 36816
rect 28354 36116 28356 36136
rect 28356 36116 28408 36136
rect 28408 36116 28410 36136
rect 28354 36080 28410 36116
rect 27526 28600 27582 28656
rect 27526 27532 27582 27568
rect 27526 27512 27528 27532
rect 27528 27512 27580 27532
rect 27580 27512 27582 27532
rect 27434 26560 27490 26616
rect 28262 32000 28318 32056
rect 27526 21936 27582 21992
rect 27342 16532 27344 16552
rect 27344 16532 27396 16552
rect 27396 16532 27398 16552
rect 27342 16496 27398 16532
rect 28740 45722 28796 45724
rect 28820 45722 28876 45724
rect 28900 45722 28956 45724
rect 28980 45722 29036 45724
rect 28740 45670 28786 45722
rect 28786 45670 28796 45722
rect 28820 45670 28850 45722
rect 28850 45670 28862 45722
rect 28862 45670 28876 45722
rect 28900 45670 28914 45722
rect 28914 45670 28926 45722
rect 28926 45670 28956 45722
rect 28980 45670 28990 45722
rect 28990 45670 29036 45722
rect 28740 45668 28796 45670
rect 28820 45668 28876 45670
rect 28900 45668 28956 45670
rect 28980 45668 29036 45670
rect 28740 44634 28796 44636
rect 28820 44634 28876 44636
rect 28900 44634 28956 44636
rect 28980 44634 29036 44636
rect 28740 44582 28786 44634
rect 28786 44582 28796 44634
rect 28820 44582 28850 44634
rect 28850 44582 28862 44634
rect 28862 44582 28876 44634
rect 28900 44582 28914 44634
rect 28914 44582 28926 44634
rect 28926 44582 28956 44634
rect 28980 44582 28990 44634
rect 28990 44582 29036 44634
rect 28740 44580 28796 44582
rect 28820 44580 28876 44582
rect 28900 44580 28956 44582
rect 28980 44580 29036 44582
rect 28740 43546 28796 43548
rect 28820 43546 28876 43548
rect 28900 43546 28956 43548
rect 28980 43546 29036 43548
rect 28740 43494 28786 43546
rect 28786 43494 28796 43546
rect 28820 43494 28850 43546
rect 28850 43494 28862 43546
rect 28862 43494 28876 43546
rect 28900 43494 28914 43546
rect 28914 43494 28926 43546
rect 28926 43494 28956 43546
rect 28980 43494 28990 43546
rect 28990 43494 29036 43546
rect 28740 43492 28796 43494
rect 28820 43492 28876 43494
rect 28900 43492 28956 43494
rect 28980 43492 29036 43494
rect 28740 42458 28796 42460
rect 28820 42458 28876 42460
rect 28900 42458 28956 42460
rect 28980 42458 29036 42460
rect 28740 42406 28786 42458
rect 28786 42406 28796 42458
rect 28820 42406 28850 42458
rect 28850 42406 28862 42458
rect 28862 42406 28876 42458
rect 28900 42406 28914 42458
rect 28914 42406 28926 42458
rect 28926 42406 28956 42458
rect 28980 42406 28990 42458
rect 28990 42406 29036 42458
rect 28740 42404 28796 42406
rect 28820 42404 28876 42406
rect 28900 42404 28956 42406
rect 28980 42404 29036 42406
rect 28740 41370 28796 41372
rect 28820 41370 28876 41372
rect 28900 41370 28956 41372
rect 28980 41370 29036 41372
rect 28740 41318 28786 41370
rect 28786 41318 28796 41370
rect 28820 41318 28850 41370
rect 28850 41318 28862 41370
rect 28862 41318 28876 41370
rect 28900 41318 28914 41370
rect 28914 41318 28926 41370
rect 28926 41318 28956 41370
rect 28980 41318 28990 41370
rect 28990 41318 29036 41370
rect 28740 41316 28796 41318
rect 28820 41316 28876 41318
rect 28900 41316 28956 41318
rect 28980 41316 29036 41318
rect 28630 40840 28686 40896
rect 28740 40282 28796 40284
rect 28820 40282 28876 40284
rect 28900 40282 28956 40284
rect 28980 40282 29036 40284
rect 28740 40230 28786 40282
rect 28786 40230 28796 40282
rect 28820 40230 28850 40282
rect 28850 40230 28862 40282
rect 28862 40230 28876 40282
rect 28900 40230 28914 40282
rect 28914 40230 28926 40282
rect 28926 40230 28956 40282
rect 28980 40230 28990 40282
rect 28990 40230 29036 40282
rect 28740 40228 28796 40230
rect 28820 40228 28876 40230
rect 28900 40228 28956 40230
rect 28980 40228 29036 40230
rect 28740 39194 28796 39196
rect 28820 39194 28876 39196
rect 28900 39194 28956 39196
rect 28980 39194 29036 39196
rect 28740 39142 28786 39194
rect 28786 39142 28796 39194
rect 28820 39142 28850 39194
rect 28850 39142 28862 39194
rect 28862 39142 28876 39194
rect 28900 39142 28914 39194
rect 28914 39142 28926 39194
rect 28926 39142 28956 39194
rect 28980 39142 28990 39194
rect 28990 39142 29036 39194
rect 28740 39140 28796 39142
rect 28820 39140 28876 39142
rect 28900 39140 28956 39142
rect 28980 39140 29036 39142
rect 28354 29960 28410 30016
rect 27526 15680 27582 15736
rect 27526 10240 27582 10296
rect 27526 8880 27582 8936
rect 27434 3440 27490 3496
rect 26146 2760 26202 2816
rect 28354 25220 28410 25256
rect 28354 25200 28356 25220
rect 28356 25200 28408 25220
rect 28408 25200 28410 25220
rect 28354 24520 28410 24576
rect 28354 21120 28410 21176
rect 28354 20440 28410 20496
rect 28446 15000 28502 15056
rect 28354 14356 28356 14376
rect 28356 14356 28408 14376
rect 28408 14356 28410 14376
rect 28354 14320 28410 14356
rect 28354 12300 28410 12336
rect 28354 12280 28356 12300
rect 28356 12280 28408 12300
rect 28408 12280 28410 12300
rect 28740 38106 28796 38108
rect 28820 38106 28876 38108
rect 28900 38106 28956 38108
rect 28980 38106 29036 38108
rect 28740 38054 28786 38106
rect 28786 38054 28796 38106
rect 28820 38054 28850 38106
rect 28850 38054 28862 38106
rect 28862 38054 28876 38106
rect 28900 38054 28914 38106
rect 28914 38054 28926 38106
rect 28926 38054 28956 38106
rect 28980 38054 28990 38106
rect 28990 38054 29036 38106
rect 28740 38052 28796 38054
rect 28820 38052 28876 38054
rect 28900 38052 28956 38054
rect 28980 38052 29036 38054
rect 28740 37018 28796 37020
rect 28820 37018 28876 37020
rect 28900 37018 28956 37020
rect 28980 37018 29036 37020
rect 28740 36966 28786 37018
rect 28786 36966 28796 37018
rect 28820 36966 28850 37018
rect 28850 36966 28862 37018
rect 28862 36966 28876 37018
rect 28900 36966 28914 37018
rect 28914 36966 28926 37018
rect 28926 36966 28956 37018
rect 28980 36966 28990 37018
rect 28990 36966 29036 37018
rect 28740 36964 28796 36966
rect 28820 36964 28876 36966
rect 28900 36964 28956 36966
rect 28980 36964 29036 36966
rect 28740 35930 28796 35932
rect 28820 35930 28876 35932
rect 28900 35930 28956 35932
rect 28980 35930 29036 35932
rect 28740 35878 28786 35930
rect 28786 35878 28796 35930
rect 28820 35878 28850 35930
rect 28850 35878 28862 35930
rect 28862 35878 28876 35930
rect 28900 35878 28914 35930
rect 28914 35878 28926 35930
rect 28926 35878 28956 35930
rect 28980 35878 28990 35930
rect 28990 35878 29036 35930
rect 28740 35876 28796 35878
rect 28820 35876 28876 35878
rect 28900 35876 28956 35878
rect 28980 35876 29036 35878
rect 28740 34842 28796 34844
rect 28820 34842 28876 34844
rect 28900 34842 28956 34844
rect 28980 34842 29036 34844
rect 28740 34790 28786 34842
rect 28786 34790 28796 34842
rect 28820 34790 28850 34842
rect 28850 34790 28862 34842
rect 28862 34790 28876 34842
rect 28900 34790 28914 34842
rect 28914 34790 28926 34842
rect 28926 34790 28956 34842
rect 28980 34790 28990 34842
rect 28990 34790 29036 34842
rect 28740 34788 28796 34790
rect 28820 34788 28876 34790
rect 28900 34788 28956 34790
rect 28980 34788 29036 34790
rect 28740 33754 28796 33756
rect 28820 33754 28876 33756
rect 28900 33754 28956 33756
rect 28980 33754 29036 33756
rect 28740 33702 28786 33754
rect 28786 33702 28796 33754
rect 28820 33702 28850 33754
rect 28850 33702 28862 33754
rect 28862 33702 28876 33754
rect 28900 33702 28914 33754
rect 28914 33702 28926 33754
rect 28926 33702 28956 33754
rect 28980 33702 28990 33754
rect 28990 33702 29036 33754
rect 28740 33700 28796 33702
rect 28820 33700 28876 33702
rect 28900 33700 28956 33702
rect 28980 33700 29036 33702
rect 28740 32666 28796 32668
rect 28820 32666 28876 32668
rect 28900 32666 28956 32668
rect 28980 32666 29036 32668
rect 28740 32614 28786 32666
rect 28786 32614 28796 32666
rect 28820 32614 28850 32666
rect 28850 32614 28862 32666
rect 28862 32614 28876 32666
rect 28900 32614 28914 32666
rect 28914 32614 28926 32666
rect 28926 32614 28956 32666
rect 28980 32614 28990 32666
rect 28990 32614 29036 32666
rect 28740 32612 28796 32614
rect 28820 32612 28876 32614
rect 28900 32612 28956 32614
rect 28980 32612 29036 32614
rect 28740 31578 28796 31580
rect 28820 31578 28876 31580
rect 28900 31578 28956 31580
rect 28980 31578 29036 31580
rect 28740 31526 28786 31578
rect 28786 31526 28796 31578
rect 28820 31526 28850 31578
rect 28850 31526 28862 31578
rect 28862 31526 28876 31578
rect 28900 31526 28914 31578
rect 28914 31526 28926 31578
rect 28926 31526 28956 31578
rect 28980 31526 28990 31578
rect 28990 31526 29036 31578
rect 28740 31524 28796 31526
rect 28820 31524 28876 31526
rect 28900 31524 28956 31526
rect 28980 31524 29036 31526
rect 28740 30490 28796 30492
rect 28820 30490 28876 30492
rect 28900 30490 28956 30492
rect 28980 30490 29036 30492
rect 28740 30438 28786 30490
rect 28786 30438 28796 30490
rect 28820 30438 28850 30490
rect 28850 30438 28862 30490
rect 28862 30438 28876 30490
rect 28900 30438 28914 30490
rect 28914 30438 28926 30490
rect 28926 30438 28956 30490
rect 28980 30438 28990 30490
rect 28990 30438 29036 30490
rect 28740 30436 28796 30438
rect 28820 30436 28876 30438
rect 28900 30436 28956 30438
rect 28980 30436 29036 30438
rect 28740 29402 28796 29404
rect 28820 29402 28876 29404
rect 28900 29402 28956 29404
rect 28980 29402 29036 29404
rect 28740 29350 28786 29402
rect 28786 29350 28796 29402
rect 28820 29350 28850 29402
rect 28850 29350 28862 29402
rect 28862 29350 28876 29402
rect 28900 29350 28914 29402
rect 28914 29350 28926 29402
rect 28926 29350 28956 29402
rect 28980 29350 28990 29402
rect 28990 29350 29036 29402
rect 28740 29348 28796 29350
rect 28820 29348 28876 29350
rect 28900 29348 28956 29350
rect 28980 29348 29036 29350
rect 28740 28314 28796 28316
rect 28820 28314 28876 28316
rect 28900 28314 28956 28316
rect 28980 28314 29036 28316
rect 28740 28262 28786 28314
rect 28786 28262 28796 28314
rect 28820 28262 28850 28314
rect 28850 28262 28862 28314
rect 28862 28262 28876 28314
rect 28900 28262 28914 28314
rect 28914 28262 28926 28314
rect 28926 28262 28956 28314
rect 28980 28262 28990 28314
rect 28990 28262 29036 28314
rect 28740 28260 28796 28262
rect 28820 28260 28876 28262
rect 28900 28260 28956 28262
rect 28980 28260 29036 28262
rect 28740 27226 28796 27228
rect 28820 27226 28876 27228
rect 28900 27226 28956 27228
rect 28980 27226 29036 27228
rect 28740 27174 28786 27226
rect 28786 27174 28796 27226
rect 28820 27174 28850 27226
rect 28850 27174 28862 27226
rect 28862 27174 28876 27226
rect 28900 27174 28914 27226
rect 28914 27174 28926 27226
rect 28926 27174 28956 27226
rect 28980 27174 28990 27226
rect 28990 27174 29036 27226
rect 28740 27172 28796 27174
rect 28820 27172 28876 27174
rect 28900 27172 28956 27174
rect 28980 27172 29036 27174
rect 28740 26138 28796 26140
rect 28820 26138 28876 26140
rect 28900 26138 28956 26140
rect 28980 26138 29036 26140
rect 28740 26086 28786 26138
rect 28786 26086 28796 26138
rect 28820 26086 28850 26138
rect 28850 26086 28862 26138
rect 28862 26086 28876 26138
rect 28900 26086 28914 26138
rect 28914 26086 28926 26138
rect 28926 26086 28956 26138
rect 28980 26086 28990 26138
rect 28990 26086 29036 26138
rect 28740 26084 28796 26086
rect 28820 26084 28876 26086
rect 28900 26084 28956 26086
rect 28980 26084 29036 26086
rect 28740 25050 28796 25052
rect 28820 25050 28876 25052
rect 28900 25050 28956 25052
rect 28980 25050 29036 25052
rect 28740 24998 28786 25050
rect 28786 24998 28796 25050
rect 28820 24998 28850 25050
rect 28850 24998 28862 25050
rect 28862 24998 28876 25050
rect 28900 24998 28914 25050
rect 28914 24998 28926 25050
rect 28926 24998 28956 25050
rect 28980 24998 28990 25050
rect 28990 24998 29036 25050
rect 28740 24996 28796 24998
rect 28820 24996 28876 24998
rect 28900 24996 28956 24998
rect 28980 24996 29036 24998
rect 28740 23962 28796 23964
rect 28820 23962 28876 23964
rect 28900 23962 28956 23964
rect 28980 23962 29036 23964
rect 28740 23910 28786 23962
rect 28786 23910 28796 23962
rect 28820 23910 28850 23962
rect 28850 23910 28862 23962
rect 28862 23910 28876 23962
rect 28900 23910 28914 23962
rect 28914 23910 28926 23962
rect 28926 23910 28956 23962
rect 28980 23910 28990 23962
rect 28990 23910 29036 23962
rect 28740 23908 28796 23910
rect 28820 23908 28876 23910
rect 28900 23908 28956 23910
rect 28980 23908 29036 23910
rect 29918 23840 29974 23896
rect 28740 22874 28796 22876
rect 28820 22874 28876 22876
rect 28900 22874 28956 22876
rect 28980 22874 29036 22876
rect 28740 22822 28786 22874
rect 28786 22822 28796 22874
rect 28820 22822 28850 22874
rect 28850 22822 28862 22874
rect 28862 22822 28876 22874
rect 28900 22822 28914 22874
rect 28914 22822 28926 22874
rect 28926 22822 28956 22874
rect 28980 22822 28990 22874
rect 28990 22822 29036 22874
rect 28740 22820 28796 22822
rect 28820 22820 28876 22822
rect 28900 22820 28956 22822
rect 28980 22820 29036 22822
rect 28740 21786 28796 21788
rect 28820 21786 28876 21788
rect 28900 21786 28956 21788
rect 28980 21786 29036 21788
rect 28740 21734 28786 21786
rect 28786 21734 28796 21786
rect 28820 21734 28850 21786
rect 28850 21734 28862 21786
rect 28862 21734 28876 21786
rect 28900 21734 28914 21786
rect 28914 21734 28926 21786
rect 28926 21734 28956 21786
rect 28980 21734 28990 21786
rect 28990 21734 29036 21786
rect 28740 21732 28796 21734
rect 28820 21732 28876 21734
rect 28900 21732 28956 21734
rect 28980 21732 29036 21734
rect 28740 20698 28796 20700
rect 28820 20698 28876 20700
rect 28900 20698 28956 20700
rect 28980 20698 29036 20700
rect 28740 20646 28786 20698
rect 28786 20646 28796 20698
rect 28820 20646 28850 20698
rect 28850 20646 28862 20698
rect 28862 20646 28876 20698
rect 28900 20646 28914 20698
rect 28914 20646 28926 20698
rect 28926 20646 28956 20698
rect 28980 20646 28990 20698
rect 28990 20646 29036 20698
rect 28740 20644 28796 20646
rect 28820 20644 28876 20646
rect 28900 20644 28956 20646
rect 28980 20644 29036 20646
rect 28740 19610 28796 19612
rect 28820 19610 28876 19612
rect 28900 19610 28956 19612
rect 28980 19610 29036 19612
rect 28740 19558 28786 19610
rect 28786 19558 28796 19610
rect 28820 19558 28850 19610
rect 28850 19558 28862 19610
rect 28862 19558 28876 19610
rect 28900 19558 28914 19610
rect 28914 19558 28926 19610
rect 28926 19558 28956 19610
rect 28980 19558 28990 19610
rect 28990 19558 29036 19610
rect 28740 19556 28796 19558
rect 28820 19556 28876 19558
rect 28900 19556 28956 19558
rect 28980 19556 29036 19558
rect 28740 18522 28796 18524
rect 28820 18522 28876 18524
rect 28900 18522 28956 18524
rect 28980 18522 29036 18524
rect 28740 18470 28786 18522
rect 28786 18470 28796 18522
rect 28820 18470 28850 18522
rect 28850 18470 28862 18522
rect 28862 18470 28876 18522
rect 28900 18470 28914 18522
rect 28914 18470 28926 18522
rect 28926 18470 28956 18522
rect 28980 18470 28990 18522
rect 28990 18470 29036 18522
rect 28740 18468 28796 18470
rect 28820 18468 28876 18470
rect 28900 18468 28956 18470
rect 28980 18468 29036 18470
rect 28740 17434 28796 17436
rect 28820 17434 28876 17436
rect 28900 17434 28956 17436
rect 28980 17434 29036 17436
rect 28740 17382 28786 17434
rect 28786 17382 28796 17434
rect 28820 17382 28850 17434
rect 28850 17382 28862 17434
rect 28862 17382 28876 17434
rect 28900 17382 28914 17434
rect 28914 17382 28926 17434
rect 28926 17382 28956 17434
rect 28980 17382 28990 17434
rect 28990 17382 29036 17434
rect 28740 17380 28796 17382
rect 28820 17380 28876 17382
rect 28900 17380 28956 17382
rect 28980 17380 29036 17382
rect 28740 16346 28796 16348
rect 28820 16346 28876 16348
rect 28900 16346 28956 16348
rect 28980 16346 29036 16348
rect 28740 16294 28786 16346
rect 28786 16294 28796 16346
rect 28820 16294 28850 16346
rect 28850 16294 28862 16346
rect 28862 16294 28876 16346
rect 28900 16294 28914 16346
rect 28914 16294 28926 16346
rect 28926 16294 28956 16346
rect 28980 16294 28990 16346
rect 28990 16294 29036 16346
rect 28740 16292 28796 16294
rect 28820 16292 28876 16294
rect 28900 16292 28956 16294
rect 28980 16292 29036 16294
rect 28740 15258 28796 15260
rect 28820 15258 28876 15260
rect 28900 15258 28956 15260
rect 28980 15258 29036 15260
rect 28740 15206 28786 15258
rect 28786 15206 28796 15258
rect 28820 15206 28850 15258
rect 28850 15206 28862 15258
rect 28862 15206 28876 15258
rect 28900 15206 28914 15258
rect 28914 15206 28926 15258
rect 28926 15206 28956 15258
rect 28980 15206 28990 15258
rect 28990 15206 29036 15258
rect 28740 15204 28796 15206
rect 28820 15204 28876 15206
rect 28900 15204 28956 15206
rect 28980 15204 29036 15206
rect 28740 14170 28796 14172
rect 28820 14170 28876 14172
rect 28900 14170 28956 14172
rect 28980 14170 29036 14172
rect 28740 14118 28786 14170
rect 28786 14118 28796 14170
rect 28820 14118 28850 14170
rect 28850 14118 28862 14170
rect 28862 14118 28876 14170
rect 28900 14118 28914 14170
rect 28914 14118 28926 14170
rect 28926 14118 28956 14170
rect 28980 14118 28990 14170
rect 28990 14118 29036 14170
rect 28740 14116 28796 14118
rect 28820 14116 28876 14118
rect 28900 14116 28956 14118
rect 28980 14116 29036 14118
rect 28740 13082 28796 13084
rect 28820 13082 28876 13084
rect 28900 13082 28956 13084
rect 28980 13082 29036 13084
rect 28740 13030 28786 13082
rect 28786 13030 28796 13082
rect 28820 13030 28850 13082
rect 28850 13030 28862 13082
rect 28862 13030 28876 13082
rect 28900 13030 28914 13082
rect 28914 13030 28926 13082
rect 28926 13030 28956 13082
rect 28980 13030 28990 13082
rect 28990 13030 29036 13082
rect 28740 13028 28796 13030
rect 28820 13028 28876 13030
rect 28900 13028 28956 13030
rect 28980 13028 29036 13030
rect 28740 11994 28796 11996
rect 28820 11994 28876 11996
rect 28900 11994 28956 11996
rect 28980 11994 29036 11996
rect 28740 11942 28786 11994
rect 28786 11942 28796 11994
rect 28820 11942 28850 11994
rect 28850 11942 28862 11994
rect 28862 11942 28876 11994
rect 28900 11942 28914 11994
rect 28914 11942 28926 11994
rect 28926 11942 28956 11994
rect 28980 11942 28990 11994
rect 28990 11942 29036 11994
rect 28740 11940 28796 11942
rect 28820 11940 28876 11942
rect 28900 11940 28956 11942
rect 28980 11940 29036 11942
rect 29918 10920 29974 10976
rect 28740 10906 28796 10908
rect 28820 10906 28876 10908
rect 28900 10906 28956 10908
rect 28980 10906 29036 10908
rect 28740 10854 28786 10906
rect 28786 10854 28796 10906
rect 28820 10854 28850 10906
rect 28850 10854 28862 10906
rect 28862 10854 28876 10906
rect 28900 10854 28914 10906
rect 28914 10854 28926 10906
rect 28926 10854 28956 10906
rect 28980 10854 28990 10906
rect 28990 10854 29036 10906
rect 28740 10852 28796 10854
rect 28820 10852 28876 10854
rect 28900 10852 28956 10854
rect 28980 10852 29036 10854
rect 28740 9818 28796 9820
rect 28820 9818 28876 9820
rect 28900 9818 28956 9820
rect 28980 9818 29036 9820
rect 28740 9766 28786 9818
rect 28786 9766 28796 9818
rect 28820 9766 28850 9818
rect 28850 9766 28862 9818
rect 28862 9766 28876 9818
rect 28900 9766 28914 9818
rect 28914 9766 28926 9818
rect 28926 9766 28956 9818
rect 28980 9766 28990 9818
rect 28990 9766 29036 9818
rect 28740 9764 28796 9766
rect 28820 9764 28876 9766
rect 28900 9764 28956 9766
rect 28980 9764 29036 9766
rect 28740 8730 28796 8732
rect 28820 8730 28876 8732
rect 28900 8730 28956 8732
rect 28980 8730 29036 8732
rect 28740 8678 28786 8730
rect 28786 8678 28796 8730
rect 28820 8678 28850 8730
rect 28850 8678 28862 8730
rect 28862 8678 28876 8730
rect 28900 8678 28914 8730
rect 28914 8678 28926 8730
rect 28926 8678 28956 8730
rect 28980 8678 28990 8730
rect 28990 8678 29036 8730
rect 28740 8676 28796 8678
rect 28820 8676 28876 8678
rect 28900 8676 28956 8678
rect 28980 8676 29036 8678
rect 28740 7642 28796 7644
rect 28820 7642 28876 7644
rect 28900 7642 28956 7644
rect 28980 7642 29036 7644
rect 28740 7590 28786 7642
rect 28786 7590 28796 7642
rect 28820 7590 28850 7642
rect 28850 7590 28862 7642
rect 28862 7590 28876 7642
rect 28900 7590 28914 7642
rect 28914 7590 28926 7642
rect 28926 7590 28956 7642
rect 28980 7590 28990 7642
rect 28990 7590 29036 7642
rect 28740 7588 28796 7590
rect 28820 7588 28876 7590
rect 28900 7588 28956 7590
rect 28980 7588 29036 7590
rect 29918 7520 29974 7576
rect 28740 6554 28796 6556
rect 28820 6554 28876 6556
rect 28900 6554 28956 6556
rect 28980 6554 29036 6556
rect 28740 6502 28786 6554
rect 28786 6502 28796 6554
rect 28820 6502 28850 6554
rect 28850 6502 28862 6554
rect 28862 6502 28876 6554
rect 28900 6502 28914 6554
rect 28914 6502 28926 6554
rect 28926 6502 28956 6554
rect 28980 6502 28990 6554
rect 28990 6502 29036 6554
rect 28740 6500 28796 6502
rect 28820 6500 28876 6502
rect 28900 6500 28956 6502
rect 28980 6500 29036 6502
rect 29918 5480 29974 5536
rect 28740 5466 28796 5468
rect 28820 5466 28876 5468
rect 28900 5466 28956 5468
rect 28980 5466 29036 5468
rect 28740 5414 28786 5466
rect 28786 5414 28796 5466
rect 28820 5414 28850 5466
rect 28850 5414 28862 5466
rect 28862 5414 28876 5466
rect 28900 5414 28914 5466
rect 28914 5414 28926 5466
rect 28926 5414 28956 5466
rect 28980 5414 28990 5466
rect 28990 5414 29036 5466
rect 28740 5412 28796 5414
rect 28820 5412 28876 5414
rect 28900 5412 28956 5414
rect 28980 5412 29036 5414
rect 28740 4378 28796 4380
rect 28820 4378 28876 4380
rect 28900 4378 28956 4380
rect 28980 4378 29036 4380
rect 28740 4326 28786 4378
rect 28786 4326 28796 4378
rect 28820 4326 28850 4378
rect 28850 4326 28862 4378
rect 28862 4326 28876 4378
rect 28900 4326 28914 4378
rect 28914 4326 28926 4378
rect 28926 4326 28956 4378
rect 28980 4326 28990 4378
rect 28990 4326 29036 4378
rect 28740 4324 28796 4326
rect 28820 4324 28876 4326
rect 28900 4324 28956 4326
rect 28980 4324 29036 4326
rect 28740 3290 28796 3292
rect 28820 3290 28876 3292
rect 28900 3290 28956 3292
rect 28980 3290 29036 3292
rect 28740 3238 28786 3290
rect 28786 3238 28796 3290
rect 28820 3238 28850 3290
rect 28850 3238 28862 3290
rect 28862 3238 28876 3290
rect 28900 3238 28914 3290
rect 28914 3238 28926 3290
rect 28926 3238 28956 3290
rect 28980 3238 28990 3290
rect 28990 3238 29036 3290
rect 28740 3236 28796 3238
rect 28820 3236 28876 3238
rect 28900 3236 28956 3238
rect 28980 3236 29036 3238
rect 28078 2488 28134 2544
rect 28740 2202 28796 2204
rect 28820 2202 28876 2204
rect 28900 2202 28956 2204
rect 28980 2202 29036 2204
rect 28740 2150 28786 2202
rect 28786 2150 28796 2202
rect 28820 2150 28850 2202
rect 28850 2150 28862 2202
rect 28862 2150 28876 2202
rect 28900 2150 28914 2202
rect 28914 2150 28926 2202
rect 28926 2150 28956 2202
rect 28980 2150 28990 2202
rect 28990 2150 29036 2202
rect 28740 2148 28796 2150
rect 28820 2148 28876 2150
rect 28900 2148 28956 2150
rect 28980 2148 29036 2150
rect 27526 1400 27582 1456
<< metal3 >>
rect 200 49738 800 49828
rect 3509 49738 3575 49741
rect 200 49736 3575 49738
rect 200 49680 3514 49736
rect 3570 49680 3575 49736
rect 200 49678 3575 49680
rect 200 49588 800 49678
rect 3509 49675 3575 49678
rect 26141 49058 26207 49061
rect 29200 49058 29800 49148
rect 26141 49056 29800 49058
rect 26141 49000 26146 49056
rect 26202 49000 29800 49056
rect 26141 48998 29800 49000
rect 26141 48995 26207 48998
rect 29200 48908 29800 48998
rect 200 48228 800 48468
rect 29200 48228 29800 48468
rect 200 47548 800 47788
rect 28257 47698 28323 47701
rect 29200 47698 29800 47788
rect 28257 47696 29800 47698
rect 28257 47640 28262 47696
rect 28318 47640 29800 47696
rect 28257 47638 29800 47640
rect 28257 47635 28323 47638
rect 29200 47548 29800 47638
rect 4419 47360 4735 47361
rect 4419 47296 4425 47360
rect 4489 47296 4505 47360
rect 4569 47296 4585 47360
rect 4649 47296 4665 47360
rect 4729 47296 4735 47360
rect 4419 47295 4735 47296
rect 11365 47360 11681 47361
rect 11365 47296 11371 47360
rect 11435 47296 11451 47360
rect 11515 47296 11531 47360
rect 11595 47296 11611 47360
rect 11675 47296 11681 47360
rect 11365 47295 11681 47296
rect 18311 47360 18627 47361
rect 18311 47296 18317 47360
rect 18381 47296 18397 47360
rect 18461 47296 18477 47360
rect 18541 47296 18557 47360
rect 18621 47296 18627 47360
rect 18311 47295 18627 47296
rect 25257 47360 25573 47361
rect 25257 47296 25263 47360
rect 25327 47296 25343 47360
rect 25407 47296 25423 47360
rect 25487 47296 25503 47360
rect 25567 47296 25573 47360
rect 25257 47295 25573 47296
rect 200 46868 800 47108
rect 26049 47018 26115 47021
rect 29200 47018 29800 47108
rect 26049 47016 29800 47018
rect 26049 46960 26054 47016
rect 26110 46960 29800 47016
rect 26049 46958 29800 46960
rect 26049 46955 26115 46958
rect 29200 46868 29800 46958
rect 7892 46816 8208 46817
rect 7892 46752 7898 46816
rect 7962 46752 7978 46816
rect 8042 46752 8058 46816
rect 8122 46752 8138 46816
rect 8202 46752 8208 46816
rect 7892 46751 8208 46752
rect 14838 46816 15154 46817
rect 14838 46752 14844 46816
rect 14908 46752 14924 46816
rect 14988 46752 15004 46816
rect 15068 46752 15084 46816
rect 15148 46752 15154 46816
rect 14838 46751 15154 46752
rect 21784 46816 22100 46817
rect 21784 46752 21790 46816
rect 21854 46752 21870 46816
rect 21934 46752 21950 46816
rect 22014 46752 22030 46816
rect 22094 46752 22100 46816
rect 21784 46751 22100 46752
rect 28730 46816 29046 46817
rect 28730 46752 28736 46816
rect 28800 46752 28816 46816
rect 28880 46752 28896 46816
rect 28960 46752 28976 46816
rect 29040 46752 29046 46816
rect 28730 46751 29046 46752
rect 200 46188 800 46428
rect 27521 46338 27587 46341
rect 29200 46338 29800 46428
rect 27521 46336 29800 46338
rect 27521 46280 27526 46336
rect 27582 46280 29800 46336
rect 27521 46278 29800 46280
rect 27521 46275 27587 46278
rect 4419 46272 4735 46273
rect 4419 46208 4425 46272
rect 4489 46208 4505 46272
rect 4569 46208 4585 46272
rect 4649 46208 4665 46272
rect 4729 46208 4735 46272
rect 4419 46207 4735 46208
rect 11365 46272 11681 46273
rect 11365 46208 11371 46272
rect 11435 46208 11451 46272
rect 11515 46208 11531 46272
rect 11595 46208 11611 46272
rect 11675 46208 11681 46272
rect 11365 46207 11681 46208
rect 18311 46272 18627 46273
rect 18311 46208 18317 46272
rect 18381 46208 18397 46272
rect 18461 46208 18477 46272
rect 18541 46208 18557 46272
rect 18621 46208 18627 46272
rect 18311 46207 18627 46208
rect 25257 46272 25573 46273
rect 25257 46208 25263 46272
rect 25327 46208 25343 46272
rect 25407 46208 25423 46272
rect 25487 46208 25503 46272
rect 25567 46208 25573 46272
rect 25257 46207 25573 46208
rect 29200 46188 29800 46278
rect 200 45508 800 45748
rect 7892 45728 8208 45729
rect 7892 45664 7898 45728
rect 7962 45664 7978 45728
rect 8042 45664 8058 45728
rect 8122 45664 8138 45728
rect 8202 45664 8208 45728
rect 7892 45663 8208 45664
rect 14838 45728 15154 45729
rect 14838 45664 14844 45728
rect 14908 45664 14924 45728
rect 14988 45664 15004 45728
rect 15068 45664 15084 45728
rect 15148 45664 15154 45728
rect 14838 45663 15154 45664
rect 21784 45728 22100 45729
rect 21784 45664 21790 45728
rect 21854 45664 21870 45728
rect 21934 45664 21950 45728
rect 22014 45664 22030 45728
rect 22094 45664 22100 45728
rect 21784 45663 22100 45664
rect 28730 45728 29046 45729
rect 28730 45664 28736 45728
rect 28800 45664 28816 45728
rect 28880 45664 28896 45728
rect 28960 45664 28976 45728
rect 29040 45664 29046 45728
rect 28730 45663 29046 45664
rect 29200 45508 29800 45748
rect 4419 45184 4735 45185
rect 4419 45120 4425 45184
rect 4489 45120 4505 45184
rect 4569 45120 4585 45184
rect 4649 45120 4665 45184
rect 4729 45120 4735 45184
rect 4419 45119 4735 45120
rect 11365 45184 11681 45185
rect 11365 45120 11371 45184
rect 11435 45120 11451 45184
rect 11515 45120 11531 45184
rect 11595 45120 11611 45184
rect 11675 45120 11681 45184
rect 11365 45119 11681 45120
rect 18311 45184 18627 45185
rect 18311 45120 18317 45184
rect 18381 45120 18397 45184
rect 18461 45120 18477 45184
rect 18541 45120 18557 45184
rect 18621 45120 18627 45184
rect 18311 45119 18627 45120
rect 25257 45184 25573 45185
rect 25257 45120 25263 45184
rect 25327 45120 25343 45184
rect 25407 45120 25423 45184
rect 25487 45120 25503 45184
rect 25567 45120 25573 45184
rect 25257 45119 25573 45120
rect 200 44978 800 45068
rect 2773 44978 2839 44981
rect 200 44976 2839 44978
rect 200 44920 2778 44976
rect 2834 44920 2839 44976
rect 200 44918 2839 44920
rect 200 44828 800 44918
rect 2773 44915 2839 44918
rect 28073 44978 28139 44981
rect 29200 44978 29800 45068
rect 28073 44976 29800 44978
rect 28073 44920 28078 44976
rect 28134 44920 29800 44976
rect 28073 44918 29800 44920
rect 28073 44915 28139 44918
rect 29200 44828 29800 44918
rect 7892 44640 8208 44641
rect 7892 44576 7898 44640
rect 7962 44576 7978 44640
rect 8042 44576 8058 44640
rect 8122 44576 8138 44640
rect 8202 44576 8208 44640
rect 7892 44575 8208 44576
rect 14838 44640 15154 44641
rect 14838 44576 14844 44640
rect 14908 44576 14924 44640
rect 14988 44576 15004 44640
rect 15068 44576 15084 44640
rect 15148 44576 15154 44640
rect 14838 44575 15154 44576
rect 21784 44640 22100 44641
rect 21784 44576 21790 44640
rect 21854 44576 21870 44640
rect 21934 44576 21950 44640
rect 22014 44576 22030 44640
rect 22094 44576 22100 44640
rect 21784 44575 22100 44576
rect 28730 44640 29046 44641
rect 28730 44576 28736 44640
rect 28800 44576 28816 44640
rect 28880 44576 28896 44640
rect 28960 44576 28976 44640
rect 29040 44576 29046 44640
rect 28730 44575 29046 44576
rect 200 44298 800 44388
rect 4153 44298 4219 44301
rect 200 44296 4219 44298
rect 200 44240 4158 44296
rect 4214 44240 4219 44296
rect 200 44238 4219 44240
rect 200 44148 800 44238
rect 4153 44235 4219 44238
rect 4419 44096 4735 44097
rect 4419 44032 4425 44096
rect 4489 44032 4505 44096
rect 4569 44032 4585 44096
rect 4649 44032 4665 44096
rect 4729 44032 4735 44096
rect 4419 44031 4735 44032
rect 11365 44096 11681 44097
rect 11365 44032 11371 44096
rect 11435 44032 11451 44096
rect 11515 44032 11531 44096
rect 11595 44032 11611 44096
rect 11675 44032 11681 44096
rect 11365 44031 11681 44032
rect 18311 44096 18627 44097
rect 18311 44032 18317 44096
rect 18381 44032 18397 44096
rect 18461 44032 18477 44096
rect 18541 44032 18557 44096
rect 18621 44032 18627 44096
rect 18311 44031 18627 44032
rect 25257 44096 25573 44097
rect 25257 44032 25263 44096
rect 25327 44032 25343 44096
rect 25407 44032 25423 44096
rect 25487 44032 25503 44096
rect 25567 44032 25573 44096
rect 25257 44031 25573 44032
rect 7892 43552 8208 43553
rect 7892 43488 7898 43552
rect 7962 43488 7978 43552
rect 8042 43488 8058 43552
rect 8122 43488 8138 43552
rect 8202 43488 8208 43552
rect 7892 43487 8208 43488
rect 14838 43552 15154 43553
rect 14838 43488 14844 43552
rect 14908 43488 14924 43552
rect 14988 43488 15004 43552
rect 15068 43488 15084 43552
rect 15148 43488 15154 43552
rect 14838 43487 15154 43488
rect 21784 43552 22100 43553
rect 21784 43488 21790 43552
rect 21854 43488 21870 43552
rect 21934 43488 21950 43552
rect 22014 43488 22030 43552
rect 22094 43488 22100 43552
rect 21784 43487 22100 43488
rect 28730 43552 29046 43553
rect 28730 43488 28736 43552
rect 28800 43488 28816 43552
rect 28880 43488 28896 43552
rect 28960 43488 28976 43552
rect 29040 43488 29046 43552
rect 28730 43487 29046 43488
rect 29200 43468 29800 43708
rect 200 42788 800 43028
rect 4419 43008 4735 43009
rect 4419 42944 4425 43008
rect 4489 42944 4505 43008
rect 4569 42944 4585 43008
rect 4649 42944 4665 43008
rect 4729 42944 4735 43008
rect 4419 42943 4735 42944
rect 11365 43008 11681 43009
rect 11365 42944 11371 43008
rect 11435 42944 11451 43008
rect 11515 42944 11531 43008
rect 11595 42944 11611 43008
rect 11675 42944 11681 43008
rect 11365 42943 11681 42944
rect 18311 43008 18627 43009
rect 18311 42944 18317 43008
rect 18381 42944 18397 43008
rect 18461 42944 18477 43008
rect 18541 42944 18557 43008
rect 18621 42944 18627 43008
rect 18311 42943 18627 42944
rect 25257 43008 25573 43009
rect 25257 42944 25263 43008
rect 25327 42944 25343 43008
rect 25407 42944 25423 43008
rect 25487 42944 25503 43008
rect 25567 42944 25573 43008
rect 25257 42943 25573 42944
rect 19425 42938 19491 42941
rect 19558 42938 19564 42940
rect 19425 42936 19564 42938
rect 19425 42880 19430 42936
rect 19486 42880 19564 42936
rect 19425 42878 19564 42880
rect 19425 42875 19491 42878
rect 19558 42876 19564 42878
rect 19628 42876 19634 42940
rect 28349 42938 28415 42941
rect 29200 42938 29800 43028
rect 28349 42936 29800 42938
rect 28349 42880 28354 42936
rect 28410 42880 29800 42936
rect 28349 42878 29800 42880
rect 28349 42875 28415 42878
rect 29200 42788 29800 42878
rect 7892 42464 8208 42465
rect 7892 42400 7898 42464
rect 7962 42400 7978 42464
rect 8042 42400 8058 42464
rect 8122 42400 8138 42464
rect 8202 42400 8208 42464
rect 7892 42399 8208 42400
rect 14838 42464 15154 42465
rect 14838 42400 14844 42464
rect 14908 42400 14924 42464
rect 14988 42400 15004 42464
rect 15068 42400 15084 42464
rect 15148 42400 15154 42464
rect 14838 42399 15154 42400
rect 21784 42464 22100 42465
rect 21784 42400 21790 42464
rect 21854 42400 21870 42464
rect 21934 42400 21950 42464
rect 22014 42400 22030 42464
rect 22094 42400 22100 42464
rect 21784 42399 22100 42400
rect 28730 42464 29046 42465
rect 28730 42400 28736 42464
rect 28800 42400 28816 42464
rect 28880 42400 28896 42464
rect 28960 42400 28976 42464
rect 29040 42400 29046 42464
rect 28730 42399 29046 42400
rect 200 42258 800 42348
rect 2773 42258 2839 42261
rect 200 42256 2839 42258
rect 200 42200 2778 42256
rect 2834 42200 2839 42256
rect 200 42198 2839 42200
rect 200 42108 800 42198
rect 2773 42195 2839 42198
rect 26049 42258 26115 42261
rect 29200 42258 29800 42348
rect 26049 42256 29800 42258
rect 26049 42200 26054 42256
rect 26110 42200 29800 42256
rect 26049 42198 29800 42200
rect 26049 42195 26115 42198
rect 29200 42108 29800 42198
rect 4419 41920 4735 41921
rect 4419 41856 4425 41920
rect 4489 41856 4505 41920
rect 4569 41856 4585 41920
rect 4649 41856 4665 41920
rect 4729 41856 4735 41920
rect 4419 41855 4735 41856
rect 11365 41920 11681 41921
rect 11365 41856 11371 41920
rect 11435 41856 11451 41920
rect 11515 41856 11531 41920
rect 11595 41856 11611 41920
rect 11675 41856 11681 41920
rect 11365 41855 11681 41856
rect 18311 41920 18627 41921
rect 18311 41856 18317 41920
rect 18381 41856 18397 41920
rect 18461 41856 18477 41920
rect 18541 41856 18557 41920
rect 18621 41856 18627 41920
rect 18311 41855 18627 41856
rect 25257 41920 25573 41921
rect 25257 41856 25263 41920
rect 25327 41856 25343 41920
rect 25407 41856 25423 41920
rect 25487 41856 25503 41920
rect 25567 41856 25573 41920
rect 25257 41855 25573 41856
rect 200 41578 800 41668
rect 1577 41578 1643 41581
rect 200 41576 1643 41578
rect 200 41520 1582 41576
rect 1638 41520 1643 41576
rect 200 41518 1643 41520
rect 200 41428 800 41518
rect 1577 41515 1643 41518
rect 27521 41578 27587 41581
rect 29200 41578 29800 41668
rect 27521 41576 29800 41578
rect 27521 41520 27526 41576
rect 27582 41520 29800 41576
rect 27521 41518 29800 41520
rect 27521 41515 27587 41518
rect 29200 41428 29800 41518
rect 7892 41376 8208 41377
rect 7892 41312 7898 41376
rect 7962 41312 7978 41376
rect 8042 41312 8058 41376
rect 8122 41312 8138 41376
rect 8202 41312 8208 41376
rect 7892 41311 8208 41312
rect 14838 41376 15154 41377
rect 14838 41312 14844 41376
rect 14908 41312 14924 41376
rect 14988 41312 15004 41376
rect 15068 41312 15084 41376
rect 15148 41312 15154 41376
rect 14838 41311 15154 41312
rect 21784 41376 22100 41377
rect 21784 41312 21790 41376
rect 21854 41312 21870 41376
rect 21934 41312 21950 41376
rect 22014 41312 22030 41376
rect 22094 41312 22100 41376
rect 21784 41311 22100 41312
rect 28730 41376 29046 41377
rect 28730 41312 28736 41376
rect 28800 41312 28816 41376
rect 28880 41312 28896 41376
rect 28960 41312 28976 41376
rect 29040 41312 29046 41376
rect 28730 41311 29046 41312
rect 200 40748 800 40988
rect 28625 40898 28691 40901
rect 29200 40898 29800 40988
rect 28625 40896 29800 40898
rect 28625 40840 28630 40896
rect 28686 40840 29800 40896
rect 28625 40838 29800 40840
rect 28625 40835 28691 40838
rect 4419 40832 4735 40833
rect 4419 40768 4425 40832
rect 4489 40768 4505 40832
rect 4569 40768 4585 40832
rect 4649 40768 4665 40832
rect 4729 40768 4735 40832
rect 4419 40767 4735 40768
rect 11365 40832 11681 40833
rect 11365 40768 11371 40832
rect 11435 40768 11451 40832
rect 11515 40768 11531 40832
rect 11595 40768 11611 40832
rect 11675 40768 11681 40832
rect 11365 40767 11681 40768
rect 18311 40832 18627 40833
rect 18311 40768 18317 40832
rect 18381 40768 18397 40832
rect 18461 40768 18477 40832
rect 18541 40768 18557 40832
rect 18621 40768 18627 40832
rect 18311 40767 18627 40768
rect 25257 40832 25573 40833
rect 25257 40768 25263 40832
rect 25327 40768 25343 40832
rect 25407 40768 25423 40832
rect 25487 40768 25503 40832
rect 25567 40768 25573 40832
rect 25257 40767 25573 40768
rect 29200 40748 29800 40838
rect 27521 40626 27587 40629
rect 27521 40624 29378 40626
rect 27521 40568 27526 40624
rect 27582 40568 29378 40624
rect 27521 40566 29378 40568
rect 27521 40563 27587 40566
rect 29318 40354 29378 40566
rect 29318 40308 29930 40354
rect 200 40068 800 40308
rect 29200 40294 29930 40308
rect 7892 40288 8208 40289
rect 7892 40224 7898 40288
rect 7962 40224 7978 40288
rect 8042 40224 8058 40288
rect 8122 40224 8138 40288
rect 8202 40224 8208 40288
rect 7892 40223 8208 40224
rect 14838 40288 15154 40289
rect 14838 40224 14844 40288
rect 14908 40224 14924 40288
rect 14988 40224 15004 40288
rect 15068 40224 15084 40288
rect 15148 40224 15154 40288
rect 14838 40223 15154 40224
rect 21784 40288 22100 40289
rect 21784 40224 21790 40288
rect 21854 40224 21870 40288
rect 21934 40224 21950 40288
rect 22014 40224 22030 40288
rect 22094 40224 22100 40288
rect 21784 40223 22100 40224
rect 28730 40288 29046 40289
rect 28730 40224 28736 40288
rect 28800 40224 28816 40288
rect 28880 40224 28896 40288
rect 28960 40224 28976 40288
rect 29040 40224 29046 40288
rect 28730 40223 29046 40224
rect 29200 40218 29800 40294
rect 29870 40218 29930 40294
rect 29200 40158 29930 40218
rect 29200 40068 29800 40158
rect 4419 39744 4735 39745
rect 4419 39680 4425 39744
rect 4489 39680 4505 39744
rect 4569 39680 4585 39744
rect 4649 39680 4665 39744
rect 4729 39680 4735 39744
rect 4419 39679 4735 39680
rect 11365 39744 11681 39745
rect 11365 39680 11371 39744
rect 11435 39680 11451 39744
rect 11515 39680 11531 39744
rect 11595 39680 11611 39744
rect 11675 39680 11681 39744
rect 11365 39679 11681 39680
rect 18311 39744 18627 39745
rect 18311 39680 18317 39744
rect 18381 39680 18397 39744
rect 18461 39680 18477 39744
rect 18541 39680 18557 39744
rect 18621 39680 18627 39744
rect 18311 39679 18627 39680
rect 25257 39744 25573 39745
rect 25257 39680 25263 39744
rect 25327 39680 25343 39744
rect 25407 39680 25423 39744
rect 25487 39680 25503 39744
rect 25567 39680 25573 39744
rect 25257 39679 25573 39680
rect 200 39388 800 39628
rect 26141 39538 26207 39541
rect 29200 39538 29800 39628
rect 26141 39536 29800 39538
rect 26141 39480 26146 39536
rect 26202 39480 29800 39536
rect 26141 39478 29800 39480
rect 26141 39475 26207 39478
rect 29200 39388 29800 39478
rect 7892 39200 8208 39201
rect 7892 39136 7898 39200
rect 7962 39136 7978 39200
rect 8042 39136 8058 39200
rect 8122 39136 8138 39200
rect 8202 39136 8208 39200
rect 7892 39135 8208 39136
rect 14838 39200 15154 39201
rect 14838 39136 14844 39200
rect 14908 39136 14924 39200
rect 14988 39136 15004 39200
rect 15068 39136 15084 39200
rect 15148 39136 15154 39200
rect 14838 39135 15154 39136
rect 21784 39200 22100 39201
rect 21784 39136 21790 39200
rect 21854 39136 21870 39200
rect 21934 39136 21950 39200
rect 22014 39136 22030 39200
rect 22094 39136 22100 39200
rect 21784 39135 22100 39136
rect 28730 39200 29046 39201
rect 28730 39136 28736 39200
rect 28800 39136 28816 39200
rect 28880 39136 28896 39200
rect 28960 39136 28976 39200
rect 29040 39136 29046 39200
rect 28730 39135 29046 39136
rect 200 38858 800 38948
rect 2773 38858 2839 38861
rect 200 38856 2839 38858
rect 200 38800 2778 38856
rect 2834 38800 2839 38856
rect 200 38798 2839 38800
rect 200 38708 800 38798
rect 2773 38795 2839 38798
rect 4419 38656 4735 38657
rect 4419 38592 4425 38656
rect 4489 38592 4505 38656
rect 4569 38592 4585 38656
rect 4649 38592 4665 38656
rect 4729 38592 4735 38656
rect 4419 38591 4735 38592
rect 11365 38656 11681 38657
rect 11365 38592 11371 38656
rect 11435 38592 11451 38656
rect 11515 38592 11531 38656
rect 11595 38592 11611 38656
rect 11675 38592 11681 38656
rect 11365 38591 11681 38592
rect 18311 38656 18627 38657
rect 18311 38592 18317 38656
rect 18381 38592 18397 38656
rect 18461 38592 18477 38656
rect 18541 38592 18557 38656
rect 18621 38592 18627 38656
rect 18311 38591 18627 38592
rect 25257 38656 25573 38657
rect 25257 38592 25263 38656
rect 25327 38592 25343 38656
rect 25407 38592 25423 38656
rect 25487 38592 25503 38656
rect 25567 38592 25573 38656
rect 25257 38591 25573 38592
rect 7892 38112 8208 38113
rect 7892 38048 7898 38112
rect 7962 38048 7978 38112
rect 8042 38048 8058 38112
rect 8122 38048 8138 38112
rect 8202 38048 8208 38112
rect 7892 38047 8208 38048
rect 14838 38112 15154 38113
rect 14838 38048 14844 38112
rect 14908 38048 14924 38112
rect 14988 38048 15004 38112
rect 15068 38048 15084 38112
rect 15148 38048 15154 38112
rect 14838 38047 15154 38048
rect 21784 38112 22100 38113
rect 21784 38048 21790 38112
rect 21854 38048 21870 38112
rect 21934 38048 21950 38112
rect 22014 38048 22030 38112
rect 22094 38048 22100 38112
rect 21784 38047 22100 38048
rect 28730 38112 29046 38113
rect 28730 38048 28736 38112
rect 28800 38048 28816 38112
rect 28880 38048 28896 38112
rect 28960 38048 28976 38112
rect 29040 38048 29046 38112
rect 28730 38047 29046 38048
rect 29200 38028 29800 38268
rect 200 37498 800 37588
rect 4419 37568 4735 37569
rect 4419 37504 4425 37568
rect 4489 37504 4505 37568
rect 4569 37504 4585 37568
rect 4649 37504 4665 37568
rect 4729 37504 4735 37568
rect 4419 37503 4735 37504
rect 11365 37568 11681 37569
rect 11365 37504 11371 37568
rect 11435 37504 11451 37568
rect 11515 37504 11531 37568
rect 11595 37504 11611 37568
rect 11675 37504 11681 37568
rect 11365 37503 11681 37504
rect 18311 37568 18627 37569
rect 18311 37504 18317 37568
rect 18381 37504 18397 37568
rect 18461 37504 18477 37568
rect 18541 37504 18557 37568
rect 18621 37504 18627 37568
rect 18311 37503 18627 37504
rect 25257 37568 25573 37569
rect 25257 37504 25263 37568
rect 25327 37504 25343 37568
rect 25407 37504 25423 37568
rect 25487 37504 25503 37568
rect 25567 37504 25573 37568
rect 25257 37503 25573 37504
rect 1577 37498 1643 37501
rect 200 37496 1643 37498
rect 200 37440 1582 37496
rect 1638 37440 1643 37496
rect 200 37438 1643 37440
rect 200 37348 800 37438
rect 1577 37435 1643 37438
rect 29200 37348 29800 37588
rect 7892 37024 8208 37025
rect 7892 36960 7898 37024
rect 7962 36960 7978 37024
rect 8042 36960 8058 37024
rect 8122 36960 8138 37024
rect 8202 36960 8208 37024
rect 7892 36959 8208 36960
rect 14838 37024 15154 37025
rect 14838 36960 14844 37024
rect 14908 36960 14924 37024
rect 14988 36960 15004 37024
rect 15068 36960 15084 37024
rect 15148 36960 15154 37024
rect 14838 36959 15154 36960
rect 21784 37024 22100 37025
rect 21784 36960 21790 37024
rect 21854 36960 21870 37024
rect 21934 36960 21950 37024
rect 22014 36960 22030 37024
rect 22094 36960 22100 37024
rect 21784 36959 22100 36960
rect 28730 37024 29046 37025
rect 28730 36960 28736 37024
rect 28800 36960 28816 37024
rect 28880 36960 28896 37024
rect 28960 36960 28976 37024
rect 29040 36960 29046 37024
rect 28730 36959 29046 36960
rect 200 36818 800 36908
rect 2865 36818 2931 36821
rect 200 36816 2931 36818
rect 200 36760 2870 36816
rect 2926 36760 2931 36816
rect 200 36758 2931 36760
rect 200 36668 800 36758
rect 2865 36755 2931 36758
rect 28349 36818 28415 36821
rect 29200 36818 29800 36908
rect 28349 36816 29800 36818
rect 28349 36760 28354 36816
rect 28410 36760 29800 36816
rect 28349 36758 29800 36760
rect 28349 36755 28415 36758
rect 29200 36668 29800 36758
rect 4419 36480 4735 36481
rect 4419 36416 4425 36480
rect 4489 36416 4505 36480
rect 4569 36416 4585 36480
rect 4649 36416 4665 36480
rect 4729 36416 4735 36480
rect 4419 36415 4735 36416
rect 11365 36480 11681 36481
rect 11365 36416 11371 36480
rect 11435 36416 11451 36480
rect 11515 36416 11531 36480
rect 11595 36416 11611 36480
rect 11675 36416 11681 36480
rect 11365 36415 11681 36416
rect 18311 36480 18627 36481
rect 18311 36416 18317 36480
rect 18381 36416 18397 36480
rect 18461 36416 18477 36480
rect 18541 36416 18557 36480
rect 18621 36416 18627 36480
rect 18311 36415 18627 36416
rect 25257 36480 25573 36481
rect 25257 36416 25263 36480
rect 25327 36416 25343 36480
rect 25407 36416 25423 36480
rect 25487 36416 25503 36480
rect 25567 36416 25573 36480
rect 25257 36415 25573 36416
rect 200 36138 800 36228
rect 2773 36138 2839 36141
rect 200 36136 2839 36138
rect 200 36080 2778 36136
rect 2834 36080 2839 36136
rect 200 36078 2839 36080
rect 200 35988 800 36078
rect 2773 36075 2839 36078
rect 28349 36138 28415 36141
rect 29200 36138 29800 36228
rect 28349 36136 29800 36138
rect 28349 36080 28354 36136
rect 28410 36080 29800 36136
rect 28349 36078 29800 36080
rect 28349 36075 28415 36078
rect 29200 35988 29800 36078
rect 7892 35936 8208 35937
rect 7892 35872 7898 35936
rect 7962 35872 7978 35936
rect 8042 35872 8058 35936
rect 8122 35872 8138 35936
rect 8202 35872 8208 35936
rect 7892 35871 8208 35872
rect 14838 35936 15154 35937
rect 14838 35872 14844 35936
rect 14908 35872 14924 35936
rect 14988 35872 15004 35936
rect 15068 35872 15084 35936
rect 15148 35872 15154 35936
rect 14838 35871 15154 35872
rect 21784 35936 22100 35937
rect 21784 35872 21790 35936
rect 21854 35872 21870 35936
rect 21934 35872 21950 35936
rect 22014 35872 22030 35936
rect 22094 35872 22100 35936
rect 21784 35871 22100 35872
rect 28730 35936 29046 35937
rect 28730 35872 28736 35936
rect 28800 35872 28816 35936
rect 28880 35872 28896 35936
rect 28960 35872 28976 35936
rect 29040 35872 29046 35936
rect 28730 35871 29046 35872
rect 200 35308 800 35548
rect 4419 35392 4735 35393
rect 4419 35328 4425 35392
rect 4489 35328 4505 35392
rect 4569 35328 4585 35392
rect 4649 35328 4665 35392
rect 4729 35328 4735 35392
rect 4419 35327 4735 35328
rect 11365 35392 11681 35393
rect 11365 35328 11371 35392
rect 11435 35328 11451 35392
rect 11515 35328 11531 35392
rect 11595 35328 11611 35392
rect 11675 35328 11681 35392
rect 11365 35327 11681 35328
rect 18311 35392 18627 35393
rect 18311 35328 18317 35392
rect 18381 35328 18397 35392
rect 18461 35328 18477 35392
rect 18541 35328 18557 35392
rect 18621 35328 18627 35392
rect 18311 35327 18627 35328
rect 25257 35392 25573 35393
rect 25257 35328 25263 35392
rect 25327 35328 25343 35392
rect 25407 35328 25423 35392
rect 25487 35328 25503 35392
rect 25567 35328 25573 35392
rect 25257 35327 25573 35328
rect 29200 35308 29800 35548
rect 200 34778 800 34868
rect 7892 34848 8208 34849
rect 7892 34784 7898 34848
rect 7962 34784 7978 34848
rect 8042 34784 8058 34848
rect 8122 34784 8138 34848
rect 8202 34784 8208 34848
rect 7892 34783 8208 34784
rect 14838 34848 15154 34849
rect 14838 34784 14844 34848
rect 14908 34784 14924 34848
rect 14988 34784 15004 34848
rect 15068 34784 15084 34848
rect 15148 34784 15154 34848
rect 14838 34783 15154 34784
rect 21784 34848 22100 34849
rect 21784 34784 21790 34848
rect 21854 34784 21870 34848
rect 21934 34784 21950 34848
rect 22014 34784 22030 34848
rect 22094 34784 22100 34848
rect 21784 34783 22100 34784
rect 28730 34848 29046 34849
rect 28730 34784 28736 34848
rect 28800 34784 28816 34848
rect 28880 34784 28896 34848
rect 28960 34784 28976 34848
rect 29040 34784 29046 34848
rect 28730 34783 29046 34784
rect 2773 34778 2839 34781
rect 200 34776 2839 34778
rect 200 34720 2778 34776
rect 2834 34720 2839 34776
rect 200 34718 2839 34720
rect 200 34628 800 34718
rect 2773 34715 2839 34718
rect 29200 34628 29800 34868
rect 4419 34304 4735 34305
rect 4419 34240 4425 34304
rect 4489 34240 4505 34304
rect 4569 34240 4585 34304
rect 4649 34240 4665 34304
rect 4729 34240 4735 34304
rect 4419 34239 4735 34240
rect 11365 34304 11681 34305
rect 11365 34240 11371 34304
rect 11435 34240 11451 34304
rect 11515 34240 11531 34304
rect 11595 34240 11611 34304
rect 11675 34240 11681 34304
rect 11365 34239 11681 34240
rect 18311 34304 18627 34305
rect 18311 34240 18317 34304
rect 18381 34240 18397 34304
rect 18461 34240 18477 34304
rect 18541 34240 18557 34304
rect 18621 34240 18627 34304
rect 18311 34239 18627 34240
rect 25257 34304 25573 34305
rect 25257 34240 25263 34304
rect 25327 34240 25343 34304
rect 25407 34240 25423 34304
rect 25487 34240 25503 34304
rect 25567 34240 25573 34304
rect 25257 34239 25573 34240
rect 200 33948 800 34188
rect 27521 34098 27587 34101
rect 29200 34098 29800 34188
rect 27521 34096 29800 34098
rect 27521 34040 27526 34096
rect 27582 34040 29800 34096
rect 27521 34038 29800 34040
rect 27521 34035 27587 34038
rect 29200 33948 29800 34038
rect 7892 33760 8208 33761
rect 7892 33696 7898 33760
rect 7962 33696 7978 33760
rect 8042 33696 8058 33760
rect 8122 33696 8138 33760
rect 8202 33696 8208 33760
rect 7892 33695 8208 33696
rect 14838 33760 15154 33761
rect 14838 33696 14844 33760
rect 14908 33696 14924 33760
rect 14988 33696 15004 33760
rect 15068 33696 15084 33760
rect 15148 33696 15154 33760
rect 14838 33695 15154 33696
rect 21784 33760 22100 33761
rect 21784 33696 21790 33760
rect 21854 33696 21870 33760
rect 21934 33696 21950 33760
rect 22014 33696 22030 33760
rect 22094 33696 22100 33760
rect 21784 33695 22100 33696
rect 28730 33760 29046 33761
rect 28730 33696 28736 33760
rect 28800 33696 28816 33760
rect 28880 33696 28896 33760
rect 28960 33696 28976 33760
rect 29040 33696 29046 33760
rect 28730 33695 29046 33696
rect 200 33418 800 33508
rect 3509 33418 3575 33421
rect 200 33416 3575 33418
rect 200 33360 3514 33416
rect 3570 33360 3575 33416
rect 200 33358 3575 33360
rect 200 33268 800 33358
rect 3509 33355 3575 33358
rect 4419 33216 4735 33217
rect 4419 33152 4425 33216
rect 4489 33152 4505 33216
rect 4569 33152 4585 33216
rect 4649 33152 4665 33216
rect 4729 33152 4735 33216
rect 4419 33151 4735 33152
rect 11365 33216 11681 33217
rect 11365 33152 11371 33216
rect 11435 33152 11451 33216
rect 11515 33152 11531 33216
rect 11595 33152 11611 33216
rect 11675 33152 11681 33216
rect 11365 33151 11681 33152
rect 18311 33216 18627 33217
rect 18311 33152 18317 33216
rect 18381 33152 18397 33216
rect 18461 33152 18477 33216
rect 18541 33152 18557 33216
rect 18621 33152 18627 33216
rect 18311 33151 18627 33152
rect 25257 33216 25573 33217
rect 25257 33152 25263 33216
rect 25327 33152 25343 33216
rect 25407 33152 25423 33216
rect 25487 33152 25503 33216
rect 25567 33152 25573 33216
rect 25257 33151 25573 33152
rect 27521 33010 27587 33013
rect 27521 33008 29378 33010
rect 27521 32952 27526 33008
rect 27582 32952 29378 33008
rect 27521 32950 29378 32952
rect 27521 32947 27587 32950
rect 29318 32874 29378 32950
rect 29318 32828 29930 32874
rect 29200 32814 29930 32828
rect 29200 32738 29800 32814
rect 29870 32738 29930 32814
rect 29200 32678 29930 32738
rect 7892 32672 8208 32673
rect 7892 32608 7898 32672
rect 7962 32608 7978 32672
rect 8042 32608 8058 32672
rect 8122 32608 8138 32672
rect 8202 32608 8208 32672
rect 7892 32607 8208 32608
rect 14838 32672 15154 32673
rect 14838 32608 14844 32672
rect 14908 32608 14924 32672
rect 14988 32608 15004 32672
rect 15068 32608 15084 32672
rect 15148 32608 15154 32672
rect 14838 32607 15154 32608
rect 21784 32672 22100 32673
rect 21784 32608 21790 32672
rect 21854 32608 21870 32672
rect 21934 32608 21950 32672
rect 22014 32608 22030 32672
rect 22094 32608 22100 32672
rect 21784 32607 22100 32608
rect 28730 32672 29046 32673
rect 28730 32608 28736 32672
rect 28800 32608 28816 32672
rect 28880 32608 28896 32672
rect 28960 32608 28976 32672
rect 29040 32608 29046 32672
rect 28730 32607 29046 32608
rect 29200 32588 29800 32678
rect 200 32058 800 32148
rect 4419 32128 4735 32129
rect 4419 32064 4425 32128
rect 4489 32064 4505 32128
rect 4569 32064 4585 32128
rect 4649 32064 4665 32128
rect 4729 32064 4735 32128
rect 4419 32063 4735 32064
rect 11365 32128 11681 32129
rect 11365 32064 11371 32128
rect 11435 32064 11451 32128
rect 11515 32064 11531 32128
rect 11595 32064 11611 32128
rect 11675 32064 11681 32128
rect 11365 32063 11681 32064
rect 18311 32128 18627 32129
rect 18311 32064 18317 32128
rect 18381 32064 18397 32128
rect 18461 32064 18477 32128
rect 18541 32064 18557 32128
rect 18621 32064 18627 32128
rect 18311 32063 18627 32064
rect 25257 32128 25573 32129
rect 25257 32064 25263 32128
rect 25327 32064 25343 32128
rect 25407 32064 25423 32128
rect 25487 32064 25503 32128
rect 25567 32064 25573 32128
rect 25257 32063 25573 32064
rect 2957 32058 3023 32061
rect 200 32056 3023 32058
rect 200 32000 2962 32056
rect 3018 32000 3023 32056
rect 200 31998 3023 32000
rect 200 31908 800 31998
rect 2957 31995 3023 31998
rect 28257 32058 28323 32061
rect 29200 32058 29800 32148
rect 28257 32056 29800 32058
rect 28257 32000 28262 32056
rect 28318 32000 29800 32056
rect 28257 31998 29800 32000
rect 28257 31995 28323 31998
rect 29200 31908 29800 31998
rect 7892 31584 8208 31585
rect 7892 31520 7898 31584
rect 7962 31520 7978 31584
rect 8042 31520 8058 31584
rect 8122 31520 8138 31584
rect 8202 31520 8208 31584
rect 7892 31519 8208 31520
rect 14838 31584 15154 31585
rect 14838 31520 14844 31584
rect 14908 31520 14924 31584
rect 14988 31520 15004 31584
rect 15068 31520 15084 31584
rect 15148 31520 15154 31584
rect 14838 31519 15154 31520
rect 21784 31584 22100 31585
rect 21784 31520 21790 31584
rect 21854 31520 21870 31584
rect 21934 31520 21950 31584
rect 22014 31520 22030 31584
rect 22094 31520 22100 31584
rect 21784 31519 22100 31520
rect 28730 31584 29046 31585
rect 28730 31520 28736 31584
rect 28800 31520 28816 31584
rect 28880 31520 28896 31584
rect 28960 31520 28976 31584
rect 29040 31520 29046 31584
rect 28730 31519 29046 31520
rect 200 31228 800 31468
rect 27521 31378 27587 31381
rect 29200 31378 29800 31468
rect 27521 31376 29800 31378
rect 27521 31320 27526 31376
rect 27582 31320 29800 31376
rect 27521 31318 29800 31320
rect 27521 31315 27587 31318
rect 29200 31228 29800 31318
rect 4419 31040 4735 31041
rect 4419 30976 4425 31040
rect 4489 30976 4505 31040
rect 4569 30976 4585 31040
rect 4649 30976 4665 31040
rect 4729 30976 4735 31040
rect 4419 30975 4735 30976
rect 11365 31040 11681 31041
rect 11365 30976 11371 31040
rect 11435 30976 11451 31040
rect 11515 30976 11531 31040
rect 11595 30976 11611 31040
rect 11675 30976 11681 31040
rect 11365 30975 11681 30976
rect 18311 31040 18627 31041
rect 18311 30976 18317 31040
rect 18381 30976 18397 31040
rect 18461 30976 18477 31040
rect 18541 30976 18557 31040
rect 18621 30976 18627 31040
rect 18311 30975 18627 30976
rect 25257 31040 25573 31041
rect 25257 30976 25263 31040
rect 25327 30976 25343 31040
rect 25407 30976 25423 31040
rect 25487 30976 25503 31040
rect 25567 30976 25573 31040
rect 25257 30975 25573 30976
rect 200 30548 800 30788
rect 26141 30698 26207 30701
rect 29200 30698 29800 30788
rect 26141 30696 29800 30698
rect 26141 30640 26146 30696
rect 26202 30640 29800 30696
rect 26141 30638 29800 30640
rect 26141 30635 26207 30638
rect 29200 30548 29800 30638
rect 7892 30496 8208 30497
rect 7892 30432 7898 30496
rect 7962 30432 7978 30496
rect 8042 30432 8058 30496
rect 8122 30432 8138 30496
rect 8202 30432 8208 30496
rect 7892 30431 8208 30432
rect 14838 30496 15154 30497
rect 14838 30432 14844 30496
rect 14908 30432 14924 30496
rect 14988 30432 15004 30496
rect 15068 30432 15084 30496
rect 15148 30432 15154 30496
rect 14838 30431 15154 30432
rect 21784 30496 22100 30497
rect 21784 30432 21790 30496
rect 21854 30432 21870 30496
rect 21934 30432 21950 30496
rect 22014 30432 22030 30496
rect 22094 30432 22100 30496
rect 21784 30431 22100 30432
rect 28730 30496 29046 30497
rect 28730 30432 28736 30496
rect 28800 30432 28816 30496
rect 28880 30432 28896 30496
rect 28960 30432 28976 30496
rect 29040 30432 29046 30496
rect 28730 30431 29046 30432
rect 200 30018 800 30108
rect 1577 30018 1643 30021
rect 200 30016 1643 30018
rect 200 29960 1582 30016
rect 1638 29960 1643 30016
rect 200 29958 1643 29960
rect 200 29868 800 29958
rect 1577 29955 1643 29958
rect 28349 30018 28415 30021
rect 29200 30018 29800 30108
rect 28349 30016 29800 30018
rect 28349 29960 28354 30016
rect 28410 29960 29800 30016
rect 28349 29958 29800 29960
rect 28349 29955 28415 29958
rect 4419 29952 4735 29953
rect 4419 29888 4425 29952
rect 4489 29888 4505 29952
rect 4569 29888 4585 29952
rect 4649 29888 4665 29952
rect 4729 29888 4735 29952
rect 4419 29887 4735 29888
rect 11365 29952 11681 29953
rect 11365 29888 11371 29952
rect 11435 29888 11451 29952
rect 11515 29888 11531 29952
rect 11595 29888 11611 29952
rect 11675 29888 11681 29952
rect 11365 29887 11681 29888
rect 18311 29952 18627 29953
rect 18311 29888 18317 29952
rect 18381 29888 18397 29952
rect 18461 29888 18477 29952
rect 18541 29888 18557 29952
rect 18621 29888 18627 29952
rect 18311 29887 18627 29888
rect 25257 29952 25573 29953
rect 25257 29888 25263 29952
rect 25327 29888 25343 29952
rect 25407 29888 25423 29952
rect 25487 29888 25503 29952
rect 25567 29888 25573 29952
rect 25257 29887 25573 29888
rect 29200 29868 29800 29958
rect 200 29188 800 29428
rect 7892 29408 8208 29409
rect 7892 29344 7898 29408
rect 7962 29344 7978 29408
rect 8042 29344 8058 29408
rect 8122 29344 8138 29408
rect 8202 29344 8208 29408
rect 7892 29343 8208 29344
rect 14838 29408 15154 29409
rect 14838 29344 14844 29408
rect 14908 29344 14924 29408
rect 14988 29344 15004 29408
rect 15068 29344 15084 29408
rect 15148 29344 15154 29408
rect 14838 29343 15154 29344
rect 21784 29408 22100 29409
rect 21784 29344 21790 29408
rect 21854 29344 21870 29408
rect 21934 29344 21950 29408
rect 22014 29344 22030 29408
rect 22094 29344 22100 29408
rect 21784 29343 22100 29344
rect 28730 29408 29046 29409
rect 28730 29344 28736 29408
rect 28800 29344 28816 29408
rect 28880 29344 28896 29408
rect 28960 29344 28976 29408
rect 29040 29344 29046 29408
rect 28730 29343 29046 29344
rect 29200 29338 29800 29428
rect 29200 29278 29930 29338
rect 29200 29202 29800 29278
rect 29870 29202 29930 29278
rect 29200 29188 29930 29202
rect 29318 29142 29930 29188
rect 24853 29066 24919 29069
rect 29318 29066 29378 29142
rect 24853 29064 29378 29066
rect 24853 29008 24858 29064
rect 24914 29008 29378 29064
rect 24853 29006 29378 29008
rect 24853 29003 24919 29006
rect 4419 28864 4735 28865
rect 4419 28800 4425 28864
rect 4489 28800 4505 28864
rect 4569 28800 4585 28864
rect 4649 28800 4665 28864
rect 4729 28800 4735 28864
rect 4419 28799 4735 28800
rect 11365 28864 11681 28865
rect 11365 28800 11371 28864
rect 11435 28800 11451 28864
rect 11515 28800 11531 28864
rect 11595 28800 11611 28864
rect 11675 28800 11681 28864
rect 11365 28799 11681 28800
rect 18311 28864 18627 28865
rect 18311 28800 18317 28864
rect 18381 28800 18397 28864
rect 18461 28800 18477 28864
rect 18541 28800 18557 28864
rect 18621 28800 18627 28864
rect 18311 28799 18627 28800
rect 25257 28864 25573 28865
rect 25257 28800 25263 28864
rect 25327 28800 25343 28864
rect 25407 28800 25423 28864
rect 25487 28800 25503 28864
rect 25567 28800 25573 28864
rect 25257 28799 25573 28800
rect 200 28508 800 28748
rect 27521 28658 27587 28661
rect 29200 28658 29800 28748
rect 27521 28656 29800 28658
rect 27521 28600 27526 28656
rect 27582 28600 29800 28656
rect 27521 28598 29800 28600
rect 27521 28595 27587 28598
rect 29200 28508 29800 28598
rect 7892 28320 8208 28321
rect 7892 28256 7898 28320
rect 7962 28256 7978 28320
rect 8042 28256 8058 28320
rect 8122 28256 8138 28320
rect 8202 28256 8208 28320
rect 7892 28255 8208 28256
rect 14838 28320 15154 28321
rect 14838 28256 14844 28320
rect 14908 28256 14924 28320
rect 14988 28256 15004 28320
rect 15068 28256 15084 28320
rect 15148 28256 15154 28320
rect 14838 28255 15154 28256
rect 21784 28320 22100 28321
rect 21784 28256 21790 28320
rect 21854 28256 21870 28320
rect 21934 28256 21950 28320
rect 22014 28256 22030 28320
rect 22094 28256 22100 28320
rect 21784 28255 22100 28256
rect 28730 28320 29046 28321
rect 28730 28256 28736 28320
rect 28800 28256 28816 28320
rect 28880 28256 28896 28320
rect 28960 28256 28976 28320
rect 29040 28256 29046 28320
rect 28730 28255 29046 28256
rect 200 27978 800 28068
rect 1577 27978 1643 27981
rect 200 27976 1643 27978
rect 200 27920 1582 27976
rect 1638 27920 1643 27976
rect 200 27918 1643 27920
rect 200 27828 800 27918
rect 1577 27915 1643 27918
rect 4419 27776 4735 27777
rect 4419 27712 4425 27776
rect 4489 27712 4505 27776
rect 4569 27712 4585 27776
rect 4649 27712 4665 27776
rect 4729 27712 4735 27776
rect 4419 27711 4735 27712
rect 11365 27776 11681 27777
rect 11365 27712 11371 27776
rect 11435 27712 11451 27776
rect 11515 27712 11531 27776
rect 11595 27712 11611 27776
rect 11675 27712 11681 27776
rect 11365 27711 11681 27712
rect 18311 27776 18627 27777
rect 18311 27712 18317 27776
rect 18381 27712 18397 27776
rect 18461 27712 18477 27776
rect 18541 27712 18557 27776
rect 18621 27712 18627 27776
rect 18311 27711 18627 27712
rect 25257 27776 25573 27777
rect 25257 27712 25263 27776
rect 25327 27712 25343 27776
rect 25407 27712 25423 27776
rect 25487 27712 25503 27776
rect 25567 27712 25573 27776
rect 25257 27711 25573 27712
rect 27521 27570 27587 27573
rect 27521 27568 29378 27570
rect 27521 27512 27526 27568
rect 27582 27512 29378 27568
rect 27521 27510 29378 27512
rect 27521 27507 27587 27510
rect 29318 27434 29378 27510
rect 29318 27388 29930 27434
rect 29200 27374 29930 27388
rect 29200 27298 29800 27374
rect 29870 27298 29930 27374
rect 29200 27238 29930 27298
rect 7892 27232 8208 27233
rect 7892 27168 7898 27232
rect 7962 27168 7978 27232
rect 8042 27168 8058 27232
rect 8122 27168 8138 27232
rect 8202 27168 8208 27232
rect 7892 27167 8208 27168
rect 14838 27232 15154 27233
rect 14838 27168 14844 27232
rect 14908 27168 14924 27232
rect 14988 27168 15004 27232
rect 15068 27168 15084 27232
rect 15148 27168 15154 27232
rect 14838 27167 15154 27168
rect 21784 27232 22100 27233
rect 21784 27168 21790 27232
rect 21854 27168 21870 27232
rect 21934 27168 21950 27232
rect 22014 27168 22030 27232
rect 22094 27168 22100 27232
rect 21784 27167 22100 27168
rect 28730 27232 29046 27233
rect 28730 27168 28736 27232
rect 28800 27168 28816 27232
rect 28880 27168 28896 27232
rect 28960 27168 28976 27232
rect 29040 27168 29046 27232
rect 28730 27167 29046 27168
rect 29200 27148 29800 27238
rect 200 26468 800 26708
rect 4419 26688 4735 26689
rect 4419 26624 4425 26688
rect 4489 26624 4505 26688
rect 4569 26624 4585 26688
rect 4649 26624 4665 26688
rect 4729 26624 4735 26688
rect 4419 26623 4735 26624
rect 11365 26688 11681 26689
rect 11365 26624 11371 26688
rect 11435 26624 11451 26688
rect 11515 26624 11531 26688
rect 11595 26624 11611 26688
rect 11675 26624 11681 26688
rect 11365 26623 11681 26624
rect 18311 26688 18627 26689
rect 18311 26624 18317 26688
rect 18381 26624 18397 26688
rect 18461 26624 18477 26688
rect 18541 26624 18557 26688
rect 18621 26624 18627 26688
rect 18311 26623 18627 26624
rect 25257 26688 25573 26689
rect 25257 26624 25263 26688
rect 25327 26624 25343 26688
rect 25407 26624 25423 26688
rect 25487 26624 25503 26688
rect 25567 26624 25573 26688
rect 25257 26623 25573 26624
rect 27429 26618 27495 26621
rect 29200 26618 29800 26708
rect 27429 26616 29800 26618
rect 27429 26560 27434 26616
rect 27490 26560 29800 26616
rect 27429 26558 29800 26560
rect 27429 26555 27495 26558
rect 29200 26468 29800 26558
rect 7892 26144 8208 26145
rect 7892 26080 7898 26144
rect 7962 26080 7978 26144
rect 8042 26080 8058 26144
rect 8122 26080 8138 26144
rect 8202 26080 8208 26144
rect 7892 26079 8208 26080
rect 14838 26144 15154 26145
rect 14838 26080 14844 26144
rect 14908 26080 14924 26144
rect 14988 26080 15004 26144
rect 15068 26080 15084 26144
rect 15148 26080 15154 26144
rect 14838 26079 15154 26080
rect 21784 26144 22100 26145
rect 21784 26080 21790 26144
rect 21854 26080 21870 26144
rect 21934 26080 21950 26144
rect 22014 26080 22030 26144
rect 22094 26080 22100 26144
rect 21784 26079 22100 26080
rect 28730 26144 29046 26145
rect 28730 26080 28736 26144
rect 28800 26080 28816 26144
rect 28880 26080 28896 26144
rect 28960 26080 28976 26144
rect 29040 26080 29046 26144
rect 28730 26079 29046 26080
rect 200 25938 800 26028
rect 2773 25938 2839 25941
rect 200 25936 2839 25938
rect 200 25880 2778 25936
rect 2834 25880 2839 25936
rect 200 25878 2839 25880
rect 200 25788 800 25878
rect 2773 25875 2839 25878
rect 29200 25788 29800 26028
rect 4419 25600 4735 25601
rect 4419 25536 4425 25600
rect 4489 25536 4505 25600
rect 4569 25536 4585 25600
rect 4649 25536 4665 25600
rect 4729 25536 4735 25600
rect 4419 25535 4735 25536
rect 11365 25600 11681 25601
rect 11365 25536 11371 25600
rect 11435 25536 11451 25600
rect 11515 25536 11531 25600
rect 11595 25536 11611 25600
rect 11675 25536 11681 25600
rect 11365 25535 11681 25536
rect 18311 25600 18627 25601
rect 18311 25536 18317 25600
rect 18381 25536 18397 25600
rect 18461 25536 18477 25600
rect 18541 25536 18557 25600
rect 18621 25536 18627 25600
rect 18311 25535 18627 25536
rect 25257 25600 25573 25601
rect 25257 25536 25263 25600
rect 25327 25536 25343 25600
rect 25407 25536 25423 25600
rect 25487 25536 25503 25600
rect 25567 25536 25573 25600
rect 25257 25535 25573 25536
rect 200 25258 800 25348
rect 1577 25258 1643 25261
rect 200 25256 1643 25258
rect 200 25200 1582 25256
rect 1638 25200 1643 25256
rect 200 25198 1643 25200
rect 200 25108 800 25198
rect 1577 25195 1643 25198
rect 28349 25258 28415 25261
rect 29200 25258 29800 25348
rect 28349 25256 29800 25258
rect 28349 25200 28354 25256
rect 28410 25200 29800 25256
rect 28349 25198 29800 25200
rect 28349 25195 28415 25198
rect 29200 25108 29800 25198
rect 7892 25056 8208 25057
rect 7892 24992 7898 25056
rect 7962 24992 7978 25056
rect 8042 24992 8058 25056
rect 8122 24992 8138 25056
rect 8202 24992 8208 25056
rect 7892 24991 8208 24992
rect 14838 25056 15154 25057
rect 14838 24992 14844 25056
rect 14908 24992 14924 25056
rect 14988 24992 15004 25056
rect 15068 24992 15084 25056
rect 15148 24992 15154 25056
rect 14838 24991 15154 24992
rect 21784 25056 22100 25057
rect 21784 24992 21790 25056
rect 21854 24992 21870 25056
rect 21934 24992 21950 25056
rect 22014 24992 22030 25056
rect 22094 24992 22100 25056
rect 21784 24991 22100 24992
rect 28730 25056 29046 25057
rect 28730 24992 28736 25056
rect 28800 24992 28816 25056
rect 28880 24992 28896 25056
rect 28960 24992 28976 25056
rect 29040 24992 29046 25056
rect 28730 24991 29046 24992
rect 18781 24714 18847 24717
rect 19558 24714 19564 24716
rect 18781 24712 19564 24714
rect 200 24428 800 24668
rect 18781 24656 18786 24712
rect 18842 24656 19564 24712
rect 18781 24654 19564 24656
rect 18781 24651 18847 24654
rect 19558 24652 19564 24654
rect 19628 24652 19634 24716
rect 28349 24578 28415 24581
rect 29200 24578 29800 24668
rect 28349 24576 29800 24578
rect 28349 24520 28354 24576
rect 28410 24520 29800 24576
rect 28349 24518 29800 24520
rect 28349 24515 28415 24518
rect 4419 24512 4735 24513
rect 4419 24448 4425 24512
rect 4489 24448 4505 24512
rect 4569 24448 4585 24512
rect 4649 24448 4665 24512
rect 4729 24448 4735 24512
rect 4419 24447 4735 24448
rect 11365 24512 11681 24513
rect 11365 24448 11371 24512
rect 11435 24448 11451 24512
rect 11515 24448 11531 24512
rect 11595 24448 11611 24512
rect 11675 24448 11681 24512
rect 11365 24447 11681 24448
rect 18311 24512 18627 24513
rect 18311 24448 18317 24512
rect 18381 24448 18397 24512
rect 18461 24448 18477 24512
rect 18541 24448 18557 24512
rect 18621 24448 18627 24512
rect 18311 24447 18627 24448
rect 25257 24512 25573 24513
rect 25257 24448 25263 24512
rect 25327 24448 25343 24512
rect 25407 24448 25423 24512
rect 25487 24448 25503 24512
rect 25567 24448 25573 24512
rect 25257 24447 25573 24448
rect 29200 24428 29800 24518
rect 200 23748 800 23988
rect 7892 23968 8208 23969
rect 7892 23904 7898 23968
rect 7962 23904 7978 23968
rect 8042 23904 8058 23968
rect 8122 23904 8138 23968
rect 8202 23904 8208 23968
rect 7892 23903 8208 23904
rect 14838 23968 15154 23969
rect 14838 23904 14844 23968
rect 14908 23904 14924 23968
rect 14988 23904 15004 23968
rect 15068 23904 15084 23968
rect 15148 23904 15154 23968
rect 14838 23903 15154 23904
rect 21784 23968 22100 23969
rect 21784 23904 21790 23968
rect 21854 23904 21870 23968
rect 21934 23904 21950 23968
rect 22014 23904 22030 23968
rect 22094 23904 22100 23968
rect 21784 23903 22100 23904
rect 28730 23968 29046 23969
rect 28730 23904 28736 23968
rect 28800 23904 28816 23968
rect 28880 23904 28896 23968
rect 28960 23904 28976 23968
rect 29040 23904 29046 23968
rect 28730 23903 29046 23904
rect 29200 23898 29800 23988
rect 29913 23898 29979 23901
rect 29200 23896 29979 23898
rect 29200 23840 29918 23896
rect 29974 23840 29979 23896
rect 29200 23838 29979 23840
rect 29200 23748 29800 23838
rect 29913 23835 29979 23838
rect 4419 23424 4735 23425
rect 4419 23360 4425 23424
rect 4489 23360 4505 23424
rect 4569 23360 4585 23424
rect 4649 23360 4665 23424
rect 4729 23360 4735 23424
rect 4419 23359 4735 23360
rect 11365 23424 11681 23425
rect 11365 23360 11371 23424
rect 11435 23360 11451 23424
rect 11515 23360 11531 23424
rect 11595 23360 11611 23424
rect 11675 23360 11681 23424
rect 11365 23359 11681 23360
rect 18311 23424 18627 23425
rect 18311 23360 18317 23424
rect 18381 23360 18397 23424
rect 18461 23360 18477 23424
rect 18541 23360 18557 23424
rect 18621 23360 18627 23424
rect 18311 23359 18627 23360
rect 25257 23424 25573 23425
rect 25257 23360 25263 23424
rect 25327 23360 25343 23424
rect 25407 23360 25423 23424
rect 25487 23360 25503 23424
rect 25567 23360 25573 23424
rect 25257 23359 25573 23360
rect 200 23068 800 23308
rect 29200 23068 29800 23308
rect 7892 22880 8208 22881
rect 7892 22816 7898 22880
rect 7962 22816 7978 22880
rect 8042 22816 8058 22880
rect 8122 22816 8138 22880
rect 8202 22816 8208 22880
rect 7892 22815 8208 22816
rect 14838 22880 15154 22881
rect 14838 22816 14844 22880
rect 14908 22816 14924 22880
rect 14988 22816 15004 22880
rect 15068 22816 15084 22880
rect 15148 22816 15154 22880
rect 14838 22815 15154 22816
rect 21784 22880 22100 22881
rect 21784 22816 21790 22880
rect 21854 22816 21870 22880
rect 21934 22816 21950 22880
rect 22014 22816 22030 22880
rect 22094 22816 22100 22880
rect 21784 22815 22100 22816
rect 28730 22880 29046 22881
rect 28730 22816 28736 22880
rect 28800 22816 28816 22880
rect 28880 22816 28896 22880
rect 28960 22816 28976 22880
rect 29040 22816 29046 22880
rect 28730 22815 29046 22816
rect 200 22388 800 22628
rect 4419 22336 4735 22337
rect 4419 22272 4425 22336
rect 4489 22272 4505 22336
rect 4569 22272 4585 22336
rect 4649 22272 4665 22336
rect 4729 22272 4735 22336
rect 4419 22271 4735 22272
rect 11365 22336 11681 22337
rect 11365 22272 11371 22336
rect 11435 22272 11451 22336
rect 11515 22272 11531 22336
rect 11595 22272 11611 22336
rect 11675 22272 11681 22336
rect 11365 22271 11681 22272
rect 18311 22336 18627 22337
rect 18311 22272 18317 22336
rect 18381 22272 18397 22336
rect 18461 22272 18477 22336
rect 18541 22272 18557 22336
rect 18621 22272 18627 22336
rect 18311 22271 18627 22272
rect 25257 22336 25573 22337
rect 25257 22272 25263 22336
rect 25327 22272 25343 22336
rect 25407 22272 25423 22336
rect 25487 22272 25503 22336
rect 25567 22272 25573 22336
rect 25257 22271 25573 22272
rect 27521 21994 27587 21997
rect 27521 21992 29930 21994
rect 27521 21936 27526 21992
rect 27582 21936 29930 21992
rect 27521 21934 29930 21936
rect 27521 21931 27587 21934
rect 29200 21858 29800 21934
rect 29870 21858 29930 21934
rect 29200 21798 29930 21858
rect 7892 21792 8208 21793
rect 7892 21728 7898 21792
rect 7962 21728 7978 21792
rect 8042 21728 8058 21792
rect 8122 21728 8138 21792
rect 8202 21728 8208 21792
rect 7892 21727 8208 21728
rect 14838 21792 15154 21793
rect 14838 21728 14844 21792
rect 14908 21728 14924 21792
rect 14988 21728 15004 21792
rect 15068 21728 15084 21792
rect 15148 21728 15154 21792
rect 14838 21727 15154 21728
rect 21784 21792 22100 21793
rect 21784 21728 21790 21792
rect 21854 21728 21870 21792
rect 21934 21728 21950 21792
rect 22014 21728 22030 21792
rect 22094 21728 22100 21792
rect 21784 21727 22100 21728
rect 28730 21792 29046 21793
rect 28730 21728 28736 21792
rect 28800 21728 28816 21792
rect 28880 21728 28896 21792
rect 28960 21728 28976 21792
rect 29040 21728 29046 21792
rect 28730 21727 29046 21728
rect 29200 21708 29800 21798
rect 200 21028 800 21268
rect 4419 21248 4735 21249
rect 4419 21184 4425 21248
rect 4489 21184 4505 21248
rect 4569 21184 4585 21248
rect 4649 21184 4665 21248
rect 4729 21184 4735 21248
rect 4419 21183 4735 21184
rect 11365 21248 11681 21249
rect 11365 21184 11371 21248
rect 11435 21184 11451 21248
rect 11515 21184 11531 21248
rect 11595 21184 11611 21248
rect 11675 21184 11681 21248
rect 11365 21183 11681 21184
rect 18311 21248 18627 21249
rect 18311 21184 18317 21248
rect 18381 21184 18397 21248
rect 18461 21184 18477 21248
rect 18541 21184 18557 21248
rect 18621 21184 18627 21248
rect 18311 21183 18627 21184
rect 25257 21248 25573 21249
rect 25257 21184 25263 21248
rect 25327 21184 25343 21248
rect 25407 21184 25423 21248
rect 25487 21184 25503 21248
rect 25567 21184 25573 21248
rect 25257 21183 25573 21184
rect 28349 21178 28415 21181
rect 29200 21178 29800 21268
rect 28349 21176 29800 21178
rect 28349 21120 28354 21176
rect 28410 21120 29800 21176
rect 28349 21118 29800 21120
rect 28349 21115 28415 21118
rect 29200 21028 29800 21118
rect 7892 20704 8208 20705
rect 7892 20640 7898 20704
rect 7962 20640 7978 20704
rect 8042 20640 8058 20704
rect 8122 20640 8138 20704
rect 8202 20640 8208 20704
rect 7892 20639 8208 20640
rect 14838 20704 15154 20705
rect 14838 20640 14844 20704
rect 14908 20640 14924 20704
rect 14988 20640 15004 20704
rect 15068 20640 15084 20704
rect 15148 20640 15154 20704
rect 14838 20639 15154 20640
rect 21784 20704 22100 20705
rect 21784 20640 21790 20704
rect 21854 20640 21870 20704
rect 21934 20640 21950 20704
rect 22014 20640 22030 20704
rect 22094 20640 22100 20704
rect 21784 20639 22100 20640
rect 28730 20704 29046 20705
rect 28730 20640 28736 20704
rect 28800 20640 28816 20704
rect 28880 20640 28896 20704
rect 28960 20640 28976 20704
rect 29040 20640 29046 20704
rect 28730 20639 29046 20640
rect 200 20348 800 20588
rect 28349 20498 28415 20501
rect 29200 20498 29800 20588
rect 28349 20496 29800 20498
rect 28349 20440 28354 20496
rect 28410 20440 29800 20496
rect 28349 20438 29800 20440
rect 28349 20435 28415 20438
rect 29200 20348 29800 20438
rect 4419 20160 4735 20161
rect 4419 20096 4425 20160
rect 4489 20096 4505 20160
rect 4569 20096 4585 20160
rect 4649 20096 4665 20160
rect 4729 20096 4735 20160
rect 4419 20095 4735 20096
rect 11365 20160 11681 20161
rect 11365 20096 11371 20160
rect 11435 20096 11451 20160
rect 11515 20096 11531 20160
rect 11595 20096 11611 20160
rect 11675 20096 11681 20160
rect 11365 20095 11681 20096
rect 18311 20160 18627 20161
rect 18311 20096 18317 20160
rect 18381 20096 18397 20160
rect 18461 20096 18477 20160
rect 18541 20096 18557 20160
rect 18621 20096 18627 20160
rect 18311 20095 18627 20096
rect 25257 20160 25573 20161
rect 25257 20096 25263 20160
rect 25327 20096 25343 20160
rect 25407 20096 25423 20160
rect 25487 20096 25503 20160
rect 25567 20096 25573 20160
rect 25257 20095 25573 20096
rect 200 19818 800 19908
rect 2773 19818 2839 19821
rect 200 19816 2839 19818
rect 200 19760 2778 19816
rect 2834 19760 2839 19816
rect 200 19758 2839 19760
rect 200 19668 800 19758
rect 2773 19755 2839 19758
rect 26141 19818 26207 19821
rect 29200 19818 29800 19908
rect 26141 19816 29800 19818
rect 26141 19760 26146 19816
rect 26202 19760 29800 19816
rect 26141 19758 29800 19760
rect 26141 19755 26207 19758
rect 29200 19668 29800 19758
rect 7892 19616 8208 19617
rect 7892 19552 7898 19616
rect 7962 19552 7978 19616
rect 8042 19552 8058 19616
rect 8122 19552 8138 19616
rect 8202 19552 8208 19616
rect 7892 19551 8208 19552
rect 14838 19616 15154 19617
rect 14838 19552 14844 19616
rect 14908 19552 14924 19616
rect 14988 19552 15004 19616
rect 15068 19552 15084 19616
rect 15148 19552 15154 19616
rect 14838 19551 15154 19552
rect 21784 19616 22100 19617
rect 21784 19552 21790 19616
rect 21854 19552 21870 19616
rect 21934 19552 21950 19616
rect 22014 19552 22030 19616
rect 22094 19552 22100 19616
rect 21784 19551 22100 19552
rect 28730 19616 29046 19617
rect 28730 19552 28736 19616
rect 28800 19552 28816 19616
rect 28880 19552 28896 19616
rect 28960 19552 28976 19616
rect 29040 19552 29046 19616
rect 28730 19551 29046 19552
rect 200 19138 800 19228
rect 3325 19138 3391 19141
rect 200 19136 3391 19138
rect 200 19080 3330 19136
rect 3386 19080 3391 19136
rect 200 19078 3391 19080
rect 200 18988 800 19078
rect 3325 19075 3391 19078
rect 18689 19138 18755 19141
rect 19149 19138 19215 19141
rect 18689 19136 19215 19138
rect 18689 19080 18694 19136
rect 18750 19080 19154 19136
rect 19210 19080 19215 19136
rect 18689 19078 19215 19080
rect 18689 19075 18755 19078
rect 19149 19075 19215 19078
rect 4419 19072 4735 19073
rect 4419 19008 4425 19072
rect 4489 19008 4505 19072
rect 4569 19008 4585 19072
rect 4649 19008 4665 19072
rect 4729 19008 4735 19072
rect 4419 19007 4735 19008
rect 11365 19072 11681 19073
rect 11365 19008 11371 19072
rect 11435 19008 11451 19072
rect 11515 19008 11531 19072
rect 11595 19008 11611 19072
rect 11675 19008 11681 19072
rect 11365 19007 11681 19008
rect 18311 19072 18627 19073
rect 18311 19008 18317 19072
rect 18381 19008 18397 19072
rect 18461 19008 18477 19072
rect 18541 19008 18557 19072
rect 18621 19008 18627 19072
rect 18311 19007 18627 19008
rect 25257 19072 25573 19073
rect 25257 19008 25263 19072
rect 25327 19008 25343 19072
rect 25407 19008 25423 19072
rect 25487 19008 25503 19072
rect 25567 19008 25573 19072
rect 25257 19007 25573 19008
rect 29200 18988 29800 19228
rect 200 18458 800 18548
rect 7892 18528 8208 18529
rect 7892 18464 7898 18528
rect 7962 18464 7978 18528
rect 8042 18464 8058 18528
rect 8122 18464 8138 18528
rect 8202 18464 8208 18528
rect 7892 18463 8208 18464
rect 14838 18528 15154 18529
rect 14838 18464 14844 18528
rect 14908 18464 14924 18528
rect 14988 18464 15004 18528
rect 15068 18464 15084 18528
rect 15148 18464 15154 18528
rect 14838 18463 15154 18464
rect 21784 18528 22100 18529
rect 21784 18464 21790 18528
rect 21854 18464 21870 18528
rect 21934 18464 21950 18528
rect 22014 18464 22030 18528
rect 22094 18464 22100 18528
rect 21784 18463 22100 18464
rect 28730 18528 29046 18529
rect 28730 18464 28736 18528
rect 28800 18464 28816 18528
rect 28880 18464 28896 18528
rect 28960 18464 28976 18528
rect 29040 18464 29046 18528
rect 28730 18463 29046 18464
rect 1577 18458 1643 18461
rect 200 18456 1643 18458
rect 200 18400 1582 18456
rect 1638 18400 1643 18456
rect 200 18398 1643 18400
rect 200 18308 800 18398
rect 1577 18395 1643 18398
rect 29200 18308 29800 18548
rect 4419 17984 4735 17985
rect 4419 17920 4425 17984
rect 4489 17920 4505 17984
rect 4569 17920 4585 17984
rect 4649 17920 4665 17984
rect 4729 17920 4735 17984
rect 4419 17919 4735 17920
rect 11365 17984 11681 17985
rect 11365 17920 11371 17984
rect 11435 17920 11451 17984
rect 11515 17920 11531 17984
rect 11595 17920 11611 17984
rect 11675 17920 11681 17984
rect 11365 17919 11681 17920
rect 18311 17984 18627 17985
rect 18311 17920 18317 17984
rect 18381 17920 18397 17984
rect 18461 17920 18477 17984
rect 18541 17920 18557 17984
rect 18621 17920 18627 17984
rect 18311 17919 18627 17920
rect 25257 17984 25573 17985
rect 25257 17920 25263 17984
rect 25327 17920 25343 17984
rect 25407 17920 25423 17984
rect 25487 17920 25503 17984
rect 25567 17920 25573 17984
rect 25257 17919 25573 17920
rect 200 17778 800 17868
rect 2773 17778 2839 17781
rect 200 17776 2839 17778
rect 200 17720 2778 17776
rect 2834 17720 2839 17776
rect 200 17718 2839 17720
rect 200 17628 800 17718
rect 2773 17715 2839 17718
rect 29200 17628 29800 17868
rect 7892 17440 8208 17441
rect 7892 17376 7898 17440
rect 7962 17376 7978 17440
rect 8042 17376 8058 17440
rect 8122 17376 8138 17440
rect 8202 17376 8208 17440
rect 7892 17375 8208 17376
rect 14838 17440 15154 17441
rect 14838 17376 14844 17440
rect 14908 17376 14924 17440
rect 14988 17376 15004 17440
rect 15068 17376 15084 17440
rect 15148 17376 15154 17440
rect 14838 17375 15154 17376
rect 21784 17440 22100 17441
rect 21784 17376 21790 17440
rect 21854 17376 21870 17440
rect 21934 17376 21950 17440
rect 22014 17376 22030 17440
rect 22094 17376 22100 17440
rect 21784 17375 22100 17376
rect 28730 17440 29046 17441
rect 28730 17376 28736 17440
rect 28800 17376 28816 17440
rect 28880 17376 28896 17440
rect 28960 17376 28976 17440
rect 29040 17376 29046 17440
rect 28730 17375 29046 17376
rect 200 16948 800 17188
rect 4419 16896 4735 16897
rect 4419 16832 4425 16896
rect 4489 16832 4505 16896
rect 4569 16832 4585 16896
rect 4649 16832 4665 16896
rect 4729 16832 4735 16896
rect 4419 16831 4735 16832
rect 11365 16896 11681 16897
rect 11365 16832 11371 16896
rect 11435 16832 11451 16896
rect 11515 16832 11531 16896
rect 11595 16832 11611 16896
rect 11675 16832 11681 16896
rect 11365 16831 11681 16832
rect 18311 16896 18627 16897
rect 18311 16832 18317 16896
rect 18381 16832 18397 16896
rect 18461 16832 18477 16896
rect 18541 16832 18557 16896
rect 18621 16832 18627 16896
rect 18311 16831 18627 16832
rect 25257 16896 25573 16897
rect 25257 16832 25263 16896
rect 25327 16832 25343 16896
rect 25407 16832 25423 16896
rect 25487 16832 25503 16896
rect 25567 16832 25573 16896
rect 25257 16831 25573 16832
rect 27337 16554 27403 16557
rect 27337 16552 29930 16554
rect 27337 16496 27342 16552
rect 27398 16496 29930 16552
rect 27337 16494 29930 16496
rect 27337 16491 27403 16494
rect 29200 16418 29800 16494
rect 29870 16418 29930 16494
rect 29200 16358 29930 16418
rect 7892 16352 8208 16353
rect 7892 16288 7898 16352
rect 7962 16288 7978 16352
rect 8042 16288 8058 16352
rect 8122 16288 8138 16352
rect 8202 16288 8208 16352
rect 7892 16287 8208 16288
rect 14838 16352 15154 16353
rect 14838 16288 14844 16352
rect 14908 16288 14924 16352
rect 14988 16288 15004 16352
rect 15068 16288 15084 16352
rect 15148 16288 15154 16352
rect 14838 16287 15154 16288
rect 21784 16352 22100 16353
rect 21784 16288 21790 16352
rect 21854 16288 21870 16352
rect 21934 16288 21950 16352
rect 22014 16288 22030 16352
rect 22094 16288 22100 16352
rect 21784 16287 22100 16288
rect 28730 16352 29046 16353
rect 28730 16288 28736 16352
rect 28800 16288 28816 16352
rect 28880 16288 28896 16352
rect 28960 16288 28976 16352
rect 29040 16288 29046 16352
rect 28730 16287 29046 16288
rect 29200 16268 29800 16358
rect 200 15738 800 15828
rect 4419 15808 4735 15809
rect 4419 15744 4425 15808
rect 4489 15744 4505 15808
rect 4569 15744 4585 15808
rect 4649 15744 4665 15808
rect 4729 15744 4735 15808
rect 4419 15743 4735 15744
rect 11365 15808 11681 15809
rect 11365 15744 11371 15808
rect 11435 15744 11451 15808
rect 11515 15744 11531 15808
rect 11595 15744 11611 15808
rect 11675 15744 11681 15808
rect 11365 15743 11681 15744
rect 18311 15808 18627 15809
rect 18311 15744 18317 15808
rect 18381 15744 18397 15808
rect 18461 15744 18477 15808
rect 18541 15744 18557 15808
rect 18621 15744 18627 15808
rect 18311 15743 18627 15744
rect 25257 15808 25573 15809
rect 25257 15744 25263 15808
rect 25327 15744 25343 15808
rect 25407 15744 25423 15808
rect 25487 15744 25503 15808
rect 25567 15744 25573 15808
rect 25257 15743 25573 15744
rect 2773 15738 2839 15741
rect 200 15736 2839 15738
rect 200 15680 2778 15736
rect 2834 15680 2839 15736
rect 200 15678 2839 15680
rect 200 15588 800 15678
rect 2773 15675 2839 15678
rect 27521 15738 27587 15741
rect 29200 15738 29800 15828
rect 27521 15736 29800 15738
rect 27521 15680 27526 15736
rect 27582 15680 29800 15736
rect 27521 15678 29800 15680
rect 27521 15675 27587 15678
rect 29200 15588 29800 15678
rect 7892 15264 8208 15265
rect 7892 15200 7898 15264
rect 7962 15200 7978 15264
rect 8042 15200 8058 15264
rect 8122 15200 8138 15264
rect 8202 15200 8208 15264
rect 7892 15199 8208 15200
rect 14838 15264 15154 15265
rect 14838 15200 14844 15264
rect 14908 15200 14924 15264
rect 14988 15200 15004 15264
rect 15068 15200 15084 15264
rect 15148 15200 15154 15264
rect 14838 15199 15154 15200
rect 21784 15264 22100 15265
rect 21784 15200 21790 15264
rect 21854 15200 21870 15264
rect 21934 15200 21950 15264
rect 22014 15200 22030 15264
rect 22094 15200 22100 15264
rect 21784 15199 22100 15200
rect 28730 15264 29046 15265
rect 28730 15200 28736 15264
rect 28800 15200 28816 15264
rect 28880 15200 28896 15264
rect 28960 15200 28976 15264
rect 29040 15200 29046 15264
rect 28730 15199 29046 15200
rect 200 14908 800 15148
rect 28441 15058 28507 15061
rect 29200 15058 29800 15148
rect 28441 15056 29800 15058
rect 28441 15000 28446 15056
rect 28502 15000 29800 15056
rect 28441 14998 29800 15000
rect 28441 14995 28507 14998
rect 29200 14908 29800 14998
rect 4419 14720 4735 14721
rect 4419 14656 4425 14720
rect 4489 14656 4505 14720
rect 4569 14656 4585 14720
rect 4649 14656 4665 14720
rect 4729 14656 4735 14720
rect 4419 14655 4735 14656
rect 11365 14720 11681 14721
rect 11365 14656 11371 14720
rect 11435 14656 11451 14720
rect 11515 14656 11531 14720
rect 11595 14656 11611 14720
rect 11675 14656 11681 14720
rect 11365 14655 11681 14656
rect 18311 14720 18627 14721
rect 18311 14656 18317 14720
rect 18381 14656 18397 14720
rect 18461 14656 18477 14720
rect 18541 14656 18557 14720
rect 18621 14656 18627 14720
rect 18311 14655 18627 14656
rect 25257 14720 25573 14721
rect 25257 14656 25263 14720
rect 25327 14656 25343 14720
rect 25407 14656 25423 14720
rect 25487 14656 25503 14720
rect 25567 14656 25573 14720
rect 25257 14655 25573 14656
rect 200 14378 800 14468
rect 2773 14378 2839 14381
rect 200 14376 2839 14378
rect 200 14320 2778 14376
rect 2834 14320 2839 14376
rect 200 14318 2839 14320
rect 200 14228 800 14318
rect 2773 14315 2839 14318
rect 28349 14378 28415 14381
rect 29200 14378 29800 14468
rect 28349 14376 29800 14378
rect 28349 14320 28354 14376
rect 28410 14320 29800 14376
rect 28349 14318 29800 14320
rect 28349 14315 28415 14318
rect 29200 14228 29800 14318
rect 7892 14176 8208 14177
rect 7892 14112 7898 14176
rect 7962 14112 7978 14176
rect 8042 14112 8058 14176
rect 8122 14112 8138 14176
rect 8202 14112 8208 14176
rect 7892 14111 8208 14112
rect 14838 14176 15154 14177
rect 14838 14112 14844 14176
rect 14908 14112 14924 14176
rect 14988 14112 15004 14176
rect 15068 14112 15084 14176
rect 15148 14112 15154 14176
rect 14838 14111 15154 14112
rect 21784 14176 22100 14177
rect 21784 14112 21790 14176
rect 21854 14112 21870 14176
rect 21934 14112 21950 14176
rect 22014 14112 22030 14176
rect 22094 14112 22100 14176
rect 21784 14111 22100 14112
rect 28730 14176 29046 14177
rect 28730 14112 28736 14176
rect 28800 14112 28816 14176
rect 28880 14112 28896 14176
rect 28960 14112 28976 14176
rect 29040 14112 29046 14176
rect 28730 14111 29046 14112
rect 200 13698 800 13788
rect 1577 13698 1643 13701
rect 200 13696 1643 13698
rect 200 13640 1582 13696
rect 1638 13640 1643 13696
rect 200 13638 1643 13640
rect 200 13548 800 13638
rect 1577 13635 1643 13638
rect 4419 13632 4735 13633
rect 4419 13568 4425 13632
rect 4489 13568 4505 13632
rect 4569 13568 4585 13632
rect 4649 13568 4665 13632
rect 4729 13568 4735 13632
rect 4419 13567 4735 13568
rect 11365 13632 11681 13633
rect 11365 13568 11371 13632
rect 11435 13568 11451 13632
rect 11515 13568 11531 13632
rect 11595 13568 11611 13632
rect 11675 13568 11681 13632
rect 11365 13567 11681 13568
rect 18311 13632 18627 13633
rect 18311 13568 18317 13632
rect 18381 13568 18397 13632
rect 18461 13568 18477 13632
rect 18541 13568 18557 13632
rect 18621 13568 18627 13632
rect 18311 13567 18627 13568
rect 25257 13632 25573 13633
rect 25257 13568 25263 13632
rect 25327 13568 25343 13632
rect 25407 13568 25423 13632
rect 25487 13568 25503 13632
rect 25567 13568 25573 13632
rect 25257 13567 25573 13568
rect 29200 13548 29800 13788
rect 200 12868 800 13108
rect 7892 13088 8208 13089
rect 7892 13024 7898 13088
rect 7962 13024 7978 13088
rect 8042 13024 8058 13088
rect 8122 13024 8138 13088
rect 8202 13024 8208 13088
rect 7892 13023 8208 13024
rect 14838 13088 15154 13089
rect 14838 13024 14844 13088
rect 14908 13024 14924 13088
rect 14988 13024 15004 13088
rect 15068 13024 15084 13088
rect 15148 13024 15154 13088
rect 14838 13023 15154 13024
rect 21784 13088 22100 13089
rect 21784 13024 21790 13088
rect 21854 13024 21870 13088
rect 21934 13024 21950 13088
rect 22014 13024 22030 13088
rect 22094 13024 22100 13088
rect 21784 13023 22100 13024
rect 28730 13088 29046 13089
rect 28730 13024 28736 13088
rect 28800 13024 28816 13088
rect 28880 13024 28896 13088
rect 28960 13024 28976 13088
rect 29040 13024 29046 13088
rect 28730 13023 29046 13024
rect 29200 12868 29800 13108
rect 4419 12544 4735 12545
rect 4419 12480 4425 12544
rect 4489 12480 4505 12544
rect 4569 12480 4585 12544
rect 4649 12480 4665 12544
rect 4729 12480 4735 12544
rect 4419 12479 4735 12480
rect 11365 12544 11681 12545
rect 11365 12480 11371 12544
rect 11435 12480 11451 12544
rect 11515 12480 11531 12544
rect 11595 12480 11611 12544
rect 11675 12480 11681 12544
rect 11365 12479 11681 12480
rect 18311 12544 18627 12545
rect 18311 12480 18317 12544
rect 18381 12480 18397 12544
rect 18461 12480 18477 12544
rect 18541 12480 18557 12544
rect 18621 12480 18627 12544
rect 18311 12479 18627 12480
rect 25257 12544 25573 12545
rect 25257 12480 25263 12544
rect 25327 12480 25343 12544
rect 25407 12480 25423 12544
rect 25487 12480 25503 12544
rect 25567 12480 25573 12544
rect 25257 12479 25573 12480
rect 200 12338 800 12428
rect 3601 12338 3667 12341
rect 200 12336 3667 12338
rect 200 12280 3606 12336
rect 3662 12280 3667 12336
rect 200 12278 3667 12280
rect 200 12188 800 12278
rect 3601 12275 3667 12278
rect 28349 12338 28415 12341
rect 29200 12338 29800 12428
rect 28349 12336 29800 12338
rect 28349 12280 28354 12336
rect 28410 12280 29800 12336
rect 28349 12278 29800 12280
rect 28349 12275 28415 12278
rect 29200 12188 29800 12278
rect 7892 12000 8208 12001
rect 7892 11936 7898 12000
rect 7962 11936 7978 12000
rect 8042 11936 8058 12000
rect 8122 11936 8138 12000
rect 8202 11936 8208 12000
rect 7892 11935 8208 11936
rect 14838 12000 15154 12001
rect 14838 11936 14844 12000
rect 14908 11936 14924 12000
rect 14988 11936 15004 12000
rect 15068 11936 15084 12000
rect 15148 11936 15154 12000
rect 14838 11935 15154 11936
rect 21784 12000 22100 12001
rect 21784 11936 21790 12000
rect 21854 11936 21870 12000
rect 21934 11936 21950 12000
rect 22014 11936 22030 12000
rect 22094 11936 22100 12000
rect 21784 11935 22100 11936
rect 28730 12000 29046 12001
rect 28730 11936 28736 12000
rect 28800 11936 28816 12000
rect 28880 11936 28896 12000
rect 28960 11936 28976 12000
rect 29040 11936 29046 12000
rect 28730 11935 29046 11936
rect 200 11658 800 11748
rect 2773 11658 2839 11661
rect 200 11656 2839 11658
rect 200 11600 2778 11656
rect 2834 11600 2839 11656
rect 200 11598 2839 11600
rect 200 11508 800 11598
rect 2773 11595 2839 11598
rect 4419 11456 4735 11457
rect 4419 11392 4425 11456
rect 4489 11392 4505 11456
rect 4569 11392 4585 11456
rect 4649 11392 4665 11456
rect 4729 11392 4735 11456
rect 4419 11391 4735 11392
rect 11365 11456 11681 11457
rect 11365 11392 11371 11456
rect 11435 11392 11451 11456
rect 11515 11392 11531 11456
rect 11595 11392 11611 11456
rect 11675 11392 11681 11456
rect 11365 11391 11681 11392
rect 18311 11456 18627 11457
rect 18311 11392 18317 11456
rect 18381 11392 18397 11456
rect 18461 11392 18477 11456
rect 18541 11392 18557 11456
rect 18621 11392 18627 11456
rect 18311 11391 18627 11392
rect 25257 11456 25573 11457
rect 25257 11392 25263 11456
rect 25327 11392 25343 11456
rect 25407 11392 25423 11456
rect 25487 11392 25503 11456
rect 25567 11392 25573 11456
rect 25257 11391 25573 11392
rect 29200 10978 29800 11068
rect 29913 10978 29979 10981
rect 29200 10976 29979 10978
rect 29200 10920 29918 10976
rect 29974 10920 29979 10976
rect 29200 10918 29979 10920
rect 7892 10912 8208 10913
rect 7892 10848 7898 10912
rect 7962 10848 7978 10912
rect 8042 10848 8058 10912
rect 8122 10848 8138 10912
rect 8202 10848 8208 10912
rect 7892 10847 8208 10848
rect 14838 10912 15154 10913
rect 14838 10848 14844 10912
rect 14908 10848 14924 10912
rect 14988 10848 15004 10912
rect 15068 10848 15084 10912
rect 15148 10848 15154 10912
rect 14838 10847 15154 10848
rect 21784 10912 22100 10913
rect 21784 10848 21790 10912
rect 21854 10848 21870 10912
rect 21934 10848 21950 10912
rect 22014 10848 22030 10912
rect 22094 10848 22100 10912
rect 21784 10847 22100 10848
rect 28730 10912 29046 10913
rect 28730 10848 28736 10912
rect 28800 10848 28816 10912
rect 28880 10848 28896 10912
rect 28960 10848 28976 10912
rect 29040 10848 29046 10912
rect 28730 10847 29046 10848
rect 29200 10828 29800 10918
rect 29913 10915 29979 10918
rect 200 10148 800 10388
rect 4419 10368 4735 10369
rect 4419 10304 4425 10368
rect 4489 10304 4505 10368
rect 4569 10304 4585 10368
rect 4649 10304 4665 10368
rect 4729 10304 4735 10368
rect 4419 10303 4735 10304
rect 11365 10368 11681 10369
rect 11365 10304 11371 10368
rect 11435 10304 11451 10368
rect 11515 10304 11531 10368
rect 11595 10304 11611 10368
rect 11675 10304 11681 10368
rect 11365 10303 11681 10304
rect 18311 10368 18627 10369
rect 18311 10304 18317 10368
rect 18381 10304 18397 10368
rect 18461 10304 18477 10368
rect 18541 10304 18557 10368
rect 18621 10304 18627 10368
rect 18311 10303 18627 10304
rect 25257 10368 25573 10369
rect 25257 10304 25263 10368
rect 25327 10304 25343 10368
rect 25407 10304 25423 10368
rect 25487 10304 25503 10368
rect 25567 10304 25573 10368
rect 25257 10303 25573 10304
rect 27521 10298 27587 10301
rect 29200 10298 29800 10388
rect 27521 10296 29800 10298
rect 27521 10240 27526 10296
rect 27582 10240 29800 10296
rect 27521 10238 29800 10240
rect 27521 10235 27587 10238
rect 29200 10148 29800 10238
rect 7892 9824 8208 9825
rect 7892 9760 7898 9824
rect 7962 9760 7978 9824
rect 8042 9760 8058 9824
rect 8122 9760 8138 9824
rect 8202 9760 8208 9824
rect 7892 9759 8208 9760
rect 14838 9824 15154 9825
rect 14838 9760 14844 9824
rect 14908 9760 14924 9824
rect 14988 9760 15004 9824
rect 15068 9760 15084 9824
rect 15148 9760 15154 9824
rect 14838 9759 15154 9760
rect 21784 9824 22100 9825
rect 21784 9760 21790 9824
rect 21854 9760 21870 9824
rect 21934 9760 21950 9824
rect 22014 9760 22030 9824
rect 22094 9760 22100 9824
rect 21784 9759 22100 9760
rect 28730 9824 29046 9825
rect 28730 9760 28736 9824
rect 28800 9760 28816 9824
rect 28880 9760 28896 9824
rect 28960 9760 28976 9824
rect 29040 9760 29046 9824
rect 28730 9759 29046 9760
rect 200 9468 800 9708
rect 29200 9468 29800 9708
rect 4419 9280 4735 9281
rect 4419 9216 4425 9280
rect 4489 9216 4505 9280
rect 4569 9216 4585 9280
rect 4649 9216 4665 9280
rect 4729 9216 4735 9280
rect 4419 9215 4735 9216
rect 11365 9280 11681 9281
rect 11365 9216 11371 9280
rect 11435 9216 11451 9280
rect 11515 9216 11531 9280
rect 11595 9216 11611 9280
rect 11675 9216 11681 9280
rect 11365 9215 11681 9216
rect 18311 9280 18627 9281
rect 18311 9216 18317 9280
rect 18381 9216 18397 9280
rect 18461 9216 18477 9280
rect 18541 9216 18557 9280
rect 18621 9216 18627 9280
rect 18311 9215 18627 9216
rect 25257 9280 25573 9281
rect 25257 9216 25263 9280
rect 25327 9216 25343 9280
rect 25407 9216 25423 9280
rect 25487 9216 25503 9280
rect 25567 9216 25573 9280
rect 25257 9215 25573 9216
rect 200 8938 800 9028
rect 2773 8938 2839 8941
rect 200 8936 2839 8938
rect 200 8880 2778 8936
rect 2834 8880 2839 8936
rect 200 8878 2839 8880
rect 200 8788 800 8878
rect 2773 8875 2839 8878
rect 27521 8938 27587 8941
rect 29200 8938 29800 9028
rect 27521 8936 29800 8938
rect 27521 8880 27526 8936
rect 27582 8880 29800 8936
rect 27521 8878 29800 8880
rect 27521 8875 27587 8878
rect 29200 8788 29800 8878
rect 7892 8736 8208 8737
rect 7892 8672 7898 8736
rect 7962 8672 7978 8736
rect 8042 8672 8058 8736
rect 8122 8672 8138 8736
rect 8202 8672 8208 8736
rect 7892 8671 8208 8672
rect 14838 8736 15154 8737
rect 14838 8672 14844 8736
rect 14908 8672 14924 8736
rect 14988 8672 15004 8736
rect 15068 8672 15084 8736
rect 15148 8672 15154 8736
rect 14838 8671 15154 8672
rect 21784 8736 22100 8737
rect 21784 8672 21790 8736
rect 21854 8672 21870 8736
rect 21934 8672 21950 8736
rect 22014 8672 22030 8736
rect 22094 8672 22100 8736
rect 21784 8671 22100 8672
rect 28730 8736 29046 8737
rect 28730 8672 28736 8736
rect 28800 8672 28816 8736
rect 28880 8672 28896 8736
rect 28960 8672 28976 8736
rect 29040 8672 29046 8736
rect 28730 8671 29046 8672
rect 200 8258 800 8348
rect 4061 8258 4127 8261
rect 200 8256 4127 8258
rect 200 8200 4066 8256
rect 4122 8200 4127 8256
rect 200 8198 4127 8200
rect 200 8108 800 8198
rect 4061 8195 4127 8198
rect 26141 8258 26207 8261
rect 29200 8258 29800 8348
rect 26141 8256 29800 8258
rect 26141 8200 26146 8256
rect 26202 8200 29800 8256
rect 26141 8198 29800 8200
rect 26141 8195 26207 8198
rect 4419 8192 4735 8193
rect 4419 8128 4425 8192
rect 4489 8128 4505 8192
rect 4569 8128 4585 8192
rect 4649 8128 4665 8192
rect 4729 8128 4735 8192
rect 4419 8127 4735 8128
rect 11365 8192 11681 8193
rect 11365 8128 11371 8192
rect 11435 8128 11451 8192
rect 11515 8128 11531 8192
rect 11595 8128 11611 8192
rect 11675 8128 11681 8192
rect 11365 8127 11681 8128
rect 18311 8192 18627 8193
rect 18311 8128 18317 8192
rect 18381 8128 18397 8192
rect 18461 8128 18477 8192
rect 18541 8128 18557 8192
rect 18621 8128 18627 8192
rect 18311 8127 18627 8128
rect 25257 8192 25573 8193
rect 25257 8128 25263 8192
rect 25327 8128 25343 8192
rect 25407 8128 25423 8192
rect 25487 8128 25503 8192
rect 25567 8128 25573 8192
rect 25257 8127 25573 8128
rect 29200 8108 29800 8198
rect 200 7578 800 7668
rect 7892 7648 8208 7649
rect 7892 7584 7898 7648
rect 7962 7584 7978 7648
rect 8042 7584 8058 7648
rect 8122 7584 8138 7648
rect 8202 7584 8208 7648
rect 7892 7583 8208 7584
rect 14838 7648 15154 7649
rect 14838 7584 14844 7648
rect 14908 7584 14924 7648
rect 14988 7584 15004 7648
rect 15068 7584 15084 7648
rect 15148 7584 15154 7648
rect 14838 7583 15154 7584
rect 21784 7648 22100 7649
rect 21784 7584 21790 7648
rect 21854 7584 21870 7648
rect 21934 7584 21950 7648
rect 22014 7584 22030 7648
rect 22094 7584 22100 7648
rect 21784 7583 22100 7584
rect 28730 7648 29046 7649
rect 28730 7584 28736 7648
rect 28800 7584 28816 7648
rect 28880 7584 28896 7648
rect 28960 7584 28976 7648
rect 29040 7584 29046 7648
rect 28730 7583 29046 7584
rect 2773 7578 2839 7581
rect 200 7576 2839 7578
rect 200 7520 2778 7576
rect 2834 7520 2839 7576
rect 200 7518 2839 7520
rect 200 7428 800 7518
rect 2773 7515 2839 7518
rect 29200 7578 29800 7668
rect 29913 7578 29979 7581
rect 29200 7576 29979 7578
rect 29200 7520 29918 7576
rect 29974 7520 29979 7576
rect 29200 7518 29979 7520
rect 29200 7428 29800 7518
rect 29913 7515 29979 7518
rect 4419 7104 4735 7105
rect 4419 7040 4425 7104
rect 4489 7040 4505 7104
rect 4569 7040 4585 7104
rect 4649 7040 4665 7104
rect 4729 7040 4735 7104
rect 4419 7039 4735 7040
rect 11365 7104 11681 7105
rect 11365 7040 11371 7104
rect 11435 7040 11451 7104
rect 11515 7040 11531 7104
rect 11595 7040 11611 7104
rect 11675 7040 11681 7104
rect 11365 7039 11681 7040
rect 18311 7104 18627 7105
rect 18311 7040 18317 7104
rect 18381 7040 18397 7104
rect 18461 7040 18477 7104
rect 18541 7040 18557 7104
rect 18621 7040 18627 7104
rect 18311 7039 18627 7040
rect 25257 7104 25573 7105
rect 25257 7040 25263 7104
rect 25327 7040 25343 7104
rect 25407 7040 25423 7104
rect 25487 7040 25503 7104
rect 25567 7040 25573 7104
rect 25257 7039 25573 7040
rect 200 6748 800 6988
rect 26141 6898 26207 6901
rect 29200 6898 29800 6988
rect 26141 6896 29800 6898
rect 26141 6840 26146 6896
rect 26202 6840 29800 6896
rect 26141 6838 29800 6840
rect 26141 6835 26207 6838
rect 29200 6748 29800 6838
rect 7892 6560 8208 6561
rect 7892 6496 7898 6560
rect 7962 6496 7978 6560
rect 8042 6496 8058 6560
rect 8122 6496 8138 6560
rect 8202 6496 8208 6560
rect 7892 6495 8208 6496
rect 14838 6560 15154 6561
rect 14838 6496 14844 6560
rect 14908 6496 14924 6560
rect 14988 6496 15004 6560
rect 15068 6496 15084 6560
rect 15148 6496 15154 6560
rect 14838 6495 15154 6496
rect 21784 6560 22100 6561
rect 21784 6496 21790 6560
rect 21854 6496 21870 6560
rect 21934 6496 21950 6560
rect 22014 6496 22030 6560
rect 22094 6496 22100 6560
rect 21784 6495 22100 6496
rect 28730 6560 29046 6561
rect 28730 6496 28736 6560
rect 28800 6496 28816 6560
rect 28880 6496 28896 6560
rect 28960 6496 28976 6560
rect 29040 6496 29046 6560
rect 28730 6495 29046 6496
rect 200 6218 800 6308
rect 3601 6218 3667 6221
rect 200 6216 3667 6218
rect 200 6160 3606 6216
rect 3662 6160 3667 6216
rect 200 6158 3667 6160
rect 200 6068 800 6158
rect 3601 6155 3667 6158
rect 4419 6016 4735 6017
rect 4419 5952 4425 6016
rect 4489 5952 4505 6016
rect 4569 5952 4585 6016
rect 4649 5952 4665 6016
rect 4729 5952 4735 6016
rect 4419 5951 4735 5952
rect 11365 6016 11681 6017
rect 11365 5952 11371 6016
rect 11435 5952 11451 6016
rect 11515 5952 11531 6016
rect 11595 5952 11611 6016
rect 11675 5952 11681 6016
rect 11365 5951 11681 5952
rect 18311 6016 18627 6017
rect 18311 5952 18317 6016
rect 18381 5952 18397 6016
rect 18461 5952 18477 6016
rect 18541 5952 18557 6016
rect 18621 5952 18627 6016
rect 18311 5951 18627 5952
rect 25257 6016 25573 6017
rect 25257 5952 25263 6016
rect 25327 5952 25343 6016
rect 25407 5952 25423 6016
rect 25487 5952 25503 6016
rect 25567 5952 25573 6016
rect 25257 5951 25573 5952
rect 29200 5538 29800 5628
rect 29913 5538 29979 5541
rect 29200 5536 29979 5538
rect 29200 5480 29918 5536
rect 29974 5480 29979 5536
rect 29200 5478 29979 5480
rect 7892 5472 8208 5473
rect 7892 5408 7898 5472
rect 7962 5408 7978 5472
rect 8042 5408 8058 5472
rect 8122 5408 8138 5472
rect 8202 5408 8208 5472
rect 7892 5407 8208 5408
rect 14838 5472 15154 5473
rect 14838 5408 14844 5472
rect 14908 5408 14924 5472
rect 14988 5408 15004 5472
rect 15068 5408 15084 5472
rect 15148 5408 15154 5472
rect 14838 5407 15154 5408
rect 21784 5472 22100 5473
rect 21784 5408 21790 5472
rect 21854 5408 21870 5472
rect 21934 5408 21950 5472
rect 22014 5408 22030 5472
rect 22094 5408 22100 5472
rect 21784 5407 22100 5408
rect 28730 5472 29046 5473
rect 28730 5408 28736 5472
rect 28800 5408 28816 5472
rect 28880 5408 28896 5472
rect 28960 5408 28976 5472
rect 29040 5408 29046 5472
rect 28730 5407 29046 5408
rect 29200 5388 29800 5478
rect 29913 5475 29979 5478
rect 200 4858 800 4948
rect 4419 4928 4735 4929
rect 4419 4864 4425 4928
rect 4489 4864 4505 4928
rect 4569 4864 4585 4928
rect 4649 4864 4665 4928
rect 4729 4864 4735 4928
rect 4419 4863 4735 4864
rect 11365 4928 11681 4929
rect 11365 4864 11371 4928
rect 11435 4864 11451 4928
rect 11515 4864 11531 4928
rect 11595 4864 11611 4928
rect 11675 4864 11681 4928
rect 11365 4863 11681 4864
rect 18311 4928 18627 4929
rect 18311 4864 18317 4928
rect 18381 4864 18397 4928
rect 18461 4864 18477 4928
rect 18541 4864 18557 4928
rect 18621 4864 18627 4928
rect 18311 4863 18627 4864
rect 25257 4928 25573 4929
rect 25257 4864 25263 4928
rect 25327 4864 25343 4928
rect 25407 4864 25423 4928
rect 25487 4864 25503 4928
rect 25567 4864 25573 4928
rect 25257 4863 25573 4864
rect 2773 4858 2839 4861
rect 200 4856 2839 4858
rect 200 4800 2778 4856
rect 2834 4800 2839 4856
rect 200 4798 2839 4800
rect 200 4708 800 4798
rect 2773 4795 2839 4798
rect 29200 4708 29800 4948
rect 7892 4384 8208 4385
rect 7892 4320 7898 4384
rect 7962 4320 7978 4384
rect 8042 4320 8058 4384
rect 8122 4320 8138 4384
rect 8202 4320 8208 4384
rect 7892 4319 8208 4320
rect 14838 4384 15154 4385
rect 14838 4320 14844 4384
rect 14908 4320 14924 4384
rect 14988 4320 15004 4384
rect 15068 4320 15084 4384
rect 15148 4320 15154 4384
rect 14838 4319 15154 4320
rect 21784 4384 22100 4385
rect 21784 4320 21790 4384
rect 21854 4320 21870 4384
rect 21934 4320 21950 4384
rect 22014 4320 22030 4384
rect 22094 4320 22100 4384
rect 21784 4319 22100 4320
rect 28730 4384 29046 4385
rect 28730 4320 28736 4384
rect 28800 4320 28816 4384
rect 28880 4320 28896 4384
rect 28960 4320 28976 4384
rect 29040 4320 29046 4384
rect 28730 4319 29046 4320
rect 200 4178 800 4268
rect 4061 4178 4127 4181
rect 200 4176 4127 4178
rect 200 4120 4066 4176
rect 4122 4120 4127 4176
rect 200 4118 4127 4120
rect 200 4028 800 4118
rect 4061 4115 4127 4118
rect 29200 4028 29800 4268
rect 4419 3840 4735 3841
rect 4419 3776 4425 3840
rect 4489 3776 4505 3840
rect 4569 3776 4585 3840
rect 4649 3776 4665 3840
rect 4729 3776 4735 3840
rect 4419 3775 4735 3776
rect 11365 3840 11681 3841
rect 11365 3776 11371 3840
rect 11435 3776 11451 3840
rect 11515 3776 11531 3840
rect 11595 3776 11611 3840
rect 11675 3776 11681 3840
rect 11365 3775 11681 3776
rect 18311 3840 18627 3841
rect 18311 3776 18317 3840
rect 18381 3776 18397 3840
rect 18461 3776 18477 3840
rect 18541 3776 18557 3840
rect 18621 3776 18627 3840
rect 18311 3775 18627 3776
rect 25257 3840 25573 3841
rect 25257 3776 25263 3840
rect 25327 3776 25343 3840
rect 25407 3776 25423 3840
rect 25487 3776 25503 3840
rect 25567 3776 25573 3840
rect 25257 3775 25573 3776
rect 200 3498 800 3588
rect 3049 3498 3115 3501
rect 200 3496 3115 3498
rect 200 3440 3054 3496
rect 3110 3440 3115 3496
rect 200 3438 3115 3440
rect 200 3348 800 3438
rect 3049 3435 3115 3438
rect 27429 3498 27495 3501
rect 29200 3498 29800 3588
rect 27429 3496 29800 3498
rect 27429 3440 27434 3496
rect 27490 3440 29800 3496
rect 27429 3438 29800 3440
rect 27429 3435 27495 3438
rect 29200 3348 29800 3438
rect 7892 3296 8208 3297
rect 7892 3232 7898 3296
rect 7962 3232 7978 3296
rect 8042 3232 8058 3296
rect 8122 3232 8138 3296
rect 8202 3232 8208 3296
rect 7892 3231 8208 3232
rect 14838 3296 15154 3297
rect 14838 3232 14844 3296
rect 14908 3232 14924 3296
rect 14988 3232 15004 3296
rect 15068 3232 15084 3296
rect 15148 3232 15154 3296
rect 14838 3231 15154 3232
rect 21784 3296 22100 3297
rect 21784 3232 21790 3296
rect 21854 3232 21870 3296
rect 21934 3232 21950 3296
rect 22014 3232 22030 3296
rect 22094 3232 22100 3296
rect 21784 3231 22100 3232
rect 28730 3296 29046 3297
rect 28730 3232 28736 3296
rect 28800 3232 28816 3296
rect 28880 3232 28896 3296
rect 28960 3232 28976 3296
rect 29040 3232 29046 3296
rect 28730 3231 29046 3232
rect 200 2818 800 2908
rect 2865 2818 2931 2821
rect 200 2816 2931 2818
rect 200 2760 2870 2816
rect 2926 2760 2931 2816
rect 200 2758 2931 2760
rect 200 2668 800 2758
rect 2865 2755 2931 2758
rect 26141 2818 26207 2821
rect 29200 2818 29800 2908
rect 26141 2816 29800 2818
rect 26141 2760 26146 2816
rect 26202 2760 29800 2816
rect 26141 2758 29800 2760
rect 26141 2755 26207 2758
rect 4419 2752 4735 2753
rect 4419 2688 4425 2752
rect 4489 2688 4505 2752
rect 4569 2688 4585 2752
rect 4649 2688 4665 2752
rect 4729 2688 4735 2752
rect 4419 2687 4735 2688
rect 11365 2752 11681 2753
rect 11365 2688 11371 2752
rect 11435 2688 11451 2752
rect 11515 2688 11531 2752
rect 11595 2688 11611 2752
rect 11675 2688 11681 2752
rect 11365 2687 11681 2688
rect 18311 2752 18627 2753
rect 18311 2688 18317 2752
rect 18381 2688 18397 2752
rect 18461 2688 18477 2752
rect 18541 2688 18557 2752
rect 18621 2688 18627 2752
rect 18311 2687 18627 2688
rect 25257 2752 25573 2753
rect 25257 2688 25263 2752
rect 25327 2688 25343 2752
rect 25407 2688 25423 2752
rect 25487 2688 25503 2752
rect 25567 2688 25573 2752
rect 25257 2687 25573 2688
rect 29200 2668 29800 2758
rect 28073 2546 28139 2549
rect 28073 2544 29378 2546
rect 28073 2488 28078 2544
rect 28134 2488 29378 2544
rect 28073 2486 29378 2488
rect 28073 2483 28139 2486
rect 29318 2274 29378 2486
rect 29318 2228 29930 2274
rect 200 2138 800 2228
rect 29200 2214 29930 2228
rect 7892 2208 8208 2209
rect 7892 2144 7898 2208
rect 7962 2144 7978 2208
rect 8042 2144 8058 2208
rect 8122 2144 8138 2208
rect 8202 2144 8208 2208
rect 7892 2143 8208 2144
rect 14838 2208 15154 2209
rect 14838 2144 14844 2208
rect 14908 2144 14924 2208
rect 14988 2144 15004 2208
rect 15068 2144 15084 2208
rect 15148 2144 15154 2208
rect 14838 2143 15154 2144
rect 21784 2208 22100 2209
rect 21784 2144 21790 2208
rect 21854 2144 21870 2208
rect 21934 2144 21950 2208
rect 22014 2144 22030 2208
rect 22094 2144 22100 2208
rect 21784 2143 22100 2144
rect 28730 2208 29046 2209
rect 28730 2144 28736 2208
rect 28800 2144 28816 2208
rect 28880 2144 28896 2208
rect 28960 2144 28976 2208
rect 29040 2144 29046 2208
rect 28730 2143 29046 2144
rect 3509 2138 3575 2141
rect 200 2136 3575 2138
rect 200 2080 3514 2136
rect 3570 2080 3575 2136
rect 200 2078 3575 2080
rect 200 1988 800 2078
rect 3509 2075 3575 2078
rect 29200 2138 29800 2214
rect 29870 2138 29930 2214
rect 29200 2078 29930 2138
rect 29200 1988 29800 2078
rect 200 1458 800 1548
rect 2773 1458 2839 1461
rect 200 1456 2839 1458
rect 200 1400 2778 1456
rect 2834 1400 2839 1456
rect 200 1398 2839 1400
rect 200 1308 800 1398
rect 2773 1395 2839 1398
rect 27521 1458 27587 1461
rect 29200 1458 29800 1548
rect 27521 1456 29800 1458
rect 27521 1400 27526 1456
rect 27582 1400 29800 1456
rect 27521 1398 29800 1400
rect 27521 1395 27587 1398
rect 29200 1308 29800 1398
rect 200 628 800 868
rect 29200 -52 29800 188
<< via3 >>
rect 4425 47356 4489 47360
rect 4425 47300 4429 47356
rect 4429 47300 4485 47356
rect 4485 47300 4489 47356
rect 4425 47296 4489 47300
rect 4505 47356 4569 47360
rect 4505 47300 4509 47356
rect 4509 47300 4565 47356
rect 4565 47300 4569 47356
rect 4505 47296 4569 47300
rect 4585 47356 4649 47360
rect 4585 47300 4589 47356
rect 4589 47300 4645 47356
rect 4645 47300 4649 47356
rect 4585 47296 4649 47300
rect 4665 47356 4729 47360
rect 4665 47300 4669 47356
rect 4669 47300 4725 47356
rect 4725 47300 4729 47356
rect 4665 47296 4729 47300
rect 11371 47356 11435 47360
rect 11371 47300 11375 47356
rect 11375 47300 11431 47356
rect 11431 47300 11435 47356
rect 11371 47296 11435 47300
rect 11451 47356 11515 47360
rect 11451 47300 11455 47356
rect 11455 47300 11511 47356
rect 11511 47300 11515 47356
rect 11451 47296 11515 47300
rect 11531 47356 11595 47360
rect 11531 47300 11535 47356
rect 11535 47300 11591 47356
rect 11591 47300 11595 47356
rect 11531 47296 11595 47300
rect 11611 47356 11675 47360
rect 11611 47300 11615 47356
rect 11615 47300 11671 47356
rect 11671 47300 11675 47356
rect 11611 47296 11675 47300
rect 18317 47356 18381 47360
rect 18317 47300 18321 47356
rect 18321 47300 18377 47356
rect 18377 47300 18381 47356
rect 18317 47296 18381 47300
rect 18397 47356 18461 47360
rect 18397 47300 18401 47356
rect 18401 47300 18457 47356
rect 18457 47300 18461 47356
rect 18397 47296 18461 47300
rect 18477 47356 18541 47360
rect 18477 47300 18481 47356
rect 18481 47300 18537 47356
rect 18537 47300 18541 47356
rect 18477 47296 18541 47300
rect 18557 47356 18621 47360
rect 18557 47300 18561 47356
rect 18561 47300 18617 47356
rect 18617 47300 18621 47356
rect 18557 47296 18621 47300
rect 25263 47356 25327 47360
rect 25263 47300 25267 47356
rect 25267 47300 25323 47356
rect 25323 47300 25327 47356
rect 25263 47296 25327 47300
rect 25343 47356 25407 47360
rect 25343 47300 25347 47356
rect 25347 47300 25403 47356
rect 25403 47300 25407 47356
rect 25343 47296 25407 47300
rect 25423 47356 25487 47360
rect 25423 47300 25427 47356
rect 25427 47300 25483 47356
rect 25483 47300 25487 47356
rect 25423 47296 25487 47300
rect 25503 47356 25567 47360
rect 25503 47300 25507 47356
rect 25507 47300 25563 47356
rect 25563 47300 25567 47356
rect 25503 47296 25567 47300
rect 7898 46812 7962 46816
rect 7898 46756 7902 46812
rect 7902 46756 7958 46812
rect 7958 46756 7962 46812
rect 7898 46752 7962 46756
rect 7978 46812 8042 46816
rect 7978 46756 7982 46812
rect 7982 46756 8038 46812
rect 8038 46756 8042 46812
rect 7978 46752 8042 46756
rect 8058 46812 8122 46816
rect 8058 46756 8062 46812
rect 8062 46756 8118 46812
rect 8118 46756 8122 46812
rect 8058 46752 8122 46756
rect 8138 46812 8202 46816
rect 8138 46756 8142 46812
rect 8142 46756 8198 46812
rect 8198 46756 8202 46812
rect 8138 46752 8202 46756
rect 14844 46812 14908 46816
rect 14844 46756 14848 46812
rect 14848 46756 14904 46812
rect 14904 46756 14908 46812
rect 14844 46752 14908 46756
rect 14924 46812 14988 46816
rect 14924 46756 14928 46812
rect 14928 46756 14984 46812
rect 14984 46756 14988 46812
rect 14924 46752 14988 46756
rect 15004 46812 15068 46816
rect 15004 46756 15008 46812
rect 15008 46756 15064 46812
rect 15064 46756 15068 46812
rect 15004 46752 15068 46756
rect 15084 46812 15148 46816
rect 15084 46756 15088 46812
rect 15088 46756 15144 46812
rect 15144 46756 15148 46812
rect 15084 46752 15148 46756
rect 21790 46812 21854 46816
rect 21790 46756 21794 46812
rect 21794 46756 21850 46812
rect 21850 46756 21854 46812
rect 21790 46752 21854 46756
rect 21870 46812 21934 46816
rect 21870 46756 21874 46812
rect 21874 46756 21930 46812
rect 21930 46756 21934 46812
rect 21870 46752 21934 46756
rect 21950 46812 22014 46816
rect 21950 46756 21954 46812
rect 21954 46756 22010 46812
rect 22010 46756 22014 46812
rect 21950 46752 22014 46756
rect 22030 46812 22094 46816
rect 22030 46756 22034 46812
rect 22034 46756 22090 46812
rect 22090 46756 22094 46812
rect 22030 46752 22094 46756
rect 28736 46812 28800 46816
rect 28736 46756 28740 46812
rect 28740 46756 28796 46812
rect 28796 46756 28800 46812
rect 28736 46752 28800 46756
rect 28816 46812 28880 46816
rect 28816 46756 28820 46812
rect 28820 46756 28876 46812
rect 28876 46756 28880 46812
rect 28816 46752 28880 46756
rect 28896 46812 28960 46816
rect 28896 46756 28900 46812
rect 28900 46756 28956 46812
rect 28956 46756 28960 46812
rect 28896 46752 28960 46756
rect 28976 46812 29040 46816
rect 28976 46756 28980 46812
rect 28980 46756 29036 46812
rect 29036 46756 29040 46812
rect 28976 46752 29040 46756
rect 4425 46268 4489 46272
rect 4425 46212 4429 46268
rect 4429 46212 4485 46268
rect 4485 46212 4489 46268
rect 4425 46208 4489 46212
rect 4505 46268 4569 46272
rect 4505 46212 4509 46268
rect 4509 46212 4565 46268
rect 4565 46212 4569 46268
rect 4505 46208 4569 46212
rect 4585 46268 4649 46272
rect 4585 46212 4589 46268
rect 4589 46212 4645 46268
rect 4645 46212 4649 46268
rect 4585 46208 4649 46212
rect 4665 46268 4729 46272
rect 4665 46212 4669 46268
rect 4669 46212 4725 46268
rect 4725 46212 4729 46268
rect 4665 46208 4729 46212
rect 11371 46268 11435 46272
rect 11371 46212 11375 46268
rect 11375 46212 11431 46268
rect 11431 46212 11435 46268
rect 11371 46208 11435 46212
rect 11451 46268 11515 46272
rect 11451 46212 11455 46268
rect 11455 46212 11511 46268
rect 11511 46212 11515 46268
rect 11451 46208 11515 46212
rect 11531 46268 11595 46272
rect 11531 46212 11535 46268
rect 11535 46212 11591 46268
rect 11591 46212 11595 46268
rect 11531 46208 11595 46212
rect 11611 46268 11675 46272
rect 11611 46212 11615 46268
rect 11615 46212 11671 46268
rect 11671 46212 11675 46268
rect 11611 46208 11675 46212
rect 18317 46268 18381 46272
rect 18317 46212 18321 46268
rect 18321 46212 18377 46268
rect 18377 46212 18381 46268
rect 18317 46208 18381 46212
rect 18397 46268 18461 46272
rect 18397 46212 18401 46268
rect 18401 46212 18457 46268
rect 18457 46212 18461 46268
rect 18397 46208 18461 46212
rect 18477 46268 18541 46272
rect 18477 46212 18481 46268
rect 18481 46212 18537 46268
rect 18537 46212 18541 46268
rect 18477 46208 18541 46212
rect 18557 46268 18621 46272
rect 18557 46212 18561 46268
rect 18561 46212 18617 46268
rect 18617 46212 18621 46268
rect 18557 46208 18621 46212
rect 25263 46268 25327 46272
rect 25263 46212 25267 46268
rect 25267 46212 25323 46268
rect 25323 46212 25327 46268
rect 25263 46208 25327 46212
rect 25343 46268 25407 46272
rect 25343 46212 25347 46268
rect 25347 46212 25403 46268
rect 25403 46212 25407 46268
rect 25343 46208 25407 46212
rect 25423 46268 25487 46272
rect 25423 46212 25427 46268
rect 25427 46212 25483 46268
rect 25483 46212 25487 46268
rect 25423 46208 25487 46212
rect 25503 46268 25567 46272
rect 25503 46212 25507 46268
rect 25507 46212 25563 46268
rect 25563 46212 25567 46268
rect 25503 46208 25567 46212
rect 7898 45724 7962 45728
rect 7898 45668 7902 45724
rect 7902 45668 7958 45724
rect 7958 45668 7962 45724
rect 7898 45664 7962 45668
rect 7978 45724 8042 45728
rect 7978 45668 7982 45724
rect 7982 45668 8038 45724
rect 8038 45668 8042 45724
rect 7978 45664 8042 45668
rect 8058 45724 8122 45728
rect 8058 45668 8062 45724
rect 8062 45668 8118 45724
rect 8118 45668 8122 45724
rect 8058 45664 8122 45668
rect 8138 45724 8202 45728
rect 8138 45668 8142 45724
rect 8142 45668 8198 45724
rect 8198 45668 8202 45724
rect 8138 45664 8202 45668
rect 14844 45724 14908 45728
rect 14844 45668 14848 45724
rect 14848 45668 14904 45724
rect 14904 45668 14908 45724
rect 14844 45664 14908 45668
rect 14924 45724 14988 45728
rect 14924 45668 14928 45724
rect 14928 45668 14984 45724
rect 14984 45668 14988 45724
rect 14924 45664 14988 45668
rect 15004 45724 15068 45728
rect 15004 45668 15008 45724
rect 15008 45668 15064 45724
rect 15064 45668 15068 45724
rect 15004 45664 15068 45668
rect 15084 45724 15148 45728
rect 15084 45668 15088 45724
rect 15088 45668 15144 45724
rect 15144 45668 15148 45724
rect 15084 45664 15148 45668
rect 21790 45724 21854 45728
rect 21790 45668 21794 45724
rect 21794 45668 21850 45724
rect 21850 45668 21854 45724
rect 21790 45664 21854 45668
rect 21870 45724 21934 45728
rect 21870 45668 21874 45724
rect 21874 45668 21930 45724
rect 21930 45668 21934 45724
rect 21870 45664 21934 45668
rect 21950 45724 22014 45728
rect 21950 45668 21954 45724
rect 21954 45668 22010 45724
rect 22010 45668 22014 45724
rect 21950 45664 22014 45668
rect 22030 45724 22094 45728
rect 22030 45668 22034 45724
rect 22034 45668 22090 45724
rect 22090 45668 22094 45724
rect 22030 45664 22094 45668
rect 28736 45724 28800 45728
rect 28736 45668 28740 45724
rect 28740 45668 28796 45724
rect 28796 45668 28800 45724
rect 28736 45664 28800 45668
rect 28816 45724 28880 45728
rect 28816 45668 28820 45724
rect 28820 45668 28876 45724
rect 28876 45668 28880 45724
rect 28816 45664 28880 45668
rect 28896 45724 28960 45728
rect 28896 45668 28900 45724
rect 28900 45668 28956 45724
rect 28956 45668 28960 45724
rect 28896 45664 28960 45668
rect 28976 45724 29040 45728
rect 28976 45668 28980 45724
rect 28980 45668 29036 45724
rect 29036 45668 29040 45724
rect 28976 45664 29040 45668
rect 4425 45180 4489 45184
rect 4425 45124 4429 45180
rect 4429 45124 4485 45180
rect 4485 45124 4489 45180
rect 4425 45120 4489 45124
rect 4505 45180 4569 45184
rect 4505 45124 4509 45180
rect 4509 45124 4565 45180
rect 4565 45124 4569 45180
rect 4505 45120 4569 45124
rect 4585 45180 4649 45184
rect 4585 45124 4589 45180
rect 4589 45124 4645 45180
rect 4645 45124 4649 45180
rect 4585 45120 4649 45124
rect 4665 45180 4729 45184
rect 4665 45124 4669 45180
rect 4669 45124 4725 45180
rect 4725 45124 4729 45180
rect 4665 45120 4729 45124
rect 11371 45180 11435 45184
rect 11371 45124 11375 45180
rect 11375 45124 11431 45180
rect 11431 45124 11435 45180
rect 11371 45120 11435 45124
rect 11451 45180 11515 45184
rect 11451 45124 11455 45180
rect 11455 45124 11511 45180
rect 11511 45124 11515 45180
rect 11451 45120 11515 45124
rect 11531 45180 11595 45184
rect 11531 45124 11535 45180
rect 11535 45124 11591 45180
rect 11591 45124 11595 45180
rect 11531 45120 11595 45124
rect 11611 45180 11675 45184
rect 11611 45124 11615 45180
rect 11615 45124 11671 45180
rect 11671 45124 11675 45180
rect 11611 45120 11675 45124
rect 18317 45180 18381 45184
rect 18317 45124 18321 45180
rect 18321 45124 18377 45180
rect 18377 45124 18381 45180
rect 18317 45120 18381 45124
rect 18397 45180 18461 45184
rect 18397 45124 18401 45180
rect 18401 45124 18457 45180
rect 18457 45124 18461 45180
rect 18397 45120 18461 45124
rect 18477 45180 18541 45184
rect 18477 45124 18481 45180
rect 18481 45124 18537 45180
rect 18537 45124 18541 45180
rect 18477 45120 18541 45124
rect 18557 45180 18621 45184
rect 18557 45124 18561 45180
rect 18561 45124 18617 45180
rect 18617 45124 18621 45180
rect 18557 45120 18621 45124
rect 25263 45180 25327 45184
rect 25263 45124 25267 45180
rect 25267 45124 25323 45180
rect 25323 45124 25327 45180
rect 25263 45120 25327 45124
rect 25343 45180 25407 45184
rect 25343 45124 25347 45180
rect 25347 45124 25403 45180
rect 25403 45124 25407 45180
rect 25343 45120 25407 45124
rect 25423 45180 25487 45184
rect 25423 45124 25427 45180
rect 25427 45124 25483 45180
rect 25483 45124 25487 45180
rect 25423 45120 25487 45124
rect 25503 45180 25567 45184
rect 25503 45124 25507 45180
rect 25507 45124 25563 45180
rect 25563 45124 25567 45180
rect 25503 45120 25567 45124
rect 7898 44636 7962 44640
rect 7898 44580 7902 44636
rect 7902 44580 7958 44636
rect 7958 44580 7962 44636
rect 7898 44576 7962 44580
rect 7978 44636 8042 44640
rect 7978 44580 7982 44636
rect 7982 44580 8038 44636
rect 8038 44580 8042 44636
rect 7978 44576 8042 44580
rect 8058 44636 8122 44640
rect 8058 44580 8062 44636
rect 8062 44580 8118 44636
rect 8118 44580 8122 44636
rect 8058 44576 8122 44580
rect 8138 44636 8202 44640
rect 8138 44580 8142 44636
rect 8142 44580 8198 44636
rect 8198 44580 8202 44636
rect 8138 44576 8202 44580
rect 14844 44636 14908 44640
rect 14844 44580 14848 44636
rect 14848 44580 14904 44636
rect 14904 44580 14908 44636
rect 14844 44576 14908 44580
rect 14924 44636 14988 44640
rect 14924 44580 14928 44636
rect 14928 44580 14984 44636
rect 14984 44580 14988 44636
rect 14924 44576 14988 44580
rect 15004 44636 15068 44640
rect 15004 44580 15008 44636
rect 15008 44580 15064 44636
rect 15064 44580 15068 44636
rect 15004 44576 15068 44580
rect 15084 44636 15148 44640
rect 15084 44580 15088 44636
rect 15088 44580 15144 44636
rect 15144 44580 15148 44636
rect 15084 44576 15148 44580
rect 21790 44636 21854 44640
rect 21790 44580 21794 44636
rect 21794 44580 21850 44636
rect 21850 44580 21854 44636
rect 21790 44576 21854 44580
rect 21870 44636 21934 44640
rect 21870 44580 21874 44636
rect 21874 44580 21930 44636
rect 21930 44580 21934 44636
rect 21870 44576 21934 44580
rect 21950 44636 22014 44640
rect 21950 44580 21954 44636
rect 21954 44580 22010 44636
rect 22010 44580 22014 44636
rect 21950 44576 22014 44580
rect 22030 44636 22094 44640
rect 22030 44580 22034 44636
rect 22034 44580 22090 44636
rect 22090 44580 22094 44636
rect 22030 44576 22094 44580
rect 28736 44636 28800 44640
rect 28736 44580 28740 44636
rect 28740 44580 28796 44636
rect 28796 44580 28800 44636
rect 28736 44576 28800 44580
rect 28816 44636 28880 44640
rect 28816 44580 28820 44636
rect 28820 44580 28876 44636
rect 28876 44580 28880 44636
rect 28816 44576 28880 44580
rect 28896 44636 28960 44640
rect 28896 44580 28900 44636
rect 28900 44580 28956 44636
rect 28956 44580 28960 44636
rect 28896 44576 28960 44580
rect 28976 44636 29040 44640
rect 28976 44580 28980 44636
rect 28980 44580 29036 44636
rect 29036 44580 29040 44636
rect 28976 44576 29040 44580
rect 4425 44092 4489 44096
rect 4425 44036 4429 44092
rect 4429 44036 4485 44092
rect 4485 44036 4489 44092
rect 4425 44032 4489 44036
rect 4505 44092 4569 44096
rect 4505 44036 4509 44092
rect 4509 44036 4565 44092
rect 4565 44036 4569 44092
rect 4505 44032 4569 44036
rect 4585 44092 4649 44096
rect 4585 44036 4589 44092
rect 4589 44036 4645 44092
rect 4645 44036 4649 44092
rect 4585 44032 4649 44036
rect 4665 44092 4729 44096
rect 4665 44036 4669 44092
rect 4669 44036 4725 44092
rect 4725 44036 4729 44092
rect 4665 44032 4729 44036
rect 11371 44092 11435 44096
rect 11371 44036 11375 44092
rect 11375 44036 11431 44092
rect 11431 44036 11435 44092
rect 11371 44032 11435 44036
rect 11451 44092 11515 44096
rect 11451 44036 11455 44092
rect 11455 44036 11511 44092
rect 11511 44036 11515 44092
rect 11451 44032 11515 44036
rect 11531 44092 11595 44096
rect 11531 44036 11535 44092
rect 11535 44036 11591 44092
rect 11591 44036 11595 44092
rect 11531 44032 11595 44036
rect 11611 44092 11675 44096
rect 11611 44036 11615 44092
rect 11615 44036 11671 44092
rect 11671 44036 11675 44092
rect 11611 44032 11675 44036
rect 18317 44092 18381 44096
rect 18317 44036 18321 44092
rect 18321 44036 18377 44092
rect 18377 44036 18381 44092
rect 18317 44032 18381 44036
rect 18397 44092 18461 44096
rect 18397 44036 18401 44092
rect 18401 44036 18457 44092
rect 18457 44036 18461 44092
rect 18397 44032 18461 44036
rect 18477 44092 18541 44096
rect 18477 44036 18481 44092
rect 18481 44036 18537 44092
rect 18537 44036 18541 44092
rect 18477 44032 18541 44036
rect 18557 44092 18621 44096
rect 18557 44036 18561 44092
rect 18561 44036 18617 44092
rect 18617 44036 18621 44092
rect 18557 44032 18621 44036
rect 25263 44092 25327 44096
rect 25263 44036 25267 44092
rect 25267 44036 25323 44092
rect 25323 44036 25327 44092
rect 25263 44032 25327 44036
rect 25343 44092 25407 44096
rect 25343 44036 25347 44092
rect 25347 44036 25403 44092
rect 25403 44036 25407 44092
rect 25343 44032 25407 44036
rect 25423 44092 25487 44096
rect 25423 44036 25427 44092
rect 25427 44036 25483 44092
rect 25483 44036 25487 44092
rect 25423 44032 25487 44036
rect 25503 44092 25567 44096
rect 25503 44036 25507 44092
rect 25507 44036 25563 44092
rect 25563 44036 25567 44092
rect 25503 44032 25567 44036
rect 7898 43548 7962 43552
rect 7898 43492 7902 43548
rect 7902 43492 7958 43548
rect 7958 43492 7962 43548
rect 7898 43488 7962 43492
rect 7978 43548 8042 43552
rect 7978 43492 7982 43548
rect 7982 43492 8038 43548
rect 8038 43492 8042 43548
rect 7978 43488 8042 43492
rect 8058 43548 8122 43552
rect 8058 43492 8062 43548
rect 8062 43492 8118 43548
rect 8118 43492 8122 43548
rect 8058 43488 8122 43492
rect 8138 43548 8202 43552
rect 8138 43492 8142 43548
rect 8142 43492 8198 43548
rect 8198 43492 8202 43548
rect 8138 43488 8202 43492
rect 14844 43548 14908 43552
rect 14844 43492 14848 43548
rect 14848 43492 14904 43548
rect 14904 43492 14908 43548
rect 14844 43488 14908 43492
rect 14924 43548 14988 43552
rect 14924 43492 14928 43548
rect 14928 43492 14984 43548
rect 14984 43492 14988 43548
rect 14924 43488 14988 43492
rect 15004 43548 15068 43552
rect 15004 43492 15008 43548
rect 15008 43492 15064 43548
rect 15064 43492 15068 43548
rect 15004 43488 15068 43492
rect 15084 43548 15148 43552
rect 15084 43492 15088 43548
rect 15088 43492 15144 43548
rect 15144 43492 15148 43548
rect 15084 43488 15148 43492
rect 21790 43548 21854 43552
rect 21790 43492 21794 43548
rect 21794 43492 21850 43548
rect 21850 43492 21854 43548
rect 21790 43488 21854 43492
rect 21870 43548 21934 43552
rect 21870 43492 21874 43548
rect 21874 43492 21930 43548
rect 21930 43492 21934 43548
rect 21870 43488 21934 43492
rect 21950 43548 22014 43552
rect 21950 43492 21954 43548
rect 21954 43492 22010 43548
rect 22010 43492 22014 43548
rect 21950 43488 22014 43492
rect 22030 43548 22094 43552
rect 22030 43492 22034 43548
rect 22034 43492 22090 43548
rect 22090 43492 22094 43548
rect 22030 43488 22094 43492
rect 28736 43548 28800 43552
rect 28736 43492 28740 43548
rect 28740 43492 28796 43548
rect 28796 43492 28800 43548
rect 28736 43488 28800 43492
rect 28816 43548 28880 43552
rect 28816 43492 28820 43548
rect 28820 43492 28876 43548
rect 28876 43492 28880 43548
rect 28816 43488 28880 43492
rect 28896 43548 28960 43552
rect 28896 43492 28900 43548
rect 28900 43492 28956 43548
rect 28956 43492 28960 43548
rect 28896 43488 28960 43492
rect 28976 43548 29040 43552
rect 28976 43492 28980 43548
rect 28980 43492 29036 43548
rect 29036 43492 29040 43548
rect 28976 43488 29040 43492
rect 4425 43004 4489 43008
rect 4425 42948 4429 43004
rect 4429 42948 4485 43004
rect 4485 42948 4489 43004
rect 4425 42944 4489 42948
rect 4505 43004 4569 43008
rect 4505 42948 4509 43004
rect 4509 42948 4565 43004
rect 4565 42948 4569 43004
rect 4505 42944 4569 42948
rect 4585 43004 4649 43008
rect 4585 42948 4589 43004
rect 4589 42948 4645 43004
rect 4645 42948 4649 43004
rect 4585 42944 4649 42948
rect 4665 43004 4729 43008
rect 4665 42948 4669 43004
rect 4669 42948 4725 43004
rect 4725 42948 4729 43004
rect 4665 42944 4729 42948
rect 11371 43004 11435 43008
rect 11371 42948 11375 43004
rect 11375 42948 11431 43004
rect 11431 42948 11435 43004
rect 11371 42944 11435 42948
rect 11451 43004 11515 43008
rect 11451 42948 11455 43004
rect 11455 42948 11511 43004
rect 11511 42948 11515 43004
rect 11451 42944 11515 42948
rect 11531 43004 11595 43008
rect 11531 42948 11535 43004
rect 11535 42948 11591 43004
rect 11591 42948 11595 43004
rect 11531 42944 11595 42948
rect 11611 43004 11675 43008
rect 11611 42948 11615 43004
rect 11615 42948 11671 43004
rect 11671 42948 11675 43004
rect 11611 42944 11675 42948
rect 18317 43004 18381 43008
rect 18317 42948 18321 43004
rect 18321 42948 18377 43004
rect 18377 42948 18381 43004
rect 18317 42944 18381 42948
rect 18397 43004 18461 43008
rect 18397 42948 18401 43004
rect 18401 42948 18457 43004
rect 18457 42948 18461 43004
rect 18397 42944 18461 42948
rect 18477 43004 18541 43008
rect 18477 42948 18481 43004
rect 18481 42948 18537 43004
rect 18537 42948 18541 43004
rect 18477 42944 18541 42948
rect 18557 43004 18621 43008
rect 18557 42948 18561 43004
rect 18561 42948 18617 43004
rect 18617 42948 18621 43004
rect 18557 42944 18621 42948
rect 25263 43004 25327 43008
rect 25263 42948 25267 43004
rect 25267 42948 25323 43004
rect 25323 42948 25327 43004
rect 25263 42944 25327 42948
rect 25343 43004 25407 43008
rect 25343 42948 25347 43004
rect 25347 42948 25403 43004
rect 25403 42948 25407 43004
rect 25343 42944 25407 42948
rect 25423 43004 25487 43008
rect 25423 42948 25427 43004
rect 25427 42948 25483 43004
rect 25483 42948 25487 43004
rect 25423 42944 25487 42948
rect 25503 43004 25567 43008
rect 25503 42948 25507 43004
rect 25507 42948 25563 43004
rect 25563 42948 25567 43004
rect 25503 42944 25567 42948
rect 19564 42876 19628 42940
rect 7898 42460 7962 42464
rect 7898 42404 7902 42460
rect 7902 42404 7958 42460
rect 7958 42404 7962 42460
rect 7898 42400 7962 42404
rect 7978 42460 8042 42464
rect 7978 42404 7982 42460
rect 7982 42404 8038 42460
rect 8038 42404 8042 42460
rect 7978 42400 8042 42404
rect 8058 42460 8122 42464
rect 8058 42404 8062 42460
rect 8062 42404 8118 42460
rect 8118 42404 8122 42460
rect 8058 42400 8122 42404
rect 8138 42460 8202 42464
rect 8138 42404 8142 42460
rect 8142 42404 8198 42460
rect 8198 42404 8202 42460
rect 8138 42400 8202 42404
rect 14844 42460 14908 42464
rect 14844 42404 14848 42460
rect 14848 42404 14904 42460
rect 14904 42404 14908 42460
rect 14844 42400 14908 42404
rect 14924 42460 14988 42464
rect 14924 42404 14928 42460
rect 14928 42404 14984 42460
rect 14984 42404 14988 42460
rect 14924 42400 14988 42404
rect 15004 42460 15068 42464
rect 15004 42404 15008 42460
rect 15008 42404 15064 42460
rect 15064 42404 15068 42460
rect 15004 42400 15068 42404
rect 15084 42460 15148 42464
rect 15084 42404 15088 42460
rect 15088 42404 15144 42460
rect 15144 42404 15148 42460
rect 15084 42400 15148 42404
rect 21790 42460 21854 42464
rect 21790 42404 21794 42460
rect 21794 42404 21850 42460
rect 21850 42404 21854 42460
rect 21790 42400 21854 42404
rect 21870 42460 21934 42464
rect 21870 42404 21874 42460
rect 21874 42404 21930 42460
rect 21930 42404 21934 42460
rect 21870 42400 21934 42404
rect 21950 42460 22014 42464
rect 21950 42404 21954 42460
rect 21954 42404 22010 42460
rect 22010 42404 22014 42460
rect 21950 42400 22014 42404
rect 22030 42460 22094 42464
rect 22030 42404 22034 42460
rect 22034 42404 22090 42460
rect 22090 42404 22094 42460
rect 22030 42400 22094 42404
rect 28736 42460 28800 42464
rect 28736 42404 28740 42460
rect 28740 42404 28796 42460
rect 28796 42404 28800 42460
rect 28736 42400 28800 42404
rect 28816 42460 28880 42464
rect 28816 42404 28820 42460
rect 28820 42404 28876 42460
rect 28876 42404 28880 42460
rect 28816 42400 28880 42404
rect 28896 42460 28960 42464
rect 28896 42404 28900 42460
rect 28900 42404 28956 42460
rect 28956 42404 28960 42460
rect 28896 42400 28960 42404
rect 28976 42460 29040 42464
rect 28976 42404 28980 42460
rect 28980 42404 29036 42460
rect 29036 42404 29040 42460
rect 28976 42400 29040 42404
rect 4425 41916 4489 41920
rect 4425 41860 4429 41916
rect 4429 41860 4485 41916
rect 4485 41860 4489 41916
rect 4425 41856 4489 41860
rect 4505 41916 4569 41920
rect 4505 41860 4509 41916
rect 4509 41860 4565 41916
rect 4565 41860 4569 41916
rect 4505 41856 4569 41860
rect 4585 41916 4649 41920
rect 4585 41860 4589 41916
rect 4589 41860 4645 41916
rect 4645 41860 4649 41916
rect 4585 41856 4649 41860
rect 4665 41916 4729 41920
rect 4665 41860 4669 41916
rect 4669 41860 4725 41916
rect 4725 41860 4729 41916
rect 4665 41856 4729 41860
rect 11371 41916 11435 41920
rect 11371 41860 11375 41916
rect 11375 41860 11431 41916
rect 11431 41860 11435 41916
rect 11371 41856 11435 41860
rect 11451 41916 11515 41920
rect 11451 41860 11455 41916
rect 11455 41860 11511 41916
rect 11511 41860 11515 41916
rect 11451 41856 11515 41860
rect 11531 41916 11595 41920
rect 11531 41860 11535 41916
rect 11535 41860 11591 41916
rect 11591 41860 11595 41916
rect 11531 41856 11595 41860
rect 11611 41916 11675 41920
rect 11611 41860 11615 41916
rect 11615 41860 11671 41916
rect 11671 41860 11675 41916
rect 11611 41856 11675 41860
rect 18317 41916 18381 41920
rect 18317 41860 18321 41916
rect 18321 41860 18377 41916
rect 18377 41860 18381 41916
rect 18317 41856 18381 41860
rect 18397 41916 18461 41920
rect 18397 41860 18401 41916
rect 18401 41860 18457 41916
rect 18457 41860 18461 41916
rect 18397 41856 18461 41860
rect 18477 41916 18541 41920
rect 18477 41860 18481 41916
rect 18481 41860 18537 41916
rect 18537 41860 18541 41916
rect 18477 41856 18541 41860
rect 18557 41916 18621 41920
rect 18557 41860 18561 41916
rect 18561 41860 18617 41916
rect 18617 41860 18621 41916
rect 18557 41856 18621 41860
rect 25263 41916 25327 41920
rect 25263 41860 25267 41916
rect 25267 41860 25323 41916
rect 25323 41860 25327 41916
rect 25263 41856 25327 41860
rect 25343 41916 25407 41920
rect 25343 41860 25347 41916
rect 25347 41860 25403 41916
rect 25403 41860 25407 41916
rect 25343 41856 25407 41860
rect 25423 41916 25487 41920
rect 25423 41860 25427 41916
rect 25427 41860 25483 41916
rect 25483 41860 25487 41916
rect 25423 41856 25487 41860
rect 25503 41916 25567 41920
rect 25503 41860 25507 41916
rect 25507 41860 25563 41916
rect 25563 41860 25567 41916
rect 25503 41856 25567 41860
rect 7898 41372 7962 41376
rect 7898 41316 7902 41372
rect 7902 41316 7958 41372
rect 7958 41316 7962 41372
rect 7898 41312 7962 41316
rect 7978 41372 8042 41376
rect 7978 41316 7982 41372
rect 7982 41316 8038 41372
rect 8038 41316 8042 41372
rect 7978 41312 8042 41316
rect 8058 41372 8122 41376
rect 8058 41316 8062 41372
rect 8062 41316 8118 41372
rect 8118 41316 8122 41372
rect 8058 41312 8122 41316
rect 8138 41372 8202 41376
rect 8138 41316 8142 41372
rect 8142 41316 8198 41372
rect 8198 41316 8202 41372
rect 8138 41312 8202 41316
rect 14844 41372 14908 41376
rect 14844 41316 14848 41372
rect 14848 41316 14904 41372
rect 14904 41316 14908 41372
rect 14844 41312 14908 41316
rect 14924 41372 14988 41376
rect 14924 41316 14928 41372
rect 14928 41316 14984 41372
rect 14984 41316 14988 41372
rect 14924 41312 14988 41316
rect 15004 41372 15068 41376
rect 15004 41316 15008 41372
rect 15008 41316 15064 41372
rect 15064 41316 15068 41372
rect 15004 41312 15068 41316
rect 15084 41372 15148 41376
rect 15084 41316 15088 41372
rect 15088 41316 15144 41372
rect 15144 41316 15148 41372
rect 15084 41312 15148 41316
rect 21790 41372 21854 41376
rect 21790 41316 21794 41372
rect 21794 41316 21850 41372
rect 21850 41316 21854 41372
rect 21790 41312 21854 41316
rect 21870 41372 21934 41376
rect 21870 41316 21874 41372
rect 21874 41316 21930 41372
rect 21930 41316 21934 41372
rect 21870 41312 21934 41316
rect 21950 41372 22014 41376
rect 21950 41316 21954 41372
rect 21954 41316 22010 41372
rect 22010 41316 22014 41372
rect 21950 41312 22014 41316
rect 22030 41372 22094 41376
rect 22030 41316 22034 41372
rect 22034 41316 22090 41372
rect 22090 41316 22094 41372
rect 22030 41312 22094 41316
rect 28736 41372 28800 41376
rect 28736 41316 28740 41372
rect 28740 41316 28796 41372
rect 28796 41316 28800 41372
rect 28736 41312 28800 41316
rect 28816 41372 28880 41376
rect 28816 41316 28820 41372
rect 28820 41316 28876 41372
rect 28876 41316 28880 41372
rect 28816 41312 28880 41316
rect 28896 41372 28960 41376
rect 28896 41316 28900 41372
rect 28900 41316 28956 41372
rect 28956 41316 28960 41372
rect 28896 41312 28960 41316
rect 28976 41372 29040 41376
rect 28976 41316 28980 41372
rect 28980 41316 29036 41372
rect 29036 41316 29040 41372
rect 28976 41312 29040 41316
rect 4425 40828 4489 40832
rect 4425 40772 4429 40828
rect 4429 40772 4485 40828
rect 4485 40772 4489 40828
rect 4425 40768 4489 40772
rect 4505 40828 4569 40832
rect 4505 40772 4509 40828
rect 4509 40772 4565 40828
rect 4565 40772 4569 40828
rect 4505 40768 4569 40772
rect 4585 40828 4649 40832
rect 4585 40772 4589 40828
rect 4589 40772 4645 40828
rect 4645 40772 4649 40828
rect 4585 40768 4649 40772
rect 4665 40828 4729 40832
rect 4665 40772 4669 40828
rect 4669 40772 4725 40828
rect 4725 40772 4729 40828
rect 4665 40768 4729 40772
rect 11371 40828 11435 40832
rect 11371 40772 11375 40828
rect 11375 40772 11431 40828
rect 11431 40772 11435 40828
rect 11371 40768 11435 40772
rect 11451 40828 11515 40832
rect 11451 40772 11455 40828
rect 11455 40772 11511 40828
rect 11511 40772 11515 40828
rect 11451 40768 11515 40772
rect 11531 40828 11595 40832
rect 11531 40772 11535 40828
rect 11535 40772 11591 40828
rect 11591 40772 11595 40828
rect 11531 40768 11595 40772
rect 11611 40828 11675 40832
rect 11611 40772 11615 40828
rect 11615 40772 11671 40828
rect 11671 40772 11675 40828
rect 11611 40768 11675 40772
rect 18317 40828 18381 40832
rect 18317 40772 18321 40828
rect 18321 40772 18377 40828
rect 18377 40772 18381 40828
rect 18317 40768 18381 40772
rect 18397 40828 18461 40832
rect 18397 40772 18401 40828
rect 18401 40772 18457 40828
rect 18457 40772 18461 40828
rect 18397 40768 18461 40772
rect 18477 40828 18541 40832
rect 18477 40772 18481 40828
rect 18481 40772 18537 40828
rect 18537 40772 18541 40828
rect 18477 40768 18541 40772
rect 18557 40828 18621 40832
rect 18557 40772 18561 40828
rect 18561 40772 18617 40828
rect 18617 40772 18621 40828
rect 18557 40768 18621 40772
rect 25263 40828 25327 40832
rect 25263 40772 25267 40828
rect 25267 40772 25323 40828
rect 25323 40772 25327 40828
rect 25263 40768 25327 40772
rect 25343 40828 25407 40832
rect 25343 40772 25347 40828
rect 25347 40772 25403 40828
rect 25403 40772 25407 40828
rect 25343 40768 25407 40772
rect 25423 40828 25487 40832
rect 25423 40772 25427 40828
rect 25427 40772 25483 40828
rect 25483 40772 25487 40828
rect 25423 40768 25487 40772
rect 25503 40828 25567 40832
rect 25503 40772 25507 40828
rect 25507 40772 25563 40828
rect 25563 40772 25567 40828
rect 25503 40768 25567 40772
rect 7898 40284 7962 40288
rect 7898 40228 7902 40284
rect 7902 40228 7958 40284
rect 7958 40228 7962 40284
rect 7898 40224 7962 40228
rect 7978 40284 8042 40288
rect 7978 40228 7982 40284
rect 7982 40228 8038 40284
rect 8038 40228 8042 40284
rect 7978 40224 8042 40228
rect 8058 40284 8122 40288
rect 8058 40228 8062 40284
rect 8062 40228 8118 40284
rect 8118 40228 8122 40284
rect 8058 40224 8122 40228
rect 8138 40284 8202 40288
rect 8138 40228 8142 40284
rect 8142 40228 8198 40284
rect 8198 40228 8202 40284
rect 8138 40224 8202 40228
rect 14844 40284 14908 40288
rect 14844 40228 14848 40284
rect 14848 40228 14904 40284
rect 14904 40228 14908 40284
rect 14844 40224 14908 40228
rect 14924 40284 14988 40288
rect 14924 40228 14928 40284
rect 14928 40228 14984 40284
rect 14984 40228 14988 40284
rect 14924 40224 14988 40228
rect 15004 40284 15068 40288
rect 15004 40228 15008 40284
rect 15008 40228 15064 40284
rect 15064 40228 15068 40284
rect 15004 40224 15068 40228
rect 15084 40284 15148 40288
rect 15084 40228 15088 40284
rect 15088 40228 15144 40284
rect 15144 40228 15148 40284
rect 15084 40224 15148 40228
rect 21790 40284 21854 40288
rect 21790 40228 21794 40284
rect 21794 40228 21850 40284
rect 21850 40228 21854 40284
rect 21790 40224 21854 40228
rect 21870 40284 21934 40288
rect 21870 40228 21874 40284
rect 21874 40228 21930 40284
rect 21930 40228 21934 40284
rect 21870 40224 21934 40228
rect 21950 40284 22014 40288
rect 21950 40228 21954 40284
rect 21954 40228 22010 40284
rect 22010 40228 22014 40284
rect 21950 40224 22014 40228
rect 22030 40284 22094 40288
rect 22030 40228 22034 40284
rect 22034 40228 22090 40284
rect 22090 40228 22094 40284
rect 22030 40224 22094 40228
rect 28736 40284 28800 40288
rect 28736 40228 28740 40284
rect 28740 40228 28796 40284
rect 28796 40228 28800 40284
rect 28736 40224 28800 40228
rect 28816 40284 28880 40288
rect 28816 40228 28820 40284
rect 28820 40228 28876 40284
rect 28876 40228 28880 40284
rect 28816 40224 28880 40228
rect 28896 40284 28960 40288
rect 28896 40228 28900 40284
rect 28900 40228 28956 40284
rect 28956 40228 28960 40284
rect 28896 40224 28960 40228
rect 28976 40284 29040 40288
rect 28976 40228 28980 40284
rect 28980 40228 29036 40284
rect 29036 40228 29040 40284
rect 28976 40224 29040 40228
rect 4425 39740 4489 39744
rect 4425 39684 4429 39740
rect 4429 39684 4485 39740
rect 4485 39684 4489 39740
rect 4425 39680 4489 39684
rect 4505 39740 4569 39744
rect 4505 39684 4509 39740
rect 4509 39684 4565 39740
rect 4565 39684 4569 39740
rect 4505 39680 4569 39684
rect 4585 39740 4649 39744
rect 4585 39684 4589 39740
rect 4589 39684 4645 39740
rect 4645 39684 4649 39740
rect 4585 39680 4649 39684
rect 4665 39740 4729 39744
rect 4665 39684 4669 39740
rect 4669 39684 4725 39740
rect 4725 39684 4729 39740
rect 4665 39680 4729 39684
rect 11371 39740 11435 39744
rect 11371 39684 11375 39740
rect 11375 39684 11431 39740
rect 11431 39684 11435 39740
rect 11371 39680 11435 39684
rect 11451 39740 11515 39744
rect 11451 39684 11455 39740
rect 11455 39684 11511 39740
rect 11511 39684 11515 39740
rect 11451 39680 11515 39684
rect 11531 39740 11595 39744
rect 11531 39684 11535 39740
rect 11535 39684 11591 39740
rect 11591 39684 11595 39740
rect 11531 39680 11595 39684
rect 11611 39740 11675 39744
rect 11611 39684 11615 39740
rect 11615 39684 11671 39740
rect 11671 39684 11675 39740
rect 11611 39680 11675 39684
rect 18317 39740 18381 39744
rect 18317 39684 18321 39740
rect 18321 39684 18377 39740
rect 18377 39684 18381 39740
rect 18317 39680 18381 39684
rect 18397 39740 18461 39744
rect 18397 39684 18401 39740
rect 18401 39684 18457 39740
rect 18457 39684 18461 39740
rect 18397 39680 18461 39684
rect 18477 39740 18541 39744
rect 18477 39684 18481 39740
rect 18481 39684 18537 39740
rect 18537 39684 18541 39740
rect 18477 39680 18541 39684
rect 18557 39740 18621 39744
rect 18557 39684 18561 39740
rect 18561 39684 18617 39740
rect 18617 39684 18621 39740
rect 18557 39680 18621 39684
rect 25263 39740 25327 39744
rect 25263 39684 25267 39740
rect 25267 39684 25323 39740
rect 25323 39684 25327 39740
rect 25263 39680 25327 39684
rect 25343 39740 25407 39744
rect 25343 39684 25347 39740
rect 25347 39684 25403 39740
rect 25403 39684 25407 39740
rect 25343 39680 25407 39684
rect 25423 39740 25487 39744
rect 25423 39684 25427 39740
rect 25427 39684 25483 39740
rect 25483 39684 25487 39740
rect 25423 39680 25487 39684
rect 25503 39740 25567 39744
rect 25503 39684 25507 39740
rect 25507 39684 25563 39740
rect 25563 39684 25567 39740
rect 25503 39680 25567 39684
rect 7898 39196 7962 39200
rect 7898 39140 7902 39196
rect 7902 39140 7958 39196
rect 7958 39140 7962 39196
rect 7898 39136 7962 39140
rect 7978 39196 8042 39200
rect 7978 39140 7982 39196
rect 7982 39140 8038 39196
rect 8038 39140 8042 39196
rect 7978 39136 8042 39140
rect 8058 39196 8122 39200
rect 8058 39140 8062 39196
rect 8062 39140 8118 39196
rect 8118 39140 8122 39196
rect 8058 39136 8122 39140
rect 8138 39196 8202 39200
rect 8138 39140 8142 39196
rect 8142 39140 8198 39196
rect 8198 39140 8202 39196
rect 8138 39136 8202 39140
rect 14844 39196 14908 39200
rect 14844 39140 14848 39196
rect 14848 39140 14904 39196
rect 14904 39140 14908 39196
rect 14844 39136 14908 39140
rect 14924 39196 14988 39200
rect 14924 39140 14928 39196
rect 14928 39140 14984 39196
rect 14984 39140 14988 39196
rect 14924 39136 14988 39140
rect 15004 39196 15068 39200
rect 15004 39140 15008 39196
rect 15008 39140 15064 39196
rect 15064 39140 15068 39196
rect 15004 39136 15068 39140
rect 15084 39196 15148 39200
rect 15084 39140 15088 39196
rect 15088 39140 15144 39196
rect 15144 39140 15148 39196
rect 15084 39136 15148 39140
rect 21790 39196 21854 39200
rect 21790 39140 21794 39196
rect 21794 39140 21850 39196
rect 21850 39140 21854 39196
rect 21790 39136 21854 39140
rect 21870 39196 21934 39200
rect 21870 39140 21874 39196
rect 21874 39140 21930 39196
rect 21930 39140 21934 39196
rect 21870 39136 21934 39140
rect 21950 39196 22014 39200
rect 21950 39140 21954 39196
rect 21954 39140 22010 39196
rect 22010 39140 22014 39196
rect 21950 39136 22014 39140
rect 22030 39196 22094 39200
rect 22030 39140 22034 39196
rect 22034 39140 22090 39196
rect 22090 39140 22094 39196
rect 22030 39136 22094 39140
rect 28736 39196 28800 39200
rect 28736 39140 28740 39196
rect 28740 39140 28796 39196
rect 28796 39140 28800 39196
rect 28736 39136 28800 39140
rect 28816 39196 28880 39200
rect 28816 39140 28820 39196
rect 28820 39140 28876 39196
rect 28876 39140 28880 39196
rect 28816 39136 28880 39140
rect 28896 39196 28960 39200
rect 28896 39140 28900 39196
rect 28900 39140 28956 39196
rect 28956 39140 28960 39196
rect 28896 39136 28960 39140
rect 28976 39196 29040 39200
rect 28976 39140 28980 39196
rect 28980 39140 29036 39196
rect 29036 39140 29040 39196
rect 28976 39136 29040 39140
rect 4425 38652 4489 38656
rect 4425 38596 4429 38652
rect 4429 38596 4485 38652
rect 4485 38596 4489 38652
rect 4425 38592 4489 38596
rect 4505 38652 4569 38656
rect 4505 38596 4509 38652
rect 4509 38596 4565 38652
rect 4565 38596 4569 38652
rect 4505 38592 4569 38596
rect 4585 38652 4649 38656
rect 4585 38596 4589 38652
rect 4589 38596 4645 38652
rect 4645 38596 4649 38652
rect 4585 38592 4649 38596
rect 4665 38652 4729 38656
rect 4665 38596 4669 38652
rect 4669 38596 4725 38652
rect 4725 38596 4729 38652
rect 4665 38592 4729 38596
rect 11371 38652 11435 38656
rect 11371 38596 11375 38652
rect 11375 38596 11431 38652
rect 11431 38596 11435 38652
rect 11371 38592 11435 38596
rect 11451 38652 11515 38656
rect 11451 38596 11455 38652
rect 11455 38596 11511 38652
rect 11511 38596 11515 38652
rect 11451 38592 11515 38596
rect 11531 38652 11595 38656
rect 11531 38596 11535 38652
rect 11535 38596 11591 38652
rect 11591 38596 11595 38652
rect 11531 38592 11595 38596
rect 11611 38652 11675 38656
rect 11611 38596 11615 38652
rect 11615 38596 11671 38652
rect 11671 38596 11675 38652
rect 11611 38592 11675 38596
rect 18317 38652 18381 38656
rect 18317 38596 18321 38652
rect 18321 38596 18377 38652
rect 18377 38596 18381 38652
rect 18317 38592 18381 38596
rect 18397 38652 18461 38656
rect 18397 38596 18401 38652
rect 18401 38596 18457 38652
rect 18457 38596 18461 38652
rect 18397 38592 18461 38596
rect 18477 38652 18541 38656
rect 18477 38596 18481 38652
rect 18481 38596 18537 38652
rect 18537 38596 18541 38652
rect 18477 38592 18541 38596
rect 18557 38652 18621 38656
rect 18557 38596 18561 38652
rect 18561 38596 18617 38652
rect 18617 38596 18621 38652
rect 18557 38592 18621 38596
rect 25263 38652 25327 38656
rect 25263 38596 25267 38652
rect 25267 38596 25323 38652
rect 25323 38596 25327 38652
rect 25263 38592 25327 38596
rect 25343 38652 25407 38656
rect 25343 38596 25347 38652
rect 25347 38596 25403 38652
rect 25403 38596 25407 38652
rect 25343 38592 25407 38596
rect 25423 38652 25487 38656
rect 25423 38596 25427 38652
rect 25427 38596 25483 38652
rect 25483 38596 25487 38652
rect 25423 38592 25487 38596
rect 25503 38652 25567 38656
rect 25503 38596 25507 38652
rect 25507 38596 25563 38652
rect 25563 38596 25567 38652
rect 25503 38592 25567 38596
rect 7898 38108 7962 38112
rect 7898 38052 7902 38108
rect 7902 38052 7958 38108
rect 7958 38052 7962 38108
rect 7898 38048 7962 38052
rect 7978 38108 8042 38112
rect 7978 38052 7982 38108
rect 7982 38052 8038 38108
rect 8038 38052 8042 38108
rect 7978 38048 8042 38052
rect 8058 38108 8122 38112
rect 8058 38052 8062 38108
rect 8062 38052 8118 38108
rect 8118 38052 8122 38108
rect 8058 38048 8122 38052
rect 8138 38108 8202 38112
rect 8138 38052 8142 38108
rect 8142 38052 8198 38108
rect 8198 38052 8202 38108
rect 8138 38048 8202 38052
rect 14844 38108 14908 38112
rect 14844 38052 14848 38108
rect 14848 38052 14904 38108
rect 14904 38052 14908 38108
rect 14844 38048 14908 38052
rect 14924 38108 14988 38112
rect 14924 38052 14928 38108
rect 14928 38052 14984 38108
rect 14984 38052 14988 38108
rect 14924 38048 14988 38052
rect 15004 38108 15068 38112
rect 15004 38052 15008 38108
rect 15008 38052 15064 38108
rect 15064 38052 15068 38108
rect 15004 38048 15068 38052
rect 15084 38108 15148 38112
rect 15084 38052 15088 38108
rect 15088 38052 15144 38108
rect 15144 38052 15148 38108
rect 15084 38048 15148 38052
rect 21790 38108 21854 38112
rect 21790 38052 21794 38108
rect 21794 38052 21850 38108
rect 21850 38052 21854 38108
rect 21790 38048 21854 38052
rect 21870 38108 21934 38112
rect 21870 38052 21874 38108
rect 21874 38052 21930 38108
rect 21930 38052 21934 38108
rect 21870 38048 21934 38052
rect 21950 38108 22014 38112
rect 21950 38052 21954 38108
rect 21954 38052 22010 38108
rect 22010 38052 22014 38108
rect 21950 38048 22014 38052
rect 22030 38108 22094 38112
rect 22030 38052 22034 38108
rect 22034 38052 22090 38108
rect 22090 38052 22094 38108
rect 22030 38048 22094 38052
rect 28736 38108 28800 38112
rect 28736 38052 28740 38108
rect 28740 38052 28796 38108
rect 28796 38052 28800 38108
rect 28736 38048 28800 38052
rect 28816 38108 28880 38112
rect 28816 38052 28820 38108
rect 28820 38052 28876 38108
rect 28876 38052 28880 38108
rect 28816 38048 28880 38052
rect 28896 38108 28960 38112
rect 28896 38052 28900 38108
rect 28900 38052 28956 38108
rect 28956 38052 28960 38108
rect 28896 38048 28960 38052
rect 28976 38108 29040 38112
rect 28976 38052 28980 38108
rect 28980 38052 29036 38108
rect 29036 38052 29040 38108
rect 28976 38048 29040 38052
rect 4425 37564 4489 37568
rect 4425 37508 4429 37564
rect 4429 37508 4485 37564
rect 4485 37508 4489 37564
rect 4425 37504 4489 37508
rect 4505 37564 4569 37568
rect 4505 37508 4509 37564
rect 4509 37508 4565 37564
rect 4565 37508 4569 37564
rect 4505 37504 4569 37508
rect 4585 37564 4649 37568
rect 4585 37508 4589 37564
rect 4589 37508 4645 37564
rect 4645 37508 4649 37564
rect 4585 37504 4649 37508
rect 4665 37564 4729 37568
rect 4665 37508 4669 37564
rect 4669 37508 4725 37564
rect 4725 37508 4729 37564
rect 4665 37504 4729 37508
rect 11371 37564 11435 37568
rect 11371 37508 11375 37564
rect 11375 37508 11431 37564
rect 11431 37508 11435 37564
rect 11371 37504 11435 37508
rect 11451 37564 11515 37568
rect 11451 37508 11455 37564
rect 11455 37508 11511 37564
rect 11511 37508 11515 37564
rect 11451 37504 11515 37508
rect 11531 37564 11595 37568
rect 11531 37508 11535 37564
rect 11535 37508 11591 37564
rect 11591 37508 11595 37564
rect 11531 37504 11595 37508
rect 11611 37564 11675 37568
rect 11611 37508 11615 37564
rect 11615 37508 11671 37564
rect 11671 37508 11675 37564
rect 11611 37504 11675 37508
rect 18317 37564 18381 37568
rect 18317 37508 18321 37564
rect 18321 37508 18377 37564
rect 18377 37508 18381 37564
rect 18317 37504 18381 37508
rect 18397 37564 18461 37568
rect 18397 37508 18401 37564
rect 18401 37508 18457 37564
rect 18457 37508 18461 37564
rect 18397 37504 18461 37508
rect 18477 37564 18541 37568
rect 18477 37508 18481 37564
rect 18481 37508 18537 37564
rect 18537 37508 18541 37564
rect 18477 37504 18541 37508
rect 18557 37564 18621 37568
rect 18557 37508 18561 37564
rect 18561 37508 18617 37564
rect 18617 37508 18621 37564
rect 18557 37504 18621 37508
rect 25263 37564 25327 37568
rect 25263 37508 25267 37564
rect 25267 37508 25323 37564
rect 25323 37508 25327 37564
rect 25263 37504 25327 37508
rect 25343 37564 25407 37568
rect 25343 37508 25347 37564
rect 25347 37508 25403 37564
rect 25403 37508 25407 37564
rect 25343 37504 25407 37508
rect 25423 37564 25487 37568
rect 25423 37508 25427 37564
rect 25427 37508 25483 37564
rect 25483 37508 25487 37564
rect 25423 37504 25487 37508
rect 25503 37564 25567 37568
rect 25503 37508 25507 37564
rect 25507 37508 25563 37564
rect 25563 37508 25567 37564
rect 25503 37504 25567 37508
rect 7898 37020 7962 37024
rect 7898 36964 7902 37020
rect 7902 36964 7958 37020
rect 7958 36964 7962 37020
rect 7898 36960 7962 36964
rect 7978 37020 8042 37024
rect 7978 36964 7982 37020
rect 7982 36964 8038 37020
rect 8038 36964 8042 37020
rect 7978 36960 8042 36964
rect 8058 37020 8122 37024
rect 8058 36964 8062 37020
rect 8062 36964 8118 37020
rect 8118 36964 8122 37020
rect 8058 36960 8122 36964
rect 8138 37020 8202 37024
rect 8138 36964 8142 37020
rect 8142 36964 8198 37020
rect 8198 36964 8202 37020
rect 8138 36960 8202 36964
rect 14844 37020 14908 37024
rect 14844 36964 14848 37020
rect 14848 36964 14904 37020
rect 14904 36964 14908 37020
rect 14844 36960 14908 36964
rect 14924 37020 14988 37024
rect 14924 36964 14928 37020
rect 14928 36964 14984 37020
rect 14984 36964 14988 37020
rect 14924 36960 14988 36964
rect 15004 37020 15068 37024
rect 15004 36964 15008 37020
rect 15008 36964 15064 37020
rect 15064 36964 15068 37020
rect 15004 36960 15068 36964
rect 15084 37020 15148 37024
rect 15084 36964 15088 37020
rect 15088 36964 15144 37020
rect 15144 36964 15148 37020
rect 15084 36960 15148 36964
rect 21790 37020 21854 37024
rect 21790 36964 21794 37020
rect 21794 36964 21850 37020
rect 21850 36964 21854 37020
rect 21790 36960 21854 36964
rect 21870 37020 21934 37024
rect 21870 36964 21874 37020
rect 21874 36964 21930 37020
rect 21930 36964 21934 37020
rect 21870 36960 21934 36964
rect 21950 37020 22014 37024
rect 21950 36964 21954 37020
rect 21954 36964 22010 37020
rect 22010 36964 22014 37020
rect 21950 36960 22014 36964
rect 22030 37020 22094 37024
rect 22030 36964 22034 37020
rect 22034 36964 22090 37020
rect 22090 36964 22094 37020
rect 22030 36960 22094 36964
rect 28736 37020 28800 37024
rect 28736 36964 28740 37020
rect 28740 36964 28796 37020
rect 28796 36964 28800 37020
rect 28736 36960 28800 36964
rect 28816 37020 28880 37024
rect 28816 36964 28820 37020
rect 28820 36964 28876 37020
rect 28876 36964 28880 37020
rect 28816 36960 28880 36964
rect 28896 37020 28960 37024
rect 28896 36964 28900 37020
rect 28900 36964 28956 37020
rect 28956 36964 28960 37020
rect 28896 36960 28960 36964
rect 28976 37020 29040 37024
rect 28976 36964 28980 37020
rect 28980 36964 29036 37020
rect 29036 36964 29040 37020
rect 28976 36960 29040 36964
rect 4425 36476 4489 36480
rect 4425 36420 4429 36476
rect 4429 36420 4485 36476
rect 4485 36420 4489 36476
rect 4425 36416 4489 36420
rect 4505 36476 4569 36480
rect 4505 36420 4509 36476
rect 4509 36420 4565 36476
rect 4565 36420 4569 36476
rect 4505 36416 4569 36420
rect 4585 36476 4649 36480
rect 4585 36420 4589 36476
rect 4589 36420 4645 36476
rect 4645 36420 4649 36476
rect 4585 36416 4649 36420
rect 4665 36476 4729 36480
rect 4665 36420 4669 36476
rect 4669 36420 4725 36476
rect 4725 36420 4729 36476
rect 4665 36416 4729 36420
rect 11371 36476 11435 36480
rect 11371 36420 11375 36476
rect 11375 36420 11431 36476
rect 11431 36420 11435 36476
rect 11371 36416 11435 36420
rect 11451 36476 11515 36480
rect 11451 36420 11455 36476
rect 11455 36420 11511 36476
rect 11511 36420 11515 36476
rect 11451 36416 11515 36420
rect 11531 36476 11595 36480
rect 11531 36420 11535 36476
rect 11535 36420 11591 36476
rect 11591 36420 11595 36476
rect 11531 36416 11595 36420
rect 11611 36476 11675 36480
rect 11611 36420 11615 36476
rect 11615 36420 11671 36476
rect 11671 36420 11675 36476
rect 11611 36416 11675 36420
rect 18317 36476 18381 36480
rect 18317 36420 18321 36476
rect 18321 36420 18377 36476
rect 18377 36420 18381 36476
rect 18317 36416 18381 36420
rect 18397 36476 18461 36480
rect 18397 36420 18401 36476
rect 18401 36420 18457 36476
rect 18457 36420 18461 36476
rect 18397 36416 18461 36420
rect 18477 36476 18541 36480
rect 18477 36420 18481 36476
rect 18481 36420 18537 36476
rect 18537 36420 18541 36476
rect 18477 36416 18541 36420
rect 18557 36476 18621 36480
rect 18557 36420 18561 36476
rect 18561 36420 18617 36476
rect 18617 36420 18621 36476
rect 18557 36416 18621 36420
rect 25263 36476 25327 36480
rect 25263 36420 25267 36476
rect 25267 36420 25323 36476
rect 25323 36420 25327 36476
rect 25263 36416 25327 36420
rect 25343 36476 25407 36480
rect 25343 36420 25347 36476
rect 25347 36420 25403 36476
rect 25403 36420 25407 36476
rect 25343 36416 25407 36420
rect 25423 36476 25487 36480
rect 25423 36420 25427 36476
rect 25427 36420 25483 36476
rect 25483 36420 25487 36476
rect 25423 36416 25487 36420
rect 25503 36476 25567 36480
rect 25503 36420 25507 36476
rect 25507 36420 25563 36476
rect 25563 36420 25567 36476
rect 25503 36416 25567 36420
rect 7898 35932 7962 35936
rect 7898 35876 7902 35932
rect 7902 35876 7958 35932
rect 7958 35876 7962 35932
rect 7898 35872 7962 35876
rect 7978 35932 8042 35936
rect 7978 35876 7982 35932
rect 7982 35876 8038 35932
rect 8038 35876 8042 35932
rect 7978 35872 8042 35876
rect 8058 35932 8122 35936
rect 8058 35876 8062 35932
rect 8062 35876 8118 35932
rect 8118 35876 8122 35932
rect 8058 35872 8122 35876
rect 8138 35932 8202 35936
rect 8138 35876 8142 35932
rect 8142 35876 8198 35932
rect 8198 35876 8202 35932
rect 8138 35872 8202 35876
rect 14844 35932 14908 35936
rect 14844 35876 14848 35932
rect 14848 35876 14904 35932
rect 14904 35876 14908 35932
rect 14844 35872 14908 35876
rect 14924 35932 14988 35936
rect 14924 35876 14928 35932
rect 14928 35876 14984 35932
rect 14984 35876 14988 35932
rect 14924 35872 14988 35876
rect 15004 35932 15068 35936
rect 15004 35876 15008 35932
rect 15008 35876 15064 35932
rect 15064 35876 15068 35932
rect 15004 35872 15068 35876
rect 15084 35932 15148 35936
rect 15084 35876 15088 35932
rect 15088 35876 15144 35932
rect 15144 35876 15148 35932
rect 15084 35872 15148 35876
rect 21790 35932 21854 35936
rect 21790 35876 21794 35932
rect 21794 35876 21850 35932
rect 21850 35876 21854 35932
rect 21790 35872 21854 35876
rect 21870 35932 21934 35936
rect 21870 35876 21874 35932
rect 21874 35876 21930 35932
rect 21930 35876 21934 35932
rect 21870 35872 21934 35876
rect 21950 35932 22014 35936
rect 21950 35876 21954 35932
rect 21954 35876 22010 35932
rect 22010 35876 22014 35932
rect 21950 35872 22014 35876
rect 22030 35932 22094 35936
rect 22030 35876 22034 35932
rect 22034 35876 22090 35932
rect 22090 35876 22094 35932
rect 22030 35872 22094 35876
rect 28736 35932 28800 35936
rect 28736 35876 28740 35932
rect 28740 35876 28796 35932
rect 28796 35876 28800 35932
rect 28736 35872 28800 35876
rect 28816 35932 28880 35936
rect 28816 35876 28820 35932
rect 28820 35876 28876 35932
rect 28876 35876 28880 35932
rect 28816 35872 28880 35876
rect 28896 35932 28960 35936
rect 28896 35876 28900 35932
rect 28900 35876 28956 35932
rect 28956 35876 28960 35932
rect 28896 35872 28960 35876
rect 28976 35932 29040 35936
rect 28976 35876 28980 35932
rect 28980 35876 29036 35932
rect 29036 35876 29040 35932
rect 28976 35872 29040 35876
rect 4425 35388 4489 35392
rect 4425 35332 4429 35388
rect 4429 35332 4485 35388
rect 4485 35332 4489 35388
rect 4425 35328 4489 35332
rect 4505 35388 4569 35392
rect 4505 35332 4509 35388
rect 4509 35332 4565 35388
rect 4565 35332 4569 35388
rect 4505 35328 4569 35332
rect 4585 35388 4649 35392
rect 4585 35332 4589 35388
rect 4589 35332 4645 35388
rect 4645 35332 4649 35388
rect 4585 35328 4649 35332
rect 4665 35388 4729 35392
rect 4665 35332 4669 35388
rect 4669 35332 4725 35388
rect 4725 35332 4729 35388
rect 4665 35328 4729 35332
rect 11371 35388 11435 35392
rect 11371 35332 11375 35388
rect 11375 35332 11431 35388
rect 11431 35332 11435 35388
rect 11371 35328 11435 35332
rect 11451 35388 11515 35392
rect 11451 35332 11455 35388
rect 11455 35332 11511 35388
rect 11511 35332 11515 35388
rect 11451 35328 11515 35332
rect 11531 35388 11595 35392
rect 11531 35332 11535 35388
rect 11535 35332 11591 35388
rect 11591 35332 11595 35388
rect 11531 35328 11595 35332
rect 11611 35388 11675 35392
rect 11611 35332 11615 35388
rect 11615 35332 11671 35388
rect 11671 35332 11675 35388
rect 11611 35328 11675 35332
rect 18317 35388 18381 35392
rect 18317 35332 18321 35388
rect 18321 35332 18377 35388
rect 18377 35332 18381 35388
rect 18317 35328 18381 35332
rect 18397 35388 18461 35392
rect 18397 35332 18401 35388
rect 18401 35332 18457 35388
rect 18457 35332 18461 35388
rect 18397 35328 18461 35332
rect 18477 35388 18541 35392
rect 18477 35332 18481 35388
rect 18481 35332 18537 35388
rect 18537 35332 18541 35388
rect 18477 35328 18541 35332
rect 18557 35388 18621 35392
rect 18557 35332 18561 35388
rect 18561 35332 18617 35388
rect 18617 35332 18621 35388
rect 18557 35328 18621 35332
rect 25263 35388 25327 35392
rect 25263 35332 25267 35388
rect 25267 35332 25323 35388
rect 25323 35332 25327 35388
rect 25263 35328 25327 35332
rect 25343 35388 25407 35392
rect 25343 35332 25347 35388
rect 25347 35332 25403 35388
rect 25403 35332 25407 35388
rect 25343 35328 25407 35332
rect 25423 35388 25487 35392
rect 25423 35332 25427 35388
rect 25427 35332 25483 35388
rect 25483 35332 25487 35388
rect 25423 35328 25487 35332
rect 25503 35388 25567 35392
rect 25503 35332 25507 35388
rect 25507 35332 25563 35388
rect 25563 35332 25567 35388
rect 25503 35328 25567 35332
rect 7898 34844 7962 34848
rect 7898 34788 7902 34844
rect 7902 34788 7958 34844
rect 7958 34788 7962 34844
rect 7898 34784 7962 34788
rect 7978 34844 8042 34848
rect 7978 34788 7982 34844
rect 7982 34788 8038 34844
rect 8038 34788 8042 34844
rect 7978 34784 8042 34788
rect 8058 34844 8122 34848
rect 8058 34788 8062 34844
rect 8062 34788 8118 34844
rect 8118 34788 8122 34844
rect 8058 34784 8122 34788
rect 8138 34844 8202 34848
rect 8138 34788 8142 34844
rect 8142 34788 8198 34844
rect 8198 34788 8202 34844
rect 8138 34784 8202 34788
rect 14844 34844 14908 34848
rect 14844 34788 14848 34844
rect 14848 34788 14904 34844
rect 14904 34788 14908 34844
rect 14844 34784 14908 34788
rect 14924 34844 14988 34848
rect 14924 34788 14928 34844
rect 14928 34788 14984 34844
rect 14984 34788 14988 34844
rect 14924 34784 14988 34788
rect 15004 34844 15068 34848
rect 15004 34788 15008 34844
rect 15008 34788 15064 34844
rect 15064 34788 15068 34844
rect 15004 34784 15068 34788
rect 15084 34844 15148 34848
rect 15084 34788 15088 34844
rect 15088 34788 15144 34844
rect 15144 34788 15148 34844
rect 15084 34784 15148 34788
rect 21790 34844 21854 34848
rect 21790 34788 21794 34844
rect 21794 34788 21850 34844
rect 21850 34788 21854 34844
rect 21790 34784 21854 34788
rect 21870 34844 21934 34848
rect 21870 34788 21874 34844
rect 21874 34788 21930 34844
rect 21930 34788 21934 34844
rect 21870 34784 21934 34788
rect 21950 34844 22014 34848
rect 21950 34788 21954 34844
rect 21954 34788 22010 34844
rect 22010 34788 22014 34844
rect 21950 34784 22014 34788
rect 22030 34844 22094 34848
rect 22030 34788 22034 34844
rect 22034 34788 22090 34844
rect 22090 34788 22094 34844
rect 22030 34784 22094 34788
rect 28736 34844 28800 34848
rect 28736 34788 28740 34844
rect 28740 34788 28796 34844
rect 28796 34788 28800 34844
rect 28736 34784 28800 34788
rect 28816 34844 28880 34848
rect 28816 34788 28820 34844
rect 28820 34788 28876 34844
rect 28876 34788 28880 34844
rect 28816 34784 28880 34788
rect 28896 34844 28960 34848
rect 28896 34788 28900 34844
rect 28900 34788 28956 34844
rect 28956 34788 28960 34844
rect 28896 34784 28960 34788
rect 28976 34844 29040 34848
rect 28976 34788 28980 34844
rect 28980 34788 29036 34844
rect 29036 34788 29040 34844
rect 28976 34784 29040 34788
rect 4425 34300 4489 34304
rect 4425 34244 4429 34300
rect 4429 34244 4485 34300
rect 4485 34244 4489 34300
rect 4425 34240 4489 34244
rect 4505 34300 4569 34304
rect 4505 34244 4509 34300
rect 4509 34244 4565 34300
rect 4565 34244 4569 34300
rect 4505 34240 4569 34244
rect 4585 34300 4649 34304
rect 4585 34244 4589 34300
rect 4589 34244 4645 34300
rect 4645 34244 4649 34300
rect 4585 34240 4649 34244
rect 4665 34300 4729 34304
rect 4665 34244 4669 34300
rect 4669 34244 4725 34300
rect 4725 34244 4729 34300
rect 4665 34240 4729 34244
rect 11371 34300 11435 34304
rect 11371 34244 11375 34300
rect 11375 34244 11431 34300
rect 11431 34244 11435 34300
rect 11371 34240 11435 34244
rect 11451 34300 11515 34304
rect 11451 34244 11455 34300
rect 11455 34244 11511 34300
rect 11511 34244 11515 34300
rect 11451 34240 11515 34244
rect 11531 34300 11595 34304
rect 11531 34244 11535 34300
rect 11535 34244 11591 34300
rect 11591 34244 11595 34300
rect 11531 34240 11595 34244
rect 11611 34300 11675 34304
rect 11611 34244 11615 34300
rect 11615 34244 11671 34300
rect 11671 34244 11675 34300
rect 11611 34240 11675 34244
rect 18317 34300 18381 34304
rect 18317 34244 18321 34300
rect 18321 34244 18377 34300
rect 18377 34244 18381 34300
rect 18317 34240 18381 34244
rect 18397 34300 18461 34304
rect 18397 34244 18401 34300
rect 18401 34244 18457 34300
rect 18457 34244 18461 34300
rect 18397 34240 18461 34244
rect 18477 34300 18541 34304
rect 18477 34244 18481 34300
rect 18481 34244 18537 34300
rect 18537 34244 18541 34300
rect 18477 34240 18541 34244
rect 18557 34300 18621 34304
rect 18557 34244 18561 34300
rect 18561 34244 18617 34300
rect 18617 34244 18621 34300
rect 18557 34240 18621 34244
rect 25263 34300 25327 34304
rect 25263 34244 25267 34300
rect 25267 34244 25323 34300
rect 25323 34244 25327 34300
rect 25263 34240 25327 34244
rect 25343 34300 25407 34304
rect 25343 34244 25347 34300
rect 25347 34244 25403 34300
rect 25403 34244 25407 34300
rect 25343 34240 25407 34244
rect 25423 34300 25487 34304
rect 25423 34244 25427 34300
rect 25427 34244 25483 34300
rect 25483 34244 25487 34300
rect 25423 34240 25487 34244
rect 25503 34300 25567 34304
rect 25503 34244 25507 34300
rect 25507 34244 25563 34300
rect 25563 34244 25567 34300
rect 25503 34240 25567 34244
rect 7898 33756 7962 33760
rect 7898 33700 7902 33756
rect 7902 33700 7958 33756
rect 7958 33700 7962 33756
rect 7898 33696 7962 33700
rect 7978 33756 8042 33760
rect 7978 33700 7982 33756
rect 7982 33700 8038 33756
rect 8038 33700 8042 33756
rect 7978 33696 8042 33700
rect 8058 33756 8122 33760
rect 8058 33700 8062 33756
rect 8062 33700 8118 33756
rect 8118 33700 8122 33756
rect 8058 33696 8122 33700
rect 8138 33756 8202 33760
rect 8138 33700 8142 33756
rect 8142 33700 8198 33756
rect 8198 33700 8202 33756
rect 8138 33696 8202 33700
rect 14844 33756 14908 33760
rect 14844 33700 14848 33756
rect 14848 33700 14904 33756
rect 14904 33700 14908 33756
rect 14844 33696 14908 33700
rect 14924 33756 14988 33760
rect 14924 33700 14928 33756
rect 14928 33700 14984 33756
rect 14984 33700 14988 33756
rect 14924 33696 14988 33700
rect 15004 33756 15068 33760
rect 15004 33700 15008 33756
rect 15008 33700 15064 33756
rect 15064 33700 15068 33756
rect 15004 33696 15068 33700
rect 15084 33756 15148 33760
rect 15084 33700 15088 33756
rect 15088 33700 15144 33756
rect 15144 33700 15148 33756
rect 15084 33696 15148 33700
rect 21790 33756 21854 33760
rect 21790 33700 21794 33756
rect 21794 33700 21850 33756
rect 21850 33700 21854 33756
rect 21790 33696 21854 33700
rect 21870 33756 21934 33760
rect 21870 33700 21874 33756
rect 21874 33700 21930 33756
rect 21930 33700 21934 33756
rect 21870 33696 21934 33700
rect 21950 33756 22014 33760
rect 21950 33700 21954 33756
rect 21954 33700 22010 33756
rect 22010 33700 22014 33756
rect 21950 33696 22014 33700
rect 22030 33756 22094 33760
rect 22030 33700 22034 33756
rect 22034 33700 22090 33756
rect 22090 33700 22094 33756
rect 22030 33696 22094 33700
rect 28736 33756 28800 33760
rect 28736 33700 28740 33756
rect 28740 33700 28796 33756
rect 28796 33700 28800 33756
rect 28736 33696 28800 33700
rect 28816 33756 28880 33760
rect 28816 33700 28820 33756
rect 28820 33700 28876 33756
rect 28876 33700 28880 33756
rect 28816 33696 28880 33700
rect 28896 33756 28960 33760
rect 28896 33700 28900 33756
rect 28900 33700 28956 33756
rect 28956 33700 28960 33756
rect 28896 33696 28960 33700
rect 28976 33756 29040 33760
rect 28976 33700 28980 33756
rect 28980 33700 29036 33756
rect 29036 33700 29040 33756
rect 28976 33696 29040 33700
rect 4425 33212 4489 33216
rect 4425 33156 4429 33212
rect 4429 33156 4485 33212
rect 4485 33156 4489 33212
rect 4425 33152 4489 33156
rect 4505 33212 4569 33216
rect 4505 33156 4509 33212
rect 4509 33156 4565 33212
rect 4565 33156 4569 33212
rect 4505 33152 4569 33156
rect 4585 33212 4649 33216
rect 4585 33156 4589 33212
rect 4589 33156 4645 33212
rect 4645 33156 4649 33212
rect 4585 33152 4649 33156
rect 4665 33212 4729 33216
rect 4665 33156 4669 33212
rect 4669 33156 4725 33212
rect 4725 33156 4729 33212
rect 4665 33152 4729 33156
rect 11371 33212 11435 33216
rect 11371 33156 11375 33212
rect 11375 33156 11431 33212
rect 11431 33156 11435 33212
rect 11371 33152 11435 33156
rect 11451 33212 11515 33216
rect 11451 33156 11455 33212
rect 11455 33156 11511 33212
rect 11511 33156 11515 33212
rect 11451 33152 11515 33156
rect 11531 33212 11595 33216
rect 11531 33156 11535 33212
rect 11535 33156 11591 33212
rect 11591 33156 11595 33212
rect 11531 33152 11595 33156
rect 11611 33212 11675 33216
rect 11611 33156 11615 33212
rect 11615 33156 11671 33212
rect 11671 33156 11675 33212
rect 11611 33152 11675 33156
rect 18317 33212 18381 33216
rect 18317 33156 18321 33212
rect 18321 33156 18377 33212
rect 18377 33156 18381 33212
rect 18317 33152 18381 33156
rect 18397 33212 18461 33216
rect 18397 33156 18401 33212
rect 18401 33156 18457 33212
rect 18457 33156 18461 33212
rect 18397 33152 18461 33156
rect 18477 33212 18541 33216
rect 18477 33156 18481 33212
rect 18481 33156 18537 33212
rect 18537 33156 18541 33212
rect 18477 33152 18541 33156
rect 18557 33212 18621 33216
rect 18557 33156 18561 33212
rect 18561 33156 18617 33212
rect 18617 33156 18621 33212
rect 18557 33152 18621 33156
rect 25263 33212 25327 33216
rect 25263 33156 25267 33212
rect 25267 33156 25323 33212
rect 25323 33156 25327 33212
rect 25263 33152 25327 33156
rect 25343 33212 25407 33216
rect 25343 33156 25347 33212
rect 25347 33156 25403 33212
rect 25403 33156 25407 33212
rect 25343 33152 25407 33156
rect 25423 33212 25487 33216
rect 25423 33156 25427 33212
rect 25427 33156 25483 33212
rect 25483 33156 25487 33212
rect 25423 33152 25487 33156
rect 25503 33212 25567 33216
rect 25503 33156 25507 33212
rect 25507 33156 25563 33212
rect 25563 33156 25567 33212
rect 25503 33152 25567 33156
rect 7898 32668 7962 32672
rect 7898 32612 7902 32668
rect 7902 32612 7958 32668
rect 7958 32612 7962 32668
rect 7898 32608 7962 32612
rect 7978 32668 8042 32672
rect 7978 32612 7982 32668
rect 7982 32612 8038 32668
rect 8038 32612 8042 32668
rect 7978 32608 8042 32612
rect 8058 32668 8122 32672
rect 8058 32612 8062 32668
rect 8062 32612 8118 32668
rect 8118 32612 8122 32668
rect 8058 32608 8122 32612
rect 8138 32668 8202 32672
rect 8138 32612 8142 32668
rect 8142 32612 8198 32668
rect 8198 32612 8202 32668
rect 8138 32608 8202 32612
rect 14844 32668 14908 32672
rect 14844 32612 14848 32668
rect 14848 32612 14904 32668
rect 14904 32612 14908 32668
rect 14844 32608 14908 32612
rect 14924 32668 14988 32672
rect 14924 32612 14928 32668
rect 14928 32612 14984 32668
rect 14984 32612 14988 32668
rect 14924 32608 14988 32612
rect 15004 32668 15068 32672
rect 15004 32612 15008 32668
rect 15008 32612 15064 32668
rect 15064 32612 15068 32668
rect 15004 32608 15068 32612
rect 15084 32668 15148 32672
rect 15084 32612 15088 32668
rect 15088 32612 15144 32668
rect 15144 32612 15148 32668
rect 15084 32608 15148 32612
rect 21790 32668 21854 32672
rect 21790 32612 21794 32668
rect 21794 32612 21850 32668
rect 21850 32612 21854 32668
rect 21790 32608 21854 32612
rect 21870 32668 21934 32672
rect 21870 32612 21874 32668
rect 21874 32612 21930 32668
rect 21930 32612 21934 32668
rect 21870 32608 21934 32612
rect 21950 32668 22014 32672
rect 21950 32612 21954 32668
rect 21954 32612 22010 32668
rect 22010 32612 22014 32668
rect 21950 32608 22014 32612
rect 22030 32668 22094 32672
rect 22030 32612 22034 32668
rect 22034 32612 22090 32668
rect 22090 32612 22094 32668
rect 22030 32608 22094 32612
rect 28736 32668 28800 32672
rect 28736 32612 28740 32668
rect 28740 32612 28796 32668
rect 28796 32612 28800 32668
rect 28736 32608 28800 32612
rect 28816 32668 28880 32672
rect 28816 32612 28820 32668
rect 28820 32612 28876 32668
rect 28876 32612 28880 32668
rect 28816 32608 28880 32612
rect 28896 32668 28960 32672
rect 28896 32612 28900 32668
rect 28900 32612 28956 32668
rect 28956 32612 28960 32668
rect 28896 32608 28960 32612
rect 28976 32668 29040 32672
rect 28976 32612 28980 32668
rect 28980 32612 29036 32668
rect 29036 32612 29040 32668
rect 28976 32608 29040 32612
rect 4425 32124 4489 32128
rect 4425 32068 4429 32124
rect 4429 32068 4485 32124
rect 4485 32068 4489 32124
rect 4425 32064 4489 32068
rect 4505 32124 4569 32128
rect 4505 32068 4509 32124
rect 4509 32068 4565 32124
rect 4565 32068 4569 32124
rect 4505 32064 4569 32068
rect 4585 32124 4649 32128
rect 4585 32068 4589 32124
rect 4589 32068 4645 32124
rect 4645 32068 4649 32124
rect 4585 32064 4649 32068
rect 4665 32124 4729 32128
rect 4665 32068 4669 32124
rect 4669 32068 4725 32124
rect 4725 32068 4729 32124
rect 4665 32064 4729 32068
rect 11371 32124 11435 32128
rect 11371 32068 11375 32124
rect 11375 32068 11431 32124
rect 11431 32068 11435 32124
rect 11371 32064 11435 32068
rect 11451 32124 11515 32128
rect 11451 32068 11455 32124
rect 11455 32068 11511 32124
rect 11511 32068 11515 32124
rect 11451 32064 11515 32068
rect 11531 32124 11595 32128
rect 11531 32068 11535 32124
rect 11535 32068 11591 32124
rect 11591 32068 11595 32124
rect 11531 32064 11595 32068
rect 11611 32124 11675 32128
rect 11611 32068 11615 32124
rect 11615 32068 11671 32124
rect 11671 32068 11675 32124
rect 11611 32064 11675 32068
rect 18317 32124 18381 32128
rect 18317 32068 18321 32124
rect 18321 32068 18377 32124
rect 18377 32068 18381 32124
rect 18317 32064 18381 32068
rect 18397 32124 18461 32128
rect 18397 32068 18401 32124
rect 18401 32068 18457 32124
rect 18457 32068 18461 32124
rect 18397 32064 18461 32068
rect 18477 32124 18541 32128
rect 18477 32068 18481 32124
rect 18481 32068 18537 32124
rect 18537 32068 18541 32124
rect 18477 32064 18541 32068
rect 18557 32124 18621 32128
rect 18557 32068 18561 32124
rect 18561 32068 18617 32124
rect 18617 32068 18621 32124
rect 18557 32064 18621 32068
rect 25263 32124 25327 32128
rect 25263 32068 25267 32124
rect 25267 32068 25323 32124
rect 25323 32068 25327 32124
rect 25263 32064 25327 32068
rect 25343 32124 25407 32128
rect 25343 32068 25347 32124
rect 25347 32068 25403 32124
rect 25403 32068 25407 32124
rect 25343 32064 25407 32068
rect 25423 32124 25487 32128
rect 25423 32068 25427 32124
rect 25427 32068 25483 32124
rect 25483 32068 25487 32124
rect 25423 32064 25487 32068
rect 25503 32124 25567 32128
rect 25503 32068 25507 32124
rect 25507 32068 25563 32124
rect 25563 32068 25567 32124
rect 25503 32064 25567 32068
rect 7898 31580 7962 31584
rect 7898 31524 7902 31580
rect 7902 31524 7958 31580
rect 7958 31524 7962 31580
rect 7898 31520 7962 31524
rect 7978 31580 8042 31584
rect 7978 31524 7982 31580
rect 7982 31524 8038 31580
rect 8038 31524 8042 31580
rect 7978 31520 8042 31524
rect 8058 31580 8122 31584
rect 8058 31524 8062 31580
rect 8062 31524 8118 31580
rect 8118 31524 8122 31580
rect 8058 31520 8122 31524
rect 8138 31580 8202 31584
rect 8138 31524 8142 31580
rect 8142 31524 8198 31580
rect 8198 31524 8202 31580
rect 8138 31520 8202 31524
rect 14844 31580 14908 31584
rect 14844 31524 14848 31580
rect 14848 31524 14904 31580
rect 14904 31524 14908 31580
rect 14844 31520 14908 31524
rect 14924 31580 14988 31584
rect 14924 31524 14928 31580
rect 14928 31524 14984 31580
rect 14984 31524 14988 31580
rect 14924 31520 14988 31524
rect 15004 31580 15068 31584
rect 15004 31524 15008 31580
rect 15008 31524 15064 31580
rect 15064 31524 15068 31580
rect 15004 31520 15068 31524
rect 15084 31580 15148 31584
rect 15084 31524 15088 31580
rect 15088 31524 15144 31580
rect 15144 31524 15148 31580
rect 15084 31520 15148 31524
rect 21790 31580 21854 31584
rect 21790 31524 21794 31580
rect 21794 31524 21850 31580
rect 21850 31524 21854 31580
rect 21790 31520 21854 31524
rect 21870 31580 21934 31584
rect 21870 31524 21874 31580
rect 21874 31524 21930 31580
rect 21930 31524 21934 31580
rect 21870 31520 21934 31524
rect 21950 31580 22014 31584
rect 21950 31524 21954 31580
rect 21954 31524 22010 31580
rect 22010 31524 22014 31580
rect 21950 31520 22014 31524
rect 22030 31580 22094 31584
rect 22030 31524 22034 31580
rect 22034 31524 22090 31580
rect 22090 31524 22094 31580
rect 22030 31520 22094 31524
rect 28736 31580 28800 31584
rect 28736 31524 28740 31580
rect 28740 31524 28796 31580
rect 28796 31524 28800 31580
rect 28736 31520 28800 31524
rect 28816 31580 28880 31584
rect 28816 31524 28820 31580
rect 28820 31524 28876 31580
rect 28876 31524 28880 31580
rect 28816 31520 28880 31524
rect 28896 31580 28960 31584
rect 28896 31524 28900 31580
rect 28900 31524 28956 31580
rect 28956 31524 28960 31580
rect 28896 31520 28960 31524
rect 28976 31580 29040 31584
rect 28976 31524 28980 31580
rect 28980 31524 29036 31580
rect 29036 31524 29040 31580
rect 28976 31520 29040 31524
rect 4425 31036 4489 31040
rect 4425 30980 4429 31036
rect 4429 30980 4485 31036
rect 4485 30980 4489 31036
rect 4425 30976 4489 30980
rect 4505 31036 4569 31040
rect 4505 30980 4509 31036
rect 4509 30980 4565 31036
rect 4565 30980 4569 31036
rect 4505 30976 4569 30980
rect 4585 31036 4649 31040
rect 4585 30980 4589 31036
rect 4589 30980 4645 31036
rect 4645 30980 4649 31036
rect 4585 30976 4649 30980
rect 4665 31036 4729 31040
rect 4665 30980 4669 31036
rect 4669 30980 4725 31036
rect 4725 30980 4729 31036
rect 4665 30976 4729 30980
rect 11371 31036 11435 31040
rect 11371 30980 11375 31036
rect 11375 30980 11431 31036
rect 11431 30980 11435 31036
rect 11371 30976 11435 30980
rect 11451 31036 11515 31040
rect 11451 30980 11455 31036
rect 11455 30980 11511 31036
rect 11511 30980 11515 31036
rect 11451 30976 11515 30980
rect 11531 31036 11595 31040
rect 11531 30980 11535 31036
rect 11535 30980 11591 31036
rect 11591 30980 11595 31036
rect 11531 30976 11595 30980
rect 11611 31036 11675 31040
rect 11611 30980 11615 31036
rect 11615 30980 11671 31036
rect 11671 30980 11675 31036
rect 11611 30976 11675 30980
rect 18317 31036 18381 31040
rect 18317 30980 18321 31036
rect 18321 30980 18377 31036
rect 18377 30980 18381 31036
rect 18317 30976 18381 30980
rect 18397 31036 18461 31040
rect 18397 30980 18401 31036
rect 18401 30980 18457 31036
rect 18457 30980 18461 31036
rect 18397 30976 18461 30980
rect 18477 31036 18541 31040
rect 18477 30980 18481 31036
rect 18481 30980 18537 31036
rect 18537 30980 18541 31036
rect 18477 30976 18541 30980
rect 18557 31036 18621 31040
rect 18557 30980 18561 31036
rect 18561 30980 18617 31036
rect 18617 30980 18621 31036
rect 18557 30976 18621 30980
rect 25263 31036 25327 31040
rect 25263 30980 25267 31036
rect 25267 30980 25323 31036
rect 25323 30980 25327 31036
rect 25263 30976 25327 30980
rect 25343 31036 25407 31040
rect 25343 30980 25347 31036
rect 25347 30980 25403 31036
rect 25403 30980 25407 31036
rect 25343 30976 25407 30980
rect 25423 31036 25487 31040
rect 25423 30980 25427 31036
rect 25427 30980 25483 31036
rect 25483 30980 25487 31036
rect 25423 30976 25487 30980
rect 25503 31036 25567 31040
rect 25503 30980 25507 31036
rect 25507 30980 25563 31036
rect 25563 30980 25567 31036
rect 25503 30976 25567 30980
rect 7898 30492 7962 30496
rect 7898 30436 7902 30492
rect 7902 30436 7958 30492
rect 7958 30436 7962 30492
rect 7898 30432 7962 30436
rect 7978 30492 8042 30496
rect 7978 30436 7982 30492
rect 7982 30436 8038 30492
rect 8038 30436 8042 30492
rect 7978 30432 8042 30436
rect 8058 30492 8122 30496
rect 8058 30436 8062 30492
rect 8062 30436 8118 30492
rect 8118 30436 8122 30492
rect 8058 30432 8122 30436
rect 8138 30492 8202 30496
rect 8138 30436 8142 30492
rect 8142 30436 8198 30492
rect 8198 30436 8202 30492
rect 8138 30432 8202 30436
rect 14844 30492 14908 30496
rect 14844 30436 14848 30492
rect 14848 30436 14904 30492
rect 14904 30436 14908 30492
rect 14844 30432 14908 30436
rect 14924 30492 14988 30496
rect 14924 30436 14928 30492
rect 14928 30436 14984 30492
rect 14984 30436 14988 30492
rect 14924 30432 14988 30436
rect 15004 30492 15068 30496
rect 15004 30436 15008 30492
rect 15008 30436 15064 30492
rect 15064 30436 15068 30492
rect 15004 30432 15068 30436
rect 15084 30492 15148 30496
rect 15084 30436 15088 30492
rect 15088 30436 15144 30492
rect 15144 30436 15148 30492
rect 15084 30432 15148 30436
rect 21790 30492 21854 30496
rect 21790 30436 21794 30492
rect 21794 30436 21850 30492
rect 21850 30436 21854 30492
rect 21790 30432 21854 30436
rect 21870 30492 21934 30496
rect 21870 30436 21874 30492
rect 21874 30436 21930 30492
rect 21930 30436 21934 30492
rect 21870 30432 21934 30436
rect 21950 30492 22014 30496
rect 21950 30436 21954 30492
rect 21954 30436 22010 30492
rect 22010 30436 22014 30492
rect 21950 30432 22014 30436
rect 22030 30492 22094 30496
rect 22030 30436 22034 30492
rect 22034 30436 22090 30492
rect 22090 30436 22094 30492
rect 22030 30432 22094 30436
rect 28736 30492 28800 30496
rect 28736 30436 28740 30492
rect 28740 30436 28796 30492
rect 28796 30436 28800 30492
rect 28736 30432 28800 30436
rect 28816 30492 28880 30496
rect 28816 30436 28820 30492
rect 28820 30436 28876 30492
rect 28876 30436 28880 30492
rect 28816 30432 28880 30436
rect 28896 30492 28960 30496
rect 28896 30436 28900 30492
rect 28900 30436 28956 30492
rect 28956 30436 28960 30492
rect 28896 30432 28960 30436
rect 28976 30492 29040 30496
rect 28976 30436 28980 30492
rect 28980 30436 29036 30492
rect 29036 30436 29040 30492
rect 28976 30432 29040 30436
rect 4425 29948 4489 29952
rect 4425 29892 4429 29948
rect 4429 29892 4485 29948
rect 4485 29892 4489 29948
rect 4425 29888 4489 29892
rect 4505 29948 4569 29952
rect 4505 29892 4509 29948
rect 4509 29892 4565 29948
rect 4565 29892 4569 29948
rect 4505 29888 4569 29892
rect 4585 29948 4649 29952
rect 4585 29892 4589 29948
rect 4589 29892 4645 29948
rect 4645 29892 4649 29948
rect 4585 29888 4649 29892
rect 4665 29948 4729 29952
rect 4665 29892 4669 29948
rect 4669 29892 4725 29948
rect 4725 29892 4729 29948
rect 4665 29888 4729 29892
rect 11371 29948 11435 29952
rect 11371 29892 11375 29948
rect 11375 29892 11431 29948
rect 11431 29892 11435 29948
rect 11371 29888 11435 29892
rect 11451 29948 11515 29952
rect 11451 29892 11455 29948
rect 11455 29892 11511 29948
rect 11511 29892 11515 29948
rect 11451 29888 11515 29892
rect 11531 29948 11595 29952
rect 11531 29892 11535 29948
rect 11535 29892 11591 29948
rect 11591 29892 11595 29948
rect 11531 29888 11595 29892
rect 11611 29948 11675 29952
rect 11611 29892 11615 29948
rect 11615 29892 11671 29948
rect 11671 29892 11675 29948
rect 11611 29888 11675 29892
rect 18317 29948 18381 29952
rect 18317 29892 18321 29948
rect 18321 29892 18377 29948
rect 18377 29892 18381 29948
rect 18317 29888 18381 29892
rect 18397 29948 18461 29952
rect 18397 29892 18401 29948
rect 18401 29892 18457 29948
rect 18457 29892 18461 29948
rect 18397 29888 18461 29892
rect 18477 29948 18541 29952
rect 18477 29892 18481 29948
rect 18481 29892 18537 29948
rect 18537 29892 18541 29948
rect 18477 29888 18541 29892
rect 18557 29948 18621 29952
rect 18557 29892 18561 29948
rect 18561 29892 18617 29948
rect 18617 29892 18621 29948
rect 18557 29888 18621 29892
rect 25263 29948 25327 29952
rect 25263 29892 25267 29948
rect 25267 29892 25323 29948
rect 25323 29892 25327 29948
rect 25263 29888 25327 29892
rect 25343 29948 25407 29952
rect 25343 29892 25347 29948
rect 25347 29892 25403 29948
rect 25403 29892 25407 29948
rect 25343 29888 25407 29892
rect 25423 29948 25487 29952
rect 25423 29892 25427 29948
rect 25427 29892 25483 29948
rect 25483 29892 25487 29948
rect 25423 29888 25487 29892
rect 25503 29948 25567 29952
rect 25503 29892 25507 29948
rect 25507 29892 25563 29948
rect 25563 29892 25567 29948
rect 25503 29888 25567 29892
rect 7898 29404 7962 29408
rect 7898 29348 7902 29404
rect 7902 29348 7958 29404
rect 7958 29348 7962 29404
rect 7898 29344 7962 29348
rect 7978 29404 8042 29408
rect 7978 29348 7982 29404
rect 7982 29348 8038 29404
rect 8038 29348 8042 29404
rect 7978 29344 8042 29348
rect 8058 29404 8122 29408
rect 8058 29348 8062 29404
rect 8062 29348 8118 29404
rect 8118 29348 8122 29404
rect 8058 29344 8122 29348
rect 8138 29404 8202 29408
rect 8138 29348 8142 29404
rect 8142 29348 8198 29404
rect 8198 29348 8202 29404
rect 8138 29344 8202 29348
rect 14844 29404 14908 29408
rect 14844 29348 14848 29404
rect 14848 29348 14904 29404
rect 14904 29348 14908 29404
rect 14844 29344 14908 29348
rect 14924 29404 14988 29408
rect 14924 29348 14928 29404
rect 14928 29348 14984 29404
rect 14984 29348 14988 29404
rect 14924 29344 14988 29348
rect 15004 29404 15068 29408
rect 15004 29348 15008 29404
rect 15008 29348 15064 29404
rect 15064 29348 15068 29404
rect 15004 29344 15068 29348
rect 15084 29404 15148 29408
rect 15084 29348 15088 29404
rect 15088 29348 15144 29404
rect 15144 29348 15148 29404
rect 15084 29344 15148 29348
rect 21790 29404 21854 29408
rect 21790 29348 21794 29404
rect 21794 29348 21850 29404
rect 21850 29348 21854 29404
rect 21790 29344 21854 29348
rect 21870 29404 21934 29408
rect 21870 29348 21874 29404
rect 21874 29348 21930 29404
rect 21930 29348 21934 29404
rect 21870 29344 21934 29348
rect 21950 29404 22014 29408
rect 21950 29348 21954 29404
rect 21954 29348 22010 29404
rect 22010 29348 22014 29404
rect 21950 29344 22014 29348
rect 22030 29404 22094 29408
rect 22030 29348 22034 29404
rect 22034 29348 22090 29404
rect 22090 29348 22094 29404
rect 22030 29344 22094 29348
rect 28736 29404 28800 29408
rect 28736 29348 28740 29404
rect 28740 29348 28796 29404
rect 28796 29348 28800 29404
rect 28736 29344 28800 29348
rect 28816 29404 28880 29408
rect 28816 29348 28820 29404
rect 28820 29348 28876 29404
rect 28876 29348 28880 29404
rect 28816 29344 28880 29348
rect 28896 29404 28960 29408
rect 28896 29348 28900 29404
rect 28900 29348 28956 29404
rect 28956 29348 28960 29404
rect 28896 29344 28960 29348
rect 28976 29404 29040 29408
rect 28976 29348 28980 29404
rect 28980 29348 29036 29404
rect 29036 29348 29040 29404
rect 28976 29344 29040 29348
rect 4425 28860 4489 28864
rect 4425 28804 4429 28860
rect 4429 28804 4485 28860
rect 4485 28804 4489 28860
rect 4425 28800 4489 28804
rect 4505 28860 4569 28864
rect 4505 28804 4509 28860
rect 4509 28804 4565 28860
rect 4565 28804 4569 28860
rect 4505 28800 4569 28804
rect 4585 28860 4649 28864
rect 4585 28804 4589 28860
rect 4589 28804 4645 28860
rect 4645 28804 4649 28860
rect 4585 28800 4649 28804
rect 4665 28860 4729 28864
rect 4665 28804 4669 28860
rect 4669 28804 4725 28860
rect 4725 28804 4729 28860
rect 4665 28800 4729 28804
rect 11371 28860 11435 28864
rect 11371 28804 11375 28860
rect 11375 28804 11431 28860
rect 11431 28804 11435 28860
rect 11371 28800 11435 28804
rect 11451 28860 11515 28864
rect 11451 28804 11455 28860
rect 11455 28804 11511 28860
rect 11511 28804 11515 28860
rect 11451 28800 11515 28804
rect 11531 28860 11595 28864
rect 11531 28804 11535 28860
rect 11535 28804 11591 28860
rect 11591 28804 11595 28860
rect 11531 28800 11595 28804
rect 11611 28860 11675 28864
rect 11611 28804 11615 28860
rect 11615 28804 11671 28860
rect 11671 28804 11675 28860
rect 11611 28800 11675 28804
rect 18317 28860 18381 28864
rect 18317 28804 18321 28860
rect 18321 28804 18377 28860
rect 18377 28804 18381 28860
rect 18317 28800 18381 28804
rect 18397 28860 18461 28864
rect 18397 28804 18401 28860
rect 18401 28804 18457 28860
rect 18457 28804 18461 28860
rect 18397 28800 18461 28804
rect 18477 28860 18541 28864
rect 18477 28804 18481 28860
rect 18481 28804 18537 28860
rect 18537 28804 18541 28860
rect 18477 28800 18541 28804
rect 18557 28860 18621 28864
rect 18557 28804 18561 28860
rect 18561 28804 18617 28860
rect 18617 28804 18621 28860
rect 18557 28800 18621 28804
rect 25263 28860 25327 28864
rect 25263 28804 25267 28860
rect 25267 28804 25323 28860
rect 25323 28804 25327 28860
rect 25263 28800 25327 28804
rect 25343 28860 25407 28864
rect 25343 28804 25347 28860
rect 25347 28804 25403 28860
rect 25403 28804 25407 28860
rect 25343 28800 25407 28804
rect 25423 28860 25487 28864
rect 25423 28804 25427 28860
rect 25427 28804 25483 28860
rect 25483 28804 25487 28860
rect 25423 28800 25487 28804
rect 25503 28860 25567 28864
rect 25503 28804 25507 28860
rect 25507 28804 25563 28860
rect 25563 28804 25567 28860
rect 25503 28800 25567 28804
rect 7898 28316 7962 28320
rect 7898 28260 7902 28316
rect 7902 28260 7958 28316
rect 7958 28260 7962 28316
rect 7898 28256 7962 28260
rect 7978 28316 8042 28320
rect 7978 28260 7982 28316
rect 7982 28260 8038 28316
rect 8038 28260 8042 28316
rect 7978 28256 8042 28260
rect 8058 28316 8122 28320
rect 8058 28260 8062 28316
rect 8062 28260 8118 28316
rect 8118 28260 8122 28316
rect 8058 28256 8122 28260
rect 8138 28316 8202 28320
rect 8138 28260 8142 28316
rect 8142 28260 8198 28316
rect 8198 28260 8202 28316
rect 8138 28256 8202 28260
rect 14844 28316 14908 28320
rect 14844 28260 14848 28316
rect 14848 28260 14904 28316
rect 14904 28260 14908 28316
rect 14844 28256 14908 28260
rect 14924 28316 14988 28320
rect 14924 28260 14928 28316
rect 14928 28260 14984 28316
rect 14984 28260 14988 28316
rect 14924 28256 14988 28260
rect 15004 28316 15068 28320
rect 15004 28260 15008 28316
rect 15008 28260 15064 28316
rect 15064 28260 15068 28316
rect 15004 28256 15068 28260
rect 15084 28316 15148 28320
rect 15084 28260 15088 28316
rect 15088 28260 15144 28316
rect 15144 28260 15148 28316
rect 15084 28256 15148 28260
rect 21790 28316 21854 28320
rect 21790 28260 21794 28316
rect 21794 28260 21850 28316
rect 21850 28260 21854 28316
rect 21790 28256 21854 28260
rect 21870 28316 21934 28320
rect 21870 28260 21874 28316
rect 21874 28260 21930 28316
rect 21930 28260 21934 28316
rect 21870 28256 21934 28260
rect 21950 28316 22014 28320
rect 21950 28260 21954 28316
rect 21954 28260 22010 28316
rect 22010 28260 22014 28316
rect 21950 28256 22014 28260
rect 22030 28316 22094 28320
rect 22030 28260 22034 28316
rect 22034 28260 22090 28316
rect 22090 28260 22094 28316
rect 22030 28256 22094 28260
rect 28736 28316 28800 28320
rect 28736 28260 28740 28316
rect 28740 28260 28796 28316
rect 28796 28260 28800 28316
rect 28736 28256 28800 28260
rect 28816 28316 28880 28320
rect 28816 28260 28820 28316
rect 28820 28260 28876 28316
rect 28876 28260 28880 28316
rect 28816 28256 28880 28260
rect 28896 28316 28960 28320
rect 28896 28260 28900 28316
rect 28900 28260 28956 28316
rect 28956 28260 28960 28316
rect 28896 28256 28960 28260
rect 28976 28316 29040 28320
rect 28976 28260 28980 28316
rect 28980 28260 29036 28316
rect 29036 28260 29040 28316
rect 28976 28256 29040 28260
rect 4425 27772 4489 27776
rect 4425 27716 4429 27772
rect 4429 27716 4485 27772
rect 4485 27716 4489 27772
rect 4425 27712 4489 27716
rect 4505 27772 4569 27776
rect 4505 27716 4509 27772
rect 4509 27716 4565 27772
rect 4565 27716 4569 27772
rect 4505 27712 4569 27716
rect 4585 27772 4649 27776
rect 4585 27716 4589 27772
rect 4589 27716 4645 27772
rect 4645 27716 4649 27772
rect 4585 27712 4649 27716
rect 4665 27772 4729 27776
rect 4665 27716 4669 27772
rect 4669 27716 4725 27772
rect 4725 27716 4729 27772
rect 4665 27712 4729 27716
rect 11371 27772 11435 27776
rect 11371 27716 11375 27772
rect 11375 27716 11431 27772
rect 11431 27716 11435 27772
rect 11371 27712 11435 27716
rect 11451 27772 11515 27776
rect 11451 27716 11455 27772
rect 11455 27716 11511 27772
rect 11511 27716 11515 27772
rect 11451 27712 11515 27716
rect 11531 27772 11595 27776
rect 11531 27716 11535 27772
rect 11535 27716 11591 27772
rect 11591 27716 11595 27772
rect 11531 27712 11595 27716
rect 11611 27772 11675 27776
rect 11611 27716 11615 27772
rect 11615 27716 11671 27772
rect 11671 27716 11675 27772
rect 11611 27712 11675 27716
rect 18317 27772 18381 27776
rect 18317 27716 18321 27772
rect 18321 27716 18377 27772
rect 18377 27716 18381 27772
rect 18317 27712 18381 27716
rect 18397 27772 18461 27776
rect 18397 27716 18401 27772
rect 18401 27716 18457 27772
rect 18457 27716 18461 27772
rect 18397 27712 18461 27716
rect 18477 27772 18541 27776
rect 18477 27716 18481 27772
rect 18481 27716 18537 27772
rect 18537 27716 18541 27772
rect 18477 27712 18541 27716
rect 18557 27772 18621 27776
rect 18557 27716 18561 27772
rect 18561 27716 18617 27772
rect 18617 27716 18621 27772
rect 18557 27712 18621 27716
rect 25263 27772 25327 27776
rect 25263 27716 25267 27772
rect 25267 27716 25323 27772
rect 25323 27716 25327 27772
rect 25263 27712 25327 27716
rect 25343 27772 25407 27776
rect 25343 27716 25347 27772
rect 25347 27716 25403 27772
rect 25403 27716 25407 27772
rect 25343 27712 25407 27716
rect 25423 27772 25487 27776
rect 25423 27716 25427 27772
rect 25427 27716 25483 27772
rect 25483 27716 25487 27772
rect 25423 27712 25487 27716
rect 25503 27772 25567 27776
rect 25503 27716 25507 27772
rect 25507 27716 25563 27772
rect 25563 27716 25567 27772
rect 25503 27712 25567 27716
rect 7898 27228 7962 27232
rect 7898 27172 7902 27228
rect 7902 27172 7958 27228
rect 7958 27172 7962 27228
rect 7898 27168 7962 27172
rect 7978 27228 8042 27232
rect 7978 27172 7982 27228
rect 7982 27172 8038 27228
rect 8038 27172 8042 27228
rect 7978 27168 8042 27172
rect 8058 27228 8122 27232
rect 8058 27172 8062 27228
rect 8062 27172 8118 27228
rect 8118 27172 8122 27228
rect 8058 27168 8122 27172
rect 8138 27228 8202 27232
rect 8138 27172 8142 27228
rect 8142 27172 8198 27228
rect 8198 27172 8202 27228
rect 8138 27168 8202 27172
rect 14844 27228 14908 27232
rect 14844 27172 14848 27228
rect 14848 27172 14904 27228
rect 14904 27172 14908 27228
rect 14844 27168 14908 27172
rect 14924 27228 14988 27232
rect 14924 27172 14928 27228
rect 14928 27172 14984 27228
rect 14984 27172 14988 27228
rect 14924 27168 14988 27172
rect 15004 27228 15068 27232
rect 15004 27172 15008 27228
rect 15008 27172 15064 27228
rect 15064 27172 15068 27228
rect 15004 27168 15068 27172
rect 15084 27228 15148 27232
rect 15084 27172 15088 27228
rect 15088 27172 15144 27228
rect 15144 27172 15148 27228
rect 15084 27168 15148 27172
rect 21790 27228 21854 27232
rect 21790 27172 21794 27228
rect 21794 27172 21850 27228
rect 21850 27172 21854 27228
rect 21790 27168 21854 27172
rect 21870 27228 21934 27232
rect 21870 27172 21874 27228
rect 21874 27172 21930 27228
rect 21930 27172 21934 27228
rect 21870 27168 21934 27172
rect 21950 27228 22014 27232
rect 21950 27172 21954 27228
rect 21954 27172 22010 27228
rect 22010 27172 22014 27228
rect 21950 27168 22014 27172
rect 22030 27228 22094 27232
rect 22030 27172 22034 27228
rect 22034 27172 22090 27228
rect 22090 27172 22094 27228
rect 22030 27168 22094 27172
rect 28736 27228 28800 27232
rect 28736 27172 28740 27228
rect 28740 27172 28796 27228
rect 28796 27172 28800 27228
rect 28736 27168 28800 27172
rect 28816 27228 28880 27232
rect 28816 27172 28820 27228
rect 28820 27172 28876 27228
rect 28876 27172 28880 27228
rect 28816 27168 28880 27172
rect 28896 27228 28960 27232
rect 28896 27172 28900 27228
rect 28900 27172 28956 27228
rect 28956 27172 28960 27228
rect 28896 27168 28960 27172
rect 28976 27228 29040 27232
rect 28976 27172 28980 27228
rect 28980 27172 29036 27228
rect 29036 27172 29040 27228
rect 28976 27168 29040 27172
rect 4425 26684 4489 26688
rect 4425 26628 4429 26684
rect 4429 26628 4485 26684
rect 4485 26628 4489 26684
rect 4425 26624 4489 26628
rect 4505 26684 4569 26688
rect 4505 26628 4509 26684
rect 4509 26628 4565 26684
rect 4565 26628 4569 26684
rect 4505 26624 4569 26628
rect 4585 26684 4649 26688
rect 4585 26628 4589 26684
rect 4589 26628 4645 26684
rect 4645 26628 4649 26684
rect 4585 26624 4649 26628
rect 4665 26684 4729 26688
rect 4665 26628 4669 26684
rect 4669 26628 4725 26684
rect 4725 26628 4729 26684
rect 4665 26624 4729 26628
rect 11371 26684 11435 26688
rect 11371 26628 11375 26684
rect 11375 26628 11431 26684
rect 11431 26628 11435 26684
rect 11371 26624 11435 26628
rect 11451 26684 11515 26688
rect 11451 26628 11455 26684
rect 11455 26628 11511 26684
rect 11511 26628 11515 26684
rect 11451 26624 11515 26628
rect 11531 26684 11595 26688
rect 11531 26628 11535 26684
rect 11535 26628 11591 26684
rect 11591 26628 11595 26684
rect 11531 26624 11595 26628
rect 11611 26684 11675 26688
rect 11611 26628 11615 26684
rect 11615 26628 11671 26684
rect 11671 26628 11675 26684
rect 11611 26624 11675 26628
rect 18317 26684 18381 26688
rect 18317 26628 18321 26684
rect 18321 26628 18377 26684
rect 18377 26628 18381 26684
rect 18317 26624 18381 26628
rect 18397 26684 18461 26688
rect 18397 26628 18401 26684
rect 18401 26628 18457 26684
rect 18457 26628 18461 26684
rect 18397 26624 18461 26628
rect 18477 26684 18541 26688
rect 18477 26628 18481 26684
rect 18481 26628 18537 26684
rect 18537 26628 18541 26684
rect 18477 26624 18541 26628
rect 18557 26684 18621 26688
rect 18557 26628 18561 26684
rect 18561 26628 18617 26684
rect 18617 26628 18621 26684
rect 18557 26624 18621 26628
rect 25263 26684 25327 26688
rect 25263 26628 25267 26684
rect 25267 26628 25323 26684
rect 25323 26628 25327 26684
rect 25263 26624 25327 26628
rect 25343 26684 25407 26688
rect 25343 26628 25347 26684
rect 25347 26628 25403 26684
rect 25403 26628 25407 26684
rect 25343 26624 25407 26628
rect 25423 26684 25487 26688
rect 25423 26628 25427 26684
rect 25427 26628 25483 26684
rect 25483 26628 25487 26684
rect 25423 26624 25487 26628
rect 25503 26684 25567 26688
rect 25503 26628 25507 26684
rect 25507 26628 25563 26684
rect 25563 26628 25567 26684
rect 25503 26624 25567 26628
rect 7898 26140 7962 26144
rect 7898 26084 7902 26140
rect 7902 26084 7958 26140
rect 7958 26084 7962 26140
rect 7898 26080 7962 26084
rect 7978 26140 8042 26144
rect 7978 26084 7982 26140
rect 7982 26084 8038 26140
rect 8038 26084 8042 26140
rect 7978 26080 8042 26084
rect 8058 26140 8122 26144
rect 8058 26084 8062 26140
rect 8062 26084 8118 26140
rect 8118 26084 8122 26140
rect 8058 26080 8122 26084
rect 8138 26140 8202 26144
rect 8138 26084 8142 26140
rect 8142 26084 8198 26140
rect 8198 26084 8202 26140
rect 8138 26080 8202 26084
rect 14844 26140 14908 26144
rect 14844 26084 14848 26140
rect 14848 26084 14904 26140
rect 14904 26084 14908 26140
rect 14844 26080 14908 26084
rect 14924 26140 14988 26144
rect 14924 26084 14928 26140
rect 14928 26084 14984 26140
rect 14984 26084 14988 26140
rect 14924 26080 14988 26084
rect 15004 26140 15068 26144
rect 15004 26084 15008 26140
rect 15008 26084 15064 26140
rect 15064 26084 15068 26140
rect 15004 26080 15068 26084
rect 15084 26140 15148 26144
rect 15084 26084 15088 26140
rect 15088 26084 15144 26140
rect 15144 26084 15148 26140
rect 15084 26080 15148 26084
rect 21790 26140 21854 26144
rect 21790 26084 21794 26140
rect 21794 26084 21850 26140
rect 21850 26084 21854 26140
rect 21790 26080 21854 26084
rect 21870 26140 21934 26144
rect 21870 26084 21874 26140
rect 21874 26084 21930 26140
rect 21930 26084 21934 26140
rect 21870 26080 21934 26084
rect 21950 26140 22014 26144
rect 21950 26084 21954 26140
rect 21954 26084 22010 26140
rect 22010 26084 22014 26140
rect 21950 26080 22014 26084
rect 22030 26140 22094 26144
rect 22030 26084 22034 26140
rect 22034 26084 22090 26140
rect 22090 26084 22094 26140
rect 22030 26080 22094 26084
rect 28736 26140 28800 26144
rect 28736 26084 28740 26140
rect 28740 26084 28796 26140
rect 28796 26084 28800 26140
rect 28736 26080 28800 26084
rect 28816 26140 28880 26144
rect 28816 26084 28820 26140
rect 28820 26084 28876 26140
rect 28876 26084 28880 26140
rect 28816 26080 28880 26084
rect 28896 26140 28960 26144
rect 28896 26084 28900 26140
rect 28900 26084 28956 26140
rect 28956 26084 28960 26140
rect 28896 26080 28960 26084
rect 28976 26140 29040 26144
rect 28976 26084 28980 26140
rect 28980 26084 29036 26140
rect 29036 26084 29040 26140
rect 28976 26080 29040 26084
rect 4425 25596 4489 25600
rect 4425 25540 4429 25596
rect 4429 25540 4485 25596
rect 4485 25540 4489 25596
rect 4425 25536 4489 25540
rect 4505 25596 4569 25600
rect 4505 25540 4509 25596
rect 4509 25540 4565 25596
rect 4565 25540 4569 25596
rect 4505 25536 4569 25540
rect 4585 25596 4649 25600
rect 4585 25540 4589 25596
rect 4589 25540 4645 25596
rect 4645 25540 4649 25596
rect 4585 25536 4649 25540
rect 4665 25596 4729 25600
rect 4665 25540 4669 25596
rect 4669 25540 4725 25596
rect 4725 25540 4729 25596
rect 4665 25536 4729 25540
rect 11371 25596 11435 25600
rect 11371 25540 11375 25596
rect 11375 25540 11431 25596
rect 11431 25540 11435 25596
rect 11371 25536 11435 25540
rect 11451 25596 11515 25600
rect 11451 25540 11455 25596
rect 11455 25540 11511 25596
rect 11511 25540 11515 25596
rect 11451 25536 11515 25540
rect 11531 25596 11595 25600
rect 11531 25540 11535 25596
rect 11535 25540 11591 25596
rect 11591 25540 11595 25596
rect 11531 25536 11595 25540
rect 11611 25596 11675 25600
rect 11611 25540 11615 25596
rect 11615 25540 11671 25596
rect 11671 25540 11675 25596
rect 11611 25536 11675 25540
rect 18317 25596 18381 25600
rect 18317 25540 18321 25596
rect 18321 25540 18377 25596
rect 18377 25540 18381 25596
rect 18317 25536 18381 25540
rect 18397 25596 18461 25600
rect 18397 25540 18401 25596
rect 18401 25540 18457 25596
rect 18457 25540 18461 25596
rect 18397 25536 18461 25540
rect 18477 25596 18541 25600
rect 18477 25540 18481 25596
rect 18481 25540 18537 25596
rect 18537 25540 18541 25596
rect 18477 25536 18541 25540
rect 18557 25596 18621 25600
rect 18557 25540 18561 25596
rect 18561 25540 18617 25596
rect 18617 25540 18621 25596
rect 18557 25536 18621 25540
rect 25263 25596 25327 25600
rect 25263 25540 25267 25596
rect 25267 25540 25323 25596
rect 25323 25540 25327 25596
rect 25263 25536 25327 25540
rect 25343 25596 25407 25600
rect 25343 25540 25347 25596
rect 25347 25540 25403 25596
rect 25403 25540 25407 25596
rect 25343 25536 25407 25540
rect 25423 25596 25487 25600
rect 25423 25540 25427 25596
rect 25427 25540 25483 25596
rect 25483 25540 25487 25596
rect 25423 25536 25487 25540
rect 25503 25596 25567 25600
rect 25503 25540 25507 25596
rect 25507 25540 25563 25596
rect 25563 25540 25567 25596
rect 25503 25536 25567 25540
rect 7898 25052 7962 25056
rect 7898 24996 7902 25052
rect 7902 24996 7958 25052
rect 7958 24996 7962 25052
rect 7898 24992 7962 24996
rect 7978 25052 8042 25056
rect 7978 24996 7982 25052
rect 7982 24996 8038 25052
rect 8038 24996 8042 25052
rect 7978 24992 8042 24996
rect 8058 25052 8122 25056
rect 8058 24996 8062 25052
rect 8062 24996 8118 25052
rect 8118 24996 8122 25052
rect 8058 24992 8122 24996
rect 8138 25052 8202 25056
rect 8138 24996 8142 25052
rect 8142 24996 8198 25052
rect 8198 24996 8202 25052
rect 8138 24992 8202 24996
rect 14844 25052 14908 25056
rect 14844 24996 14848 25052
rect 14848 24996 14904 25052
rect 14904 24996 14908 25052
rect 14844 24992 14908 24996
rect 14924 25052 14988 25056
rect 14924 24996 14928 25052
rect 14928 24996 14984 25052
rect 14984 24996 14988 25052
rect 14924 24992 14988 24996
rect 15004 25052 15068 25056
rect 15004 24996 15008 25052
rect 15008 24996 15064 25052
rect 15064 24996 15068 25052
rect 15004 24992 15068 24996
rect 15084 25052 15148 25056
rect 15084 24996 15088 25052
rect 15088 24996 15144 25052
rect 15144 24996 15148 25052
rect 15084 24992 15148 24996
rect 21790 25052 21854 25056
rect 21790 24996 21794 25052
rect 21794 24996 21850 25052
rect 21850 24996 21854 25052
rect 21790 24992 21854 24996
rect 21870 25052 21934 25056
rect 21870 24996 21874 25052
rect 21874 24996 21930 25052
rect 21930 24996 21934 25052
rect 21870 24992 21934 24996
rect 21950 25052 22014 25056
rect 21950 24996 21954 25052
rect 21954 24996 22010 25052
rect 22010 24996 22014 25052
rect 21950 24992 22014 24996
rect 22030 25052 22094 25056
rect 22030 24996 22034 25052
rect 22034 24996 22090 25052
rect 22090 24996 22094 25052
rect 22030 24992 22094 24996
rect 28736 25052 28800 25056
rect 28736 24996 28740 25052
rect 28740 24996 28796 25052
rect 28796 24996 28800 25052
rect 28736 24992 28800 24996
rect 28816 25052 28880 25056
rect 28816 24996 28820 25052
rect 28820 24996 28876 25052
rect 28876 24996 28880 25052
rect 28816 24992 28880 24996
rect 28896 25052 28960 25056
rect 28896 24996 28900 25052
rect 28900 24996 28956 25052
rect 28956 24996 28960 25052
rect 28896 24992 28960 24996
rect 28976 25052 29040 25056
rect 28976 24996 28980 25052
rect 28980 24996 29036 25052
rect 29036 24996 29040 25052
rect 28976 24992 29040 24996
rect 19564 24652 19628 24716
rect 4425 24508 4489 24512
rect 4425 24452 4429 24508
rect 4429 24452 4485 24508
rect 4485 24452 4489 24508
rect 4425 24448 4489 24452
rect 4505 24508 4569 24512
rect 4505 24452 4509 24508
rect 4509 24452 4565 24508
rect 4565 24452 4569 24508
rect 4505 24448 4569 24452
rect 4585 24508 4649 24512
rect 4585 24452 4589 24508
rect 4589 24452 4645 24508
rect 4645 24452 4649 24508
rect 4585 24448 4649 24452
rect 4665 24508 4729 24512
rect 4665 24452 4669 24508
rect 4669 24452 4725 24508
rect 4725 24452 4729 24508
rect 4665 24448 4729 24452
rect 11371 24508 11435 24512
rect 11371 24452 11375 24508
rect 11375 24452 11431 24508
rect 11431 24452 11435 24508
rect 11371 24448 11435 24452
rect 11451 24508 11515 24512
rect 11451 24452 11455 24508
rect 11455 24452 11511 24508
rect 11511 24452 11515 24508
rect 11451 24448 11515 24452
rect 11531 24508 11595 24512
rect 11531 24452 11535 24508
rect 11535 24452 11591 24508
rect 11591 24452 11595 24508
rect 11531 24448 11595 24452
rect 11611 24508 11675 24512
rect 11611 24452 11615 24508
rect 11615 24452 11671 24508
rect 11671 24452 11675 24508
rect 11611 24448 11675 24452
rect 18317 24508 18381 24512
rect 18317 24452 18321 24508
rect 18321 24452 18377 24508
rect 18377 24452 18381 24508
rect 18317 24448 18381 24452
rect 18397 24508 18461 24512
rect 18397 24452 18401 24508
rect 18401 24452 18457 24508
rect 18457 24452 18461 24508
rect 18397 24448 18461 24452
rect 18477 24508 18541 24512
rect 18477 24452 18481 24508
rect 18481 24452 18537 24508
rect 18537 24452 18541 24508
rect 18477 24448 18541 24452
rect 18557 24508 18621 24512
rect 18557 24452 18561 24508
rect 18561 24452 18617 24508
rect 18617 24452 18621 24508
rect 18557 24448 18621 24452
rect 25263 24508 25327 24512
rect 25263 24452 25267 24508
rect 25267 24452 25323 24508
rect 25323 24452 25327 24508
rect 25263 24448 25327 24452
rect 25343 24508 25407 24512
rect 25343 24452 25347 24508
rect 25347 24452 25403 24508
rect 25403 24452 25407 24508
rect 25343 24448 25407 24452
rect 25423 24508 25487 24512
rect 25423 24452 25427 24508
rect 25427 24452 25483 24508
rect 25483 24452 25487 24508
rect 25423 24448 25487 24452
rect 25503 24508 25567 24512
rect 25503 24452 25507 24508
rect 25507 24452 25563 24508
rect 25563 24452 25567 24508
rect 25503 24448 25567 24452
rect 7898 23964 7962 23968
rect 7898 23908 7902 23964
rect 7902 23908 7958 23964
rect 7958 23908 7962 23964
rect 7898 23904 7962 23908
rect 7978 23964 8042 23968
rect 7978 23908 7982 23964
rect 7982 23908 8038 23964
rect 8038 23908 8042 23964
rect 7978 23904 8042 23908
rect 8058 23964 8122 23968
rect 8058 23908 8062 23964
rect 8062 23908 8118 23964
rect 8118 23908 8122 23964
rect 8058 23904 8122 23908
rect 8138 23964 8202 23968
rect 8138 23908 8142 23964
rect 8142 23908 8198 23964
rect 8198 23908 8202 23964
rect 8138 23904 8202 23908
rect 14844 23964 14908 23968
rect 14844 23908 14848 23964
rect 14848 23908 14904 23964
rect 14904 23908 14908 23964
rect 14844 23904 14908 23908
rect 14924 23964 14988 23968
rect 14924 23908 14928 23964
rect 14928 23908 14984 23964
rect 14984 23908 14988 23964
rect 14924 23904 14988 23908
rect 15004 23964 15068 23968
rect 15004 23908 15008 23964
rect 15008 23908 15064 23964
rect 15064 23908 15068 23964
rect 15004 23904 15068 23908
rect 15084 23964 15148 23968
rect 15084 23908 15088 23964
rect 15088 23908 15144 23964
rect 15144 23908 15148 23964
rect 15084 23904 15148 23908
rect 21790 23964 21854 23968
rect 21790 23908 21794 23964
rect 21794 23908 21850 23964
rect 21850 23908 21854 23964
rect 21790 23904 21854 23908
rect 21870 23964 21934 23968
rect 21870 23908 21874 23964
rect 21874 23908 21930 23964
rect 21930 23908 21934 23964
rect 21870 23904 21934 23908
rect 21950 23964 22014 23968
rect 21950 23908 21954 23964
rect 21954 23908 22010 23964
rect 22010 23908 22014 23964
rect 21950 23904 22014 23908
rect 22030 23964 22094 23968
rect 22030 23908 22034 23964
rect 22034 23908 22090 23964
rect 22090 23908 22094 23964
rect 22030 23904 22094 23908
rect 28736 23964 28800 23968
rect 28736 23908 28740 23964
rect 28740 23908 28796 23964
rect 28796 23908 28800 23964
rect 28736 23904 28800 23908
rect 28816 23964 28880 23968
rect 28816 23908 28820 23964
rect 28820 23908 28876 23964
rect 28876 23908 28880 23964
rect 28816 23904 28880 23908
rect 28896 23964 28960 23968
rect 28896 23908 28900 23964
rect 28900 23908 28956 23964
rect 28956 23908 28960 23964
rect 28896 23904 28960 23908
rect 28976 23964 29040 23968
rect 28976 23908 28980 23964
rect 28980 23908 29036 23964
rect 29036 23908 29040 23964
rect 28976 23904 29040 23908
rect 4425 23420 4489 23424
rect 4425 23364 4429 23420
rect 4429 23364 4485 23420
rect 4485 23364 4489 23420
rect 4425 23360 4489 23364
rect 4505 23420 4569 23424
rect 4505 23364 4509 23420
rect 4509 23364 4565 23420
rect 4565 23364 4569 23420
rect 4505 23360 4569 23364
rect 4585 23420 4649 23424
rect 4585 23364 4589 23420
rect 4589 23364 4645 23420
rect 4645 23364 4649 23420
rect 4585 23360 4649 23364
rect 4665 23420 4729 23424
rect 4665 23364 4669 23420
rect 4669 23364 4725 23420
rect 4725 23364 4729 23420
rect 4665 23360 4729 23364
rect 11371 23420 11435 23424
rect 11371 23364 11375 23420
rect 11375 23364 11431 23420
rect 11431 23364 11435 23420
rect 11371 23360 11435 23364
rect 11451 23420 11515 23424
rect 11451 23364 11455 23420
rect 11455 23364 11511 23420
rect 11511 23364 11515 23420
rect 11451 23360 11515 23364
rect 11531 23420 11595 23424
rect 11531 23364 11535 23420
rect 11535 23364 11591 23420
rect 11591 23364 11595 23420
rect 11531 23360 11595 23364
rect 11611 23420 11675 23424
rect 11611 23364 11615 23420
rect 11615 23364 11671 23420
rect 11671 23364 11675 23420
rect 11611 23360 11675 23364
rect 18317 23420 18381 23424
rect 18317 23364 18321 23420
rect 18321 23364 18377 23420
rect 18377 23364 18381 23420
rect 18317 23360 18381 23364
rect 18397 23420 18461 23424
rect 18397 23364 18401 23420
rect 18401 23364 18457 23420
rect 18457 23364 18461 23420
rect 18397 23360 18461 23364
rect 18477 23420 18541 23424
rect 18477 23364 18481 23420
rect 18481 23364 18537 23420
rect 18537 23364 18541 23420
rect 18477 23360 18541 23364
rect 18557 23420 18621 23424
rect 18557 23364 18561 23420
rect 18561 23364 18617 23420
rect 18617 23364 18621 23420
rect 18557 23360 18621 23364
rect 25263 23420 25327 23424
rect 25263 23364 25267 23420
rect 25267 23364 25323 23420
rect 25323 23364 25327 23420
rect 25263 23360 25327 23364
rect 25343 23420 25407 23424
rect 25343 23364 25347 23420
rect 25347 23364 25403 23420
rect 25403 23364 25407 23420
rect 25343 23360 25407 23364
rect 25423 23420 25487 23424
rect 25423 23364 25427 23420
rect 25427 23364 25483 23420
rect 25483 23364 25487 23420
rect 25423 23360 25487 23364
rect 25503 23420 25567 23424
rect 25503 23364 25507 23420
rect 25507 23364 25563 23420
rect 25563 23364 25567 23420
rect 25503 23360 25567 23364
rect 7898 22876 7962 22880
rect 7898 22820 7902 22876
rect 7902 22820 7958 22876
rect 7958 22820 7962 22876
rect 7898 22816 7962 22820
rect 7978 22876 8042 22880
rect 7978 22820 7982 22876
rect 7982 22820 8038 22876
rect 8038 22820 8042 22876
rect 7978 22816 8042 22820
rect 8058 22876 8122 22880
rect 8058 22820 8062 22876
rect 8062 22820 8118 22876
rect 8118 22820 8122 22876
rect 8058 22816 8122 22820
rect 8138 22876 8202 22880
rect 8138 22820 8142 22876
rect 8142 22820 8198 22876
rect 8198 22820 8202 22876
rect 8138 22816 8202 22820
rect 14844 22876 14908 22880
rect 14844 22820 14848 22876
rect 14848 22820 14904 22876
rect 14904 22820 14908 22876
rect 14844 22816 14908 22820
rect 14924 22876 14988 22880
rect 14924 22820 14928 22876
rect 14928 22820 14984 22876
rect 14984 22820 14988 22876
rect 14924 22816 14988 22820
rect 15004 22876 15068 22880
rect 15004 22820 15008 22876
rect 15008 22820 15064 22876
rect 15064 22820 15068 22876
rect 15004 22816 15068 22820
rect 15084 22876 15148 22880
rect 15084 22820 15088 22876
rect 15088 22820 15144 22876
rect 15144 22820 15148 22876
rect 15084 22816 15148 22820
rect 21790 22876 21854 22880
rect 21790 22820 21794 22876
rect 21794 22820 21850 22876
rect 21850 22820 21854 22876
rect 21790 22816 21854 22820
rect 21870 22876 21934 22880
rect 21870 22820 21874 22876
rect 21874 22820 21930 22876
rect 21930 22820 21934 22876
rect 21870 22816 21934 22820
rect 21950 22876 22014 22880
rect 21950 22820 21954 22876
rect 21954 22820 22010 22876
rect 22010 22820 22014 22876
rect 21950 22816 22014 22820
rect 22030 22876 22094 22880
rect 22030 22820 22034 22876
rect 22034 22820 22090 22876
rect 22090 22820 22094 22876
rect 22030 22816 22094 22820
rect 28736 22876 28800 22880
rect 28736 22820 28740 22876
rect 28740 22820 28796 22876
rect 28796 22820 28800 22876
rect 28736 22816 28800 22820
rect 28816 22876 28880 22880
rect 28816 22820 28820 22876
rect 28820 22820 28876 22876
rect 28876 22820 28880 22876
rect 28816 22816 28880 22820
rect 28896 22876 28960 22880
rect 28896 22820 28900 22876
rect 28900 22820 28956 22876
rect 28956 22820 28960 22876
rect 28896 22816 28960 22820
rect 28976 22876 29040 22880
rect 28976 22820 28980 22876
rect 28980 22820 29036 22876
rect 29036 22820 29040 22876
rect 28976 22816 29040 22820
rect 4425 22332 4489 22336
rect 4425 22276 4429 22332
rect 4429 22276 4485 22332
rect 4485 22276 4489 22332
rect 4425 22272 4489 22276
rect 4505 22332 4569 22336
rect 4505 22276 4509 22332
rect 4509 22276 4565 22332
rect 4565 22276 4569 22332
rect 4505 22272 4569 22276
rect 4585 22332 4649 22336
rect 4585 22276 4589 22332
rect 4589 22276 4645 22332
rect 4645 22276 4649 22332
rect 4585 22272 4649 22276
rect 4665 22332 4729 22336
rect 4665 22276 4669 22332
rect 4669 22276 4725 22332
rect 4725 22276 4729 22332
rect 4665 22272 4729 22276
rect 11371 22332 11435 22336
rect 11371 22276 11375 22332
rect 11375 22276 11431 22332
rect 11431 22276 11435 22332
rect 11371 22272 11435 22276
rect 11451 22332 11515 22336
rect 11451 22276 11455 22332
rect 11455 22276 11511 22332
rect 11511 22276 11515 22332
rect 11451 22272 11515 22276
rect 11531 22332 11595 22336
rect 11531 22276 11535 22332
rect 11535 22276 11591 22332
rect 11591 22276 11595 22332
rect 11531 22272 11595 22276
rect 11611 22332 11675 22336
rect 11611 22276 11615 22332
rect 11615 22276 11671 22332
rect 11671 22276 11675 22332
rect 11611 22272 11675 22276
rect 18317 22332 18381 22336
rect 18317 22276 18321 22332
rect 18321 22276 18377 22332
rect 18377 22276 18381 22332
rect 18317 22272 18381 22276
rect 18397 22332 18461 22336
rect 18397 22276 18401 22332
rect 18401 22276 18457 22332
rect 18457 22276 18461 22332
rect 18397 22272 18461 22276
rect 18477 22332 18541 22336
rect 18477 22276 18481 22332
rect 18481 22276 18537 22332
rect 18537 22276 18541 22332
rect 18477 22272 18541 22276
rect 18557 22332 18621 22336
rect 18557 22276 18561 22332
rect 18561 22276 18617 22332
rect 18617 22276 18621 22332
rect 18557 22272 18621 22276
rect 25263 22332 25327 22336
rect 25263 22276 25267 22332
rect 25267 22276 25323 22332
rect 25323 22276 25327 22332
rect 25263 22272 25327 22276
rect 25343 22332 25407 22336
rect 25343 22276 25347 22332
rect 25347 22276 25403 22332
rect 25403 22276 25407 22332
rect 25343 22272 25407 22276
rect 25423 22332 25487 22336
rect 25423 22276 25427 22332
rect 25427 22276 25483 22332
rect 25483 22276 25487 22332
rect 25423 22272 25487 22276
rect 25503 22332 25567 22336
rect 25503 22276 25507 22332
rect 25507 22276 25563 22332
rect 25563 22276 25567 22332
rect 25503 22272 25567 22276
rect 7898 21788 7962 21792
rect 7898 21732 7902 21788
rect 7902 21732 7958 21788
rect 7958 21732 7962 21788
rect 7898 21728 7962 21732
rect 7978 21788 8042 21792
rect 7978 21732 7982 21788
rect 7982 21732 8038 21788
rect 8038 21732 8042 21788
rect 7978 21728 8042 21732
rect 8058 21788 8122 21792
rect 8058 21732 8062 21788
rect 8062 21732 8118 21788
rect 8118 21732 8122 21788
rect 8058 21728 8122 21732
rect 8138 21788 8202 21792
rect 8138 21732 8142 21788
rect 8142 21732 8198 21788
rect 8198 21732 8202 21788
rect 8138 21728 8202 21732
rect 14844 21788 14908 21792
rect 14844 21732 14848 21788
rect 14848 21732 14904 21788
rect 14904 21732 14908 21788
rect 14844 21728 14908 21732
rect 14924 21788 14988 21792
rect 14924 21732 14928 21788
rect 14928 21732 14984 21788
rect 14984 21732 14988 21788
rect 14924 21728 14988 21732
rect 15004 21788 15068 21792
rect 15004 21732 15008 21788
rect 15008 21732 15064 21788
rect 15064 21732 15068 21788
rect 15004 21728 15068 21732
rect 15084 21788 15148 21792
rect 15084 21732 15088 21788
rect 15088 21732 15144 21788
rect 15144 21732 15148 21788
rect 15084 21728 15148 21732
rect 21790 21788 21854 21792
rect 21790 21732 21794 21788
rect 21794 21732 21850 21788
rect 21850 21732 21854 21788
rect 21790 21728 21854 21732
rect 21870 21788 21934 21792
rect 21870 21732 21874 21788
rect 21874 21732 21930 21788
rect 21930 21732 21934 21788
rect 21870 21728 21934 21732
rect 21950 21788 22014 21792
rect 21950 21732 21954 21788
rect 21954 21732 22010 21788
rect 22010 21732 22014 21788
rect 21950 21728 22014 21732
rect 22030 21788 22094 21792
rect 22030 21732 22034 21788
rect 22034 21732 22090 21788
rect 22090 21732 22094 21788
rect 22030 21728 22094 21732
rect 28736 21788 28800 21792
rect 28736 21732 28740 21788
rect 28740 21732 28796 21788
rect 28796 21732 28800 21788
rect 28736 21728 28800 21732
rect 28816 21788 28880 21792
rect 28816 21732 28820 21788
rect 28820 21732 28876 21788
rect 28876 21732 28880 21788
rect 28816 21728 28880 21732
rect 28896 21788 28960 21792
rect 28896 21732 28900 21788
rect 28900 21732 28956 21788
rect 28956 21732 28960 21788
rect 28896 21728 28960 21732
rect 28976 21788 29040 21792
rect 28976 21732 28980 21788
rect 28980 21732 29036 21788
rect 29036 21732 29040 21788
rect 28976 21728 29040 21732
rect 4425 21244 4489 21248
rect 4425 21188 4429 21244
rect 4429 21188 4485 21244
rect 4485 21188 4489 21244
rect 4425 21184 4489 21188
rect 4505 21244 4569 21248
rect 4505 21188 4509 21244
rect 4509 21188 4565 21244
rect 4565 21188 4569 21244
rect 4505 21184 4569 21188
rect 4585 21244 4649 21248
rect 4585 21188 4589 21244
rect 4589 21188 4645 21244
rect 4645 21188 4649 21244
rect 4585 21184 4649 21188
rect 4665 21244 4729 21248
rect 4665 21188 4669 21244
rect 4669 21188 4725 21244
rect 4725 21188 4729 21244
rect 4665 21184 4729 21188
rect 11371 21244 11435 21248
rect 11371 21188 11375 21244
rect 11375 21188 11431 21244
rect 11431 21188 11435 21244
rect 11371 21184 11435 21188
rect 11451 21244 11515 21248
rect 11451 21188 11455 21244
rect 11455 21188 11511 21244
rect 11511 21188 11515 21244
rect 11451 21184 11515 21188
rect 11531 21244 11595 21248
rect 11531 21188 11535 21244
rect 11535 21188 11591 21244
rect 11591 21188 11595 21244
rect 11531 21184 11595 21188
rect 11611 21244 11675 21248
rect 11611 21188 11615 21244
rect 11615 21188 11671 21244
rect 11671 21188 11675 21244
rect 11611 21184 11675 21188
rect 18317 21244 18381 21248
rect 18317 21188 18321 21244
rect 18321 21188 18377 21244
rect 18377 21188 18381 21244
rect 18317 21184 18381 21188
rect 18397 21244 18461 21248
rect 18397 21188 18401 21244
rect 18401 21188 18457 21244
rect 18457 21188 18461 21244
rect 18397 21184 18461 21188
rect 18477 21244 18541 21248
rect 18477 21188 18481 21244
rect 18481 21188 18537 21244
rect 18537 21188 18541 21244
rect 18477 21184 18541 21188
rect 18557 21244 18621 21248
rect 18557 21188 18561 21244
rect 18561 21188 18617 21244
rect 18617 21188 18621 21244
rect 18557 21184 18621 21188
rect 25263 21244 25327 21248
rect 25263 21188 25267 21244
rect 25267 21188 25323 21244
rect 25323 21188 25327 21244
rect 25263 21184 25327 21188
rect 25343 21244 25407 21248
rect 25343 21188 25347 21244
rect 25347 21188 25403 21244
rect 25403 21188 25407 21244
rect 25343 21184 25407 21188
rect 25423 21244 25487 21248
rect 25423 21188 25427 21244
rect 25427 21188 25483 21244
rect 25483 21188 25487 21244
rect 25423 21184 25487 21188
rect 25503 21244 25567 21248
rect 25503 21188 25507 21244
rect 25507 21188 25563 21244
rect 25563 21188 25567 21244
rect 25503 21184 25567 21188
rect 7898 20700 7962 20704
rect 7898 20644 7902 20700
rect 7902 20644 7958 20700
rect 7958 20644 7962 20700
rect 7898 20640 7962 20644
rect 7978 20700 8042 20704
rect 7978 20644 7982 20700
rect 7982 20644 8038 20700
rect 8038 20644 8042 20700
rect 7978 20640 8042 20644
rect 8058 20700 8122 20704
rect 8058 20644 8062 20700
rect 8062 20644 8118 20700
rect 8118 20644 8122 20700
rect 8058 20640 8122 20644
rect 8138 20700 8202 20704
rect 8138 20644 8142 20700
rect 8142 20644 8198 20700
rect 8198 20644 8202 20700
rect 8138 20640 8202 20644
rect 14844 20700 14908 20704
rect 14844 20644 14848 20700
rect 14848 20644 14904 20700
rect 14904 20644 14908 20700
rect 14844 20640 14908 20644
rect 14924 20700 14988 20704
rect 14924 20644 14928 20700
rect 14928 20644 14984 20700
rect 14984 20644 14988 20700
rect 14924 20640 14988 20644
rect 15004 20700 15068 20704
rect 15004 20644 15008 20700
rect 15008 20644 15064 20700
rect 15064 20644 15068 20700
rect 15004 20640 15068 20644
rect 15084 20700 15148 20704
rect 15084 20644 15088 20700
rect 15088 20644 15144 20700
rect 15144 20644 15148 20700
rect 15084 20640 15148 20644
rect 21790 20700 21854 20704
rect 21790 20644 21794 20700
rect 21794 20644 21850 20700
rect 21850 20644 21854 20700
rect 21790 20640 21854 20644
rect 21870 20700 21934 20704
rect 21870 20644 21874 20700
rect 21874 20644 21930 20700
rect 21930 20644 21934 20700
rect 21870 20640 21934 20644
rect 21950 20700 22014 20704
rect 21950 20644 21954 20700
rect 21954 20644 22010 20700
rect 22010 20644 22014 20700
rect 21950 20640 22014 20644
rect 22030 20700 22094 20704
rect 22030 20644 22034 20700
rect 22034 20644 22090 20700
rect 22090 20644 22094 20700
rect 22030 20640 22094 20644
rect 28736 20700 28800 20704
rect 28736 20644 28740 20700
rect 28740 20644 28796 20700
rect 28796 20644 28800 20700
rect 28736 20640 28800 20644
rect 28816 20700 28880 20704
rect 28816 20644 28820 20700
rect 28820 20644 28876 20700
rect 28876 20644 28880 20700
rect 28816 20640 28880 20644
rect 28896 20700 28960 20704
rect 28896 20644 28900 20700
rect 28900 20644 28956 20700
rect 28956 20644 28960 20700
rect 28896 20640 28960 20644
rect 28976 20700 29040 20704
rect 28976 20644 28980 20700
rect 28980 20644 29036 20700
rect 29036 20644 29040 20700
rect 28976 20640 29040 20644
rect 4425 20156 4489 20160
rect 4425 20100 4429 20156
rect 4429 20100 4485 20156
rect 4485 20100 4489 20156
rect 4425 20096 4489 20100
rect 4505 20156 4569 20160
rect 4505 20100 4509 20156
rect 4509 20100 4565 20156
rect 4565 20100 4569 20156
rect 4505 20096 4569 20100
rect 4585 20156 4649 20160
rect 4585 20100 4589 20156
rect 4589 20100 4645 20156
rect 4645 20100 4649 20156
rect 4585 20096 4649 20100
rect 4665 20156 4729 20160
rect 4665 20100 4669 20156
rect 4669 20100 4725 20156
rect 4725 20100 4729 20156
rect 4665 20096 4729 20100
rect 11371 20156 11435 20160
rect 11371 20100 11375 20156
rect 11375 20100 11431 20156
rect 11431 20100 11435 20156
rect 11371 20096 11435 20100
rect 11451 20156 11515 20160
rect 11451 20100 11455 20156
rect 11455 20100 11511 20156
rect 11511 20100 11515 20156
rect 11451 20096 11515 20100
rect 11531 20156 11595 20160
rect 11531 20100 11535 20156
rect 11535 20100 11591 20156
rect 11591 20100 11595 20156
rect 11531 20096 11595 20100
rect 11611 20156 11675 20160
rect 11611 20100 11615 20156
rect 11615 20100 11671 20156
rect 11671 20100 11675 20156
rect 11611 20096 11675 20100
rect 18317 20156 18381 20160
rect 18317 20100 18321 20156
rect 18321 20100 18377 20156
rect 18377 20100 18381 20156
rect 18317 20096 18381 20100
rect 18397 20156 18461 20160
rect 18397 20100 18401 20156
rect 18401 20100 18457 20156
rect 18457 20100 18461 20156
rect 18397 20096 18461 20100
rect 18477 20156 18541 20160
rect 18477 20100 18481 20156
rect 18481 20100 18537 20156
rect 18537 20100 18541 20156
rect 18477 20096 18541 20100
rect 18557 20156 18621 20160
rect 18557 20100 18561 20156
rect 18561 20100 18617 20156
rect 18617 20100 18621 20156
rect 18557 20096 18621 20100
rect 25263 20156 25327 20160
rect 25263 20100 25267 20156
rect 25267 20100 25323 20156
rect 25323 20100 25327 20156
rect 25263 20096 25327 20100
rect 25343 20156 25407 20160
rect 25343 20100 25347 20156
rect 25347 20100 25403 20156
rect 25403 20100 25407 20156
rect 25343 20096 25407 20100
rect 25423 20156 25487 20160
rect 25423 20100 25427 20156
rect 25427 20100 25483 20156
rect 25483 20100 25487 20156
rect 25423 20096 25487 20100
rect 25503 20156 25567 20160
rect 25503 20100 25507 20156
rect 25507 20100 25563 20156
rect 25563 20100 25567 20156
rect 25503 20096 25567 20100
rect 7898 19612 7962 19616
rect 7898 19556 7902 19612
rect 7902 19556 7958 19612
rect 7958 19556 7962 19612
rect 7898 19552 7962 19556
rect 7978 19612 8042 19616
rect 7978 19556 7982 19612
rect 7982 19556 8038 19612
rect 8038 19556 8042 19612
rect 7978 19552 8042 19556
rect 8058 19612 8122 19616
rect 8058 19556 8062 19612
rect 8062 19556 8118 19612
rect 8118 19556 8122 19612
rect 8058 19552 8122 19556
rect 8138 19612 8202 19616
rect 8138 19556 8142 19612
rect 8142 19556 8198 19612
rect 8198 19556 8202 19612
rect 8138 19552 8202 19556
rect 14844 19612 14908 19616
rect 14844 19556 14848 19612
rect 14848 19556 14904 19612
rect 14904 19556 14908 19612
rect 14844 19552 14908 19556
rect 14924 19612 14988 19616
rect 14924 19556 14928 19612
rect 14928 19556 14984 19612
rect 14984 19556 14988 19612
rect 14924 19552 14988 19556
rect 15004 19612 15068 19616
rect 15004 19556 15008 19612
rect 15008 19556 15064 19612
rect 15064 19556 15068 19612
rect 15004 19552 15068 19556
rect 15084 19612 15148 19616
rect 15084 19556 15088 19612
rect 15088 19556 15144 19612
rect 15144 19556 15148 19612
rect 15084 19552 15148 19556
rect 21790 19612 21854 19616
rect 21790 19556 21794 19612
rect 21794 19556 21850 19612
rect 21850 19556 21854 19612
rect 21790 19552 21854 19556
rect 21870 19612 21934 19616
rect 21870 19556 21874 19612
rect 21874 19556 21930 19612
rect 21930 19556 21934 19612
rect 21870 19552 21934 19556
rect 21950 19612 22014 19616
rect 21950 19556 21954 19612
rect 21954 19556 22010 19612
rect 22010 19556 22014 19612
rect 21950 19552 22014 19556
rect 22030 19612 22094 19616
rect 22030 19556 22034 19612
rect 22034 19556 22090 19612
rect 22090 19556 22094 19612
rect 22030 19552 22094 19556
rect 28736 19612 28800 19616
rect 28736 19556 28740 19612
rect 28740 19556 28796 19612
rect 28796 19556 28800 19612
rect 28736 19552 28800 19556
rect 28816 19612 28880 19616
rect 28816 19556 28820 19612
rect 28820 19556 28876 19612
rect 28876 19556 28880 19612
rect 28816 19552 28880 19556
rect 28896 19612 28960 19616
rect 28896 19556 28900 19612
rect 28900 19556 28956 19612
rect 28956 19556 28960 19612
rect 28896 19552 28960 19556
rect 28976 19612 29040 19616
rect 28976 19556 28980 19612
rect 28980 19556 29036 19612
rect 29036 19556 29040 19612
rect 28976 19552 29040 19556
rect 4425 19068 4489 19072
rect 4425 19012 4429 19068
rect 4429 19012 4485 19068
rect 4485 19012 4489 19068
rect 4425 19008 4489 19012
rect 4505 19068 4569 19072
rect 4505 19012 4509 19068
rect 4509 19012 4565 19068
rect 4565 19012 4569 19068
rect 4505 19008 4569 19012
rect 4585 19068 4649 19072
rect 4585 19012 4589 19068
rect 4589 19012 4645 19068
rect 4645 19012 4649 19068
rect 4585 19008 4649 19012
rect 4665 19068 4729 19072
rect 4665 19012 4669 19068
rect 4669 19012 4725 19068
rect 4725 19012 4729 19068
rect 4665 19008 4729 19012
rect 11371 19068 11435 19072
rect 11371 19012 11375 19068
rect 11375 19012 11431 19068
rect 11431 19012 11435 19068
rect 11371 19008 11435 19012
rect 11451 19068 11515 19072
rect 11451 19012 11455 19068
rect 11455 19012 11511 19068
rect 11511 19012 11515 19068
rect 11451 19008 11515 19012
rect 11531 19068 11595 19072
rect 11531 19012 11535 19068
rect 11535 19012 11591 19068
rect 11591 19012 11595 19068
rect 11531 19008 11595 19012
rect 11611 19068 11675 19072
rect 11611 19012 11615 19068
rect 11615 19012 11671 19068
rect 11671 19012 11675 19068
rect 11611 19008 11675 19012
rect 18317 19068 18381 19072
rect 18317 19012 18321 19068
rect 18321 19012 18377 19068
rect 18377 19012 18381 19068
rect 18317 19008 18381 19012
rect 18397 19068 18461 19072
rect 18397 19012 18401 19068
rect 18401 19012 18457 19068
rect 18457 19012 18461 19068
rect 18397 19008 18461 19012
rect 18477 19068 18541 19072
rect 18477 19012 18481 19068
rect 18481 19012 18537 19068
rect 18537 19012 18541 19068
rect 18477 19008 18541 19012
rect 18557 19068 18621 19072
rect 18557 19012 18561 19068
rect 18561 19012 18617 19068
rect 18617 19012 18621 19068
rect 18557 19008 18621 19012
rect 25263 19068 25327 19072
rect 25263 19012 25267 19068
rect 25267 19012 25323 19068
rect 25323 19012 25327 19068
rect 25263 19008 25327 19012
rect 25343 19068 25407 19072
rect 25343 19012 25347 19068
rect 25347 19012 25403 19068
rect 25403 19012 25407 19068
rect 25343 19008 25407 19012
rect 25423 19068 25487 19072
rect 25423 19012 25427 19068
rect 25427 19012 25483 19068
rect 25483 19012 25487 19068
rect 25423 19008 25487 19012
rect 25503 19068 25567 19072
rect 25503 19012 25507 19068
rect 25507 19012 25563 19068
rect 25563 19012 25567 19068
rect 25503 19008 25567 19012
rect 7898 18524 7962 18528
rect 7898 18468 7902 18524
rect 7902 18468 7958 18524
rect 7958 18468 7962 18524
rect 7898 18464 7962 18468
rect 7978 18524 8042 18528
rect 7978 18468 7982 18524
rect 7982 18468 8038 18524
rect 8038 18468 8042 18524
rect 7978 18464 8042 18468
rect 8058 18524 8122 18528
rect 8058 18468 8062 18524
rect 8062 18468 8118 18524
rect 8118 18468 8122 18524
rect 8058 18464 8122 18468
rect 8138 18524 8202 18528
rect 8138 18468 8142 18524
rect 8142 18468 8198 18524
rect 8198 18468 8202 18524
rect 8138 18464 8202 18468
rect 14844 18524 14908 18528
rect 14844 18468 14848 18524
rect 14848 18468 14904 18524
rect 14904 18468 14908 18524
rect 14844 18464 14908 18468
rect 14924 18524 14988 18528
rect 14924 18468 14928 18524
rect 14928 18468 14984 18524
rect 14984 18468 14988 18524
rect 14924 18464 14988 18468
rect 15004 18524 15068 18528
rect 15004 18468 15008 18524
rect 15008 18468 15064 18524
rect 15064 18468 15068 18524
rect 15004 18464 15068 18468
rect 15084 18524 15148 18528
rect 15084 18468 15088 18524
rect 15088 18468 15144 18524
rect 15144 18468 15148 18524
rect 15084 18464 15148 18468
rect 21790 18524 21854 18528
rect 21790 18468 21794 18524
rect 21794 18468 21850 18524
rect 21850 18468 21854 18524
rect 21790 18464 21854 18468
rect 21870 18524 21934 18528
rect 21870 18468 21874 18524
rect 21874 18468 21930 18524
rect 21930 18468 21934 18524
rect 21870 18464 21934 18468
rect 21950 18524 22014 18528
rect 21950 18468 21954 18524
rect 21954 18468 22010 18524
rect 22010 18468 22014 18524
rect 21950 18464 22014 18468
rect 22030 18524 22094 18528
rect 22030 18468 22034 18524
rect 22034 18468 22090 18524
rect 22090 18468 22094 18524
rect 22030 18464 22094 18468
rect 28736 18524 28800 18528
rect 28736 18468 28740 18524
rect 28740 18468 28796 18524
rect 28796 18468 28800 18524
rect 28736 18464 28800 18468
rect 28816 18524 28880 18528
rect 28816 18468 28820 18524
rect 28820 18468 28876 18524
rect 28876 18468 28880 18524
rect 28816 18464 28880 18468
rect 28896 18524 28960 18528
rect 28896 18468 28900 18524
rect 28900 18468 28956 18524
rect 28956 18468 28960 18524
rect 28896 18464 28960 18468
rect 28976 18524 29040 18528
rect 28976 18468 28980 18524
rect 28980 18468 29036 18524
rect 29036 18468 29040 18524
rect 28976 18464 29040 18468
rect 4425 17980 4489 17984
rect 4425 17924 4429 17980
rect 4429 17924 4485 17980
rect 4485 17924 4489 17980
rect 4425 17920 4489 17924
rect 4505 17980 4569 17984
rect 4505 17924 4509 17980
rect 4509 17924 4565 17980
rect 4565 17924 4569 17980
rect 4505 17920 4569 17924
rect 4585 17980 4649 17984
rect 4585 17924 4589 17980
rect 4589 17924 4645 17980
rect 4645 17924 4649 17980
rect 4585 17920 4649 17924
rect 4665 17980 4729 17984
rect 4665 17924 4669 17980
rect 4669 17924 4725 17980
rect 4725 17924 4729 17980
rect 4665 17920 4729 17924
rect 11371 17980 11435 17984
rect 11371 17924 11375 17980
rect 11375 17924 11431 17980
rect 11431 17924 11435 17980
rect 11371 17920 11435 17924
rect 11451 17980 11515 17984
rect 11451 17924 11455 17980
rect 11455 17924 11511 17980
rect 11511 17924 11515 17980
rect 11451 17920 11515 17924
rect 11531 17980 11595 17984
rect 11531 17924 11535 17980
rect 11535 17924 11591 17980
rect 11591 17924 11595 17980
rect 11531 17920 11595 17924
rect 11611 17980 11675 17984
rect 11611 17924 11615 17980
rect 11615 17924 11671 17980
rect 11671 17924 11675 17980
rect 11611 17920 11675 17924
rect 18317 17980 18381 17984
rect 18317 17924 18321 17980
rect 18321 17924 18377 17980
rect 18377 17924 18381 17980
rect 18317 17920 18381 17924
rect 18397 17980 18461 17984
rect 18397 17924 18401 17980
rect 18401 17924 18457 17980
rect 18457 17924 18461 17980
rect 18397 17920 18461 17924
rect 18477 17980 18541 17984
rect 18477 17924 18481 17980
rect 18481 17924 18537 17980
rect 18537 17924 18541 17980
rect 18477 17920 18541 17924
rect 18557 17980 18621 17984
rect 18557 17924 18561 17980
rect 18561 17924 18617 17980
rect 18617 17924 18621 17980
rect 18557 17920 18621 17924
rect 25263 17980 25327 17984
rect 25263 17924 25267 17980
rect 25267 17924 25323 17980
rect 25323 17924 25327 17980
rect 25263 17920 25327 17924
rect 25343 17980 25407 17984
rect 25343 17924 25347 17980
rect 25347 17924 25403 17980
rect 25403 17924 25407 17980
rect 25343 17920 25407 17924
rect 25423 17980 25487 17984
rect 25423 17924 25427 17980
rect 25427 17924 25483 17980
rect 25483 17924 25487 17980
rect 25423 17920 25487 17924
rect 25503 17980 25567 17984
rect 25503 17924 25507 17980
rect 25507 17924 25563 17980
rect 25563 17924 25567 17980
rect 25503 17920 25567 17924
rect 7898 17436 7962 17440
rect 7898 17380 7902 17436
rect 7902 17380 7958 17436
rect 7958 17380 7962 17436
rect 7898 17376 7962 17380
rect 7978 17436 8042 17440
rect 7978 17380 7982 17436
rect 7982 17380 8038 17436
rect 8038 17380 8042 17436
rect 7978 17376 8042 17380
rect 8058 17436 8122 17440
rect 8058 17380 8062 17436
rect 8062 17380 8118 17436
rect 8118 17380 8122 17436
rect 8058 17376 8122 17380
rect 8138 17436 8202 17440
rect 8138 17380 8142 17436
rect 8142 17380 8198 17436
rect 8198 17380 8202 17436
rect 8138 17376 8202 17380
rect 14844 17436 14908 17440
rect 14844 17380 14848 17436
rect 14848 17380 14904 17436
rect 14904 17380 14908 17436
rect 14844 17376 14908 17380
rect 14924 17436 14988 17440
rect 14924 17380 14928 17436
rect 14928 17380 14984 17436
rect 14984 17380 14988 17436
rect 14924 17376 14988 17380
rect 15004 17436 15068 17440
rect 15004 17380 15008 17436
rect 15008 17380 15064 17436
rect 15064 17380 15068 17436
rect 15004 17376 15068 17380
rect 15084 17436 15148 17440
rect 15084 17380 15088 17436
rect 15088 17380 15144 17436
rect 15144 17380 15148 17436
rect 15084 17376 15148 17380
rect 21790 17436 21854 17440
rect 21790 17380 21794 17436
rect 21794 17380 21850 17436
rect 21850 17380 21854 17436
rect 21790 17376 21854 17380
rect 21870 17436 21934 17440
rect 21870 17380 21874 17436
rect 21874 17380 21930 17436
rect 21930 17380 21934 17436
rect 21870 17376 21934 17380
rect 21950 17436 22014 17440
rect 21950 17380 21954 17436
rect 21954 17380 22010 17436
rect 22010 17380 22014 17436
rect 21950 17376 22014 17380
rect 22030 17436 22094 17440
rect 22030 17380 22034 17436
rect 22034 17380 22090 17436
rect 22090 17380 22094 17436
rect 22030 17376 22094 17380
rect 28736 17436 28800 17440
rect 28736 17380 28740 17436
rect 28740 17380 28796 17436
rect 28796 17380 28800 17436
rect 28736 17376 28800 17380
rect 28816 17436 28880 17440
rect 28816 17380 28820 17436
rect 28820 17380 28876 17436
rect 28876 17380 28880 17436
rect 28816 17376 28880 17380
rect 28896 17436 28960 17440
rect 28896 17380 28900 17436
rect 28900 17380 28956 17436
rect 28956 17380 28960 17436
rect 28896 17376 28960 17380
rect 28976 17436 29040 17440
rect 28976 17380 28980 17436
rect 28980 17380 29036 17436
rect 29036 17380 29040 17436
rect 28976 17376 29040 17380
rect 4425 16892 4489 16896
rect 4425 16836 4429 16892
rect 4429 16836 4485 16892
rect 4485 16836 4489 16892
rect 4425 16832 4489 16836
rect 4505 16892 4569 16896
rect 4505 16836 4509 16892
rect 4509 16836 4565 16892
rect 4565 16836 4569 16892
rect 4505 16832 4569 16836
rect 4585 16892 4649 16896
rect 4585 16836 4589 16892
rect 4589 16836 4645 16892
rect 4645 16836 4649 16892
rect 4585 16832 4649 16836
rect 4665 16892 4729 16896
rect 4665 16836 4669 16892
rect 4669 16836 4725 16892
rect 4725 16836 4729 16892
rect 4665 16832 4729 16836
rect 11371 16892 11435 16896
rect 11371 16836 11375 16892
rect 11375 16836 11431 16892
rect 11431 16836 11435 16892
rect 11371 16832 11435 16836
rect 11451 16892 11515 16896
rect 11451 16836 11455 16892
rect 11455 16836 11511 16892
rect 11511 16836 11515 16892
rect 11451 16832 11515 16836
rect 11531 16892 11595 16896
rect 11531 16836 11535 16892
rect 11535 16836 11591 16892
rect 11591 16836 11595 16892
rect 11531 16832 11595 16836
rect 11611 16892 11675 16896
rect 11611 16836 11615 16892
rect 11615 16836 11671 16892
rect 11671 16836 11675 16892
rect 11611 16832 11675 16836
rect 18317 16892 18381 16896
rect 18317 16836 18321 16892
rect 18321 16836 18377 16892
rect 18377 16836 18381 16892
rect 18317 16832 18381 16836
rect 18397 16892 18461 16896
rect 18397 16836 18401 16892
rect 18401 16836 18457 16892
rect 18457 16836 18461 16892
rect 18397 16832 18461 16836
rect 18477 16892 18541 16896
rect 18477 16836 18481 16892
rect 18481 16836 18537 16892
rect 18537 16836 18541 16892
rect 18477 16832 18541 16836
rect 18557 16892 18621 16896
rect 18557 16836 18561 16892
rect 18561 16836 18617 16892
rect 18617 16836 18621 16892
rect 18557 16832 18621 16836
rect 25263 16892 25327 16896
rect 25263 16836 25267 16892
rect 25267 16836 25323 16892
rect 25323 16836 25327 16892
rect 25263 16832 25327 16836
rect 25343 16892 25407 16896
rect 25343 16836 25347 16892
rect 25347 16836 25403 16892
rect 25403 16836 25407 16892
rect 25343 16832 25407 16836
rect 25423 16892 25487 16896
rect 25423 16836 25427 16892
rect 25427 16836 25483 16892
rect 25483 16836 25487 16892
rect 25423 16832 25487 16836
rect 25503 16892 25567 16896
rect 25503 16836 25507 16892
rect 25507 16836 25563 16892
rect 25563 16836 25567 16892
rect 25503 16832 25567 16836
rect 7898 16348 7962 16352
rect 7898 16292 7902 16348
rect 7902 16292 7958 16348
rect 7958 16292 7962 16348
rect 7898 16288 7962 16292
rect 7978 16348 8042 16352
rect 7978 16292 7982 16348
rect 7982 16292 8038 16348
rect 8038 16292 8042 16348
rect 7978 16288 8042 16292
rect 8058 16348 8122 16352
rect 8058 16292 8062 16348
rect 8062 16292 8118 16348
rect 8118 16292 8122 16348
rect 8058 16288 8122 16292
rect 8138 16348 8202 16352
rect 8138 16292 8142 16348
rect 8142 16292 8198 16348
rect 8198 16292 8202 16348
rect 8138 16288 8202 16292
rect 14844 16348 14908 16352
rect 14844 16292 14848 16348
rect 14848 16292 14904 16348
rect 14904 16292 14908 16348
rect 14844 16288 14908 16292
rect 14924 16348 14988 16352
rect 14924 16292 14928 16348
rect 14928 16292 14984 16348
rect 14984 16292 14988 16348
rect 14924 16288 14988 16292
rect 15004 16348 15068 16352
rect 15004 16292 15008 16348
rect 15008 16292 15064 16348
rect 15064 16292 15068 16348
rect 15004 16288 15068 16292
rect 15084 16348 15148 16352
rect 15084 16292 15088 16348
rect 15088 16292 15144 16348
rect 15144 16292 15148 16348
rect 15084 16288 15148 16292
rect 21790 16348 21854 16352
rect 21790 16292 21794 16348
rect 21794 16292 21850 16348
rect 21850 16292 21854 16348
rect 21790 16288 21854 16292
rect 21870 16348 21934 16352
rect 21870 16292 21874 16348
rect 21874 16292 21930 16348
rect 21930 16292 21934 16348
rect 21870 16288 21934 16292
rect 21950 16348 22014 16352
rect 21950 16292 21954 16348
rect 21954 16292 22010 16348
rect 22010 16292 22014 16348
rect 21950 16288 22014 16292
rect 22030 16348 22094 16352
rect 22030 16292 22034 16348
rect 22034 16292 22090 16348
rect 22090 16292 22094 16348
rect 22030 16288 22094 16292
rect 28736 16348 28800 16352
rect 28736 16292 28740 16348
rect 28740 16292 28796 16348
rect 28796 16292 28800 16348
rect 28736 16288 28800 16292
rect 28816 16348 28880 16352
rect 28816 16292 28820 16348
rect 28820 16292 28876 16348
rect 28876 16292 28880 16348
rect 28816 16288 28880 16292
rect 28896 16348 28960 16352
rect 28896 16292 28900 16348
rect 28900 16292 28956 16348
rect 28956 16292 28960 16348
rect 28896 16288 28960 16292
rect 28976 16348 29040 16352
rect 28976 16292 28980 16348
rect 28980 16292 29036 16348
rect 29036 16292 29040 16348
rect 28976 16288 29040 16292
rect 4425 15804 4489 15808
rect 4425 15748 4429 15804
rect 4429 15748 4485 15804
rect 4485 15748 4489 15804
rect 4425 15744 4489 15748
rect 4505 15804 4569 15808
rect 4505 15748 4509 15804
rect 4509 15748 4565 15804
rect 4565 15748 4569 15804
rect 4505 15744 4569 15748
rect 4585 15804 4649 15808
rect 4585 15748 4589 15804
rect 4589 15748 4645 15804
rect 4645 15748 4649 15804
rect 4585 15744 4649 15748
rect 4665 15804 4729 15808
rect 4665 15748 4669 15804
rect 4669 15748 4725 15804
rect 4725 15748 4729 15804
rect 4665 15744 4729 15748
rect 11371 15804 11435 15808
rect 11371 15748 11375 15804
rect 11375 15748 11431 15804
rect 11431 15748 11435 15804
rect 11371 15744 11435 15748
rect 11451 15804 11515 15808
rect 11451 15748 11455 15804
rect 11455 15748 11511 15804
rect 11511 15748 11515 15804
rect 11451 15744 11515 15748
rect 11531 15804 11595 15808
rect 11531 15748 11535 15804
rect 11535 15748 11591 15804
rect 11591 15748 11595 15804
rect 11531 15744 11595 15748
rect 11611 15804 11675 15808
rect 11611 15748 11615 15804
rect 11615 15748 11671 15804
rect 11671 15748 11675 15804
rect 11611 15744 11675 15748
rect 18317 15804 18381 15808
rect 18317 15748 18321 15804
rect 18321 15748 18377 15804
rect 18377 15748 18381 15804
rect 18317 15744 18381 15748
rect 18397 15804 18461 15808
rect 18397 15748 18401 15804
rect 18401 15748 18457 15804
rect 18457 15748 18461 15804
rect 18397 15744 18461 15748
rect 18477 15804 18541 15808
rect 18477 15748 18481 15804
rect 18481 15748 18537 15804
rect 18537 15748 18541 15804
rect 18477 15744 18541 15748
rect 18557 15804 18621 15808
rect 18557 15748 18561 15804
rect 18561 15748 18617 15804
rect 18617 15748 18621 15804
rect 18557 15744 18621 15748
rect 25263 15804 25327 15808
rect 25263 15748 25267 15804
rect 25267 15748 25323 15804
rect 25323 15748 25327 15804
rect 25263 15744 25327 15748
rect 25343 15804 25407 15808
rect 25343 15748 25347 15804
rect 25347 15748 25403 15804
rect 25403 15748 25407 15804
rect 25343 15744 25407 15748
rect 25423 15804 25487 15808
rect 25423 15748 25427 15804
rect 25427 15748 25483 15804
rect 25483 15748 25487 15804
rect 25423 15744 25487 15748
rect 25503 15804 25567 15808
rect 25503 15748 25507 15804
rect 25507 15748 25563 15804
rect 25563 15748 25567 15804
rect 25503 15744 25567 15748
rect 7898 15260 7962 15264
rect 7898 15204 7902 15260
rect 7902 15204 7958 15260
rect 7958 15204 7962 15260
rect 7898 15200 7962 15204
rect 7978 15260 8042 15264
rect 7978 15204 7982 15260
rect 7982 15204 8038 15260
rect 8038 15204 8042 15260
rect 7978 15200 8042 15204
rect 8058 15260 8122 15264
rect 8058 15204 8062 15260
rect 8062 15204 8118 15260
rect 8118 15204 8122 15260
rect 8058 15200 8122 15204
rect 8138 15260 8202 15264
rect 8138 15204 8142 15260
rect 8142 15204 8198 15260
rect 8198 15204 8202 15260
rect 8138 15200 8202 15204
rect 14844 15260 14908 15264
rect 14844 15204 14848 15260
rect 14848 15204 14904 15260
rect 14904 15204 14908 15260
rect 14844 15200 14908 15204
rect 14924 15260 14988 15264
rect 14924 15204 14928 15260
rect 14928 15204 14984 15260
rect 14984 15204 14988 15260
rect 14924 15200 14988 15204
rect 15004 15260 15068 15264
rect 15004 15204 15008 15260
rect 15008 15204 15064 15260
rect 15064 15204 15068 15260
rect 15004 15200 15068 15204
rect 15084 15260 15148 15264
rect 15084 15204 15088 15260
rect 15088 15204 15144 15260
rect 15144 15204 15148 15260
rect 15084 15200 15148 15204
rect 21790 15260 21854 15264
rect 21790 15204 21794 15260
rect 21794 15204 21850 15260
rect 21850 15204 21854 15260
rect 21790 15200 21854 15204
rect 21870 15260 21934 15264
rect 21870 15204 21874 15260
rect 21874 15204 21930 15260
rect 21930 15204 21934 15260
rect 21870 15200 21934 15204
rect 21950 15260 22014 15264
rect 21950 15204 21954 15260
rect 21954 15204 22010 15260
rect 22010 15204 22014 15260
rect 21950 15200 22014 15204
rect 22030 15260 22094 15264
rect 22030 15204 22034 15260
rect 22034 15204 22090 15260
rect 22090 15204 22094 15260
rect 22030 15200 22094 15204
rect 28736 15260 28800 15264
rect 28736 15204 28740 15260
rect 28740 15204 28796 15260
rect 28796 15204 28800 15260
rect 28736 15200 28800 15204
rect 28816 15260 28880 15264
rect 28816 15204 28820 15260
rect 28820 15204 28876 15260
rect 28876 15204 28880 15260
rect 28816 15200 28880 15204
rect 28896 15260 28960 15264
rect 28896 15204 28900 15260
rect 28900 15204 28956 15260
rect 28956 15204 28960 15260
rect 28896 15200 28960 15204
rect 28976 15260 29040 15264
rect 28976 15204 28980 15260
rect 28980 15204 29036 15260
rect 29036 15204 29040 15260
rect 28976 15200 29040 15204
rect 4425 14716 4489 14720
rect 4425 14660 4429 14716
rect 4429 14660 4485 14716
rect 4485 14660 4489 14716
rect 4425 14656 4489 14660
rect 4505 14716 4569 14720
rect 4505 14660 4509 14716
rect 4509 14660 4565 14716
rect 4565 14660 4569 14716
rect 4505 14656 4569 14660
rect 4585 14716 4649 14720
rect 4585 14660 4589 14716
rect 4589 14660 4645 14716
rect 4645 14660 4649 14716
rect 4585 14656 4649 14660
rect 4665 14716 4729 14720
rect 4665 14660 4669 14716
rect 4669 14660 4725 14716
rect 4725 14660 4729 14716
rect 4665 14656 4729 14660
rect 11371 14716 11435 14720
rect 11371 14660 11375 14716
rect 11375 14660 11431 14716
rect 11431 14660 11435 14716
rect 11371 14656 11435 14660
rect 11451 14716 11515 14720
rect 11451 14660 11455 14716
rect 11455 14660 11511 14716
rect 11511 14660 11515 14716
rect 11451 14656 11515 14660
rect 11531 14716 11595 14720
rect 11531 14660 11535 14716
rect 11535 14660 11591 14716
rect 11591 14660 11595 14716
rect 11531 14656 11595 14660
rect 11611 14716 11675 14720
rect 11611 14660 11615 14716
rect 11615 14660 11671 14716
rect 11671 14660 11675 14716
rect 11611 14656 11675 14660
rect 18317 14716 18381 14720
rect 18317 14660 18321 14716
rect 18321 14660 18377 14716
rect 18377 14660 18381 14716
rect 18317 14656 18381 14660
rect 18397 14716 18461 14720
rect 18397 14660 18401 14716
rect 18401 14660 18457 14716
rect 18457 14660 18461 14716
rect 18397 14656 18461 14660
rect 18477 14716 18541 14720
rect 18477 14660 18481 14716
rect 18481 14660 18537 14716
rect 18537 14660 18541 14716
rect 18477 14656 18541 14660
rect 18557 14716 18621 14720
rect 18557 14660 18561 14716
rect 18561 14660 18617 14716
rect 18617 14660 18621 14716
rect 18557 14656 18621 14660
rect 25263 14716 25327 14720
rect 25263 14660 25267 14716
rect 25267 14660 25323 14716
rect 25323 14660 25327 14716
rect 25263 14656 25327 14660
rect 25343 14716 25407 14720
rect 25343 14660 25347 14716
rect 25347 14660 25403 14716
rect 25403 14660 25407 14716
rect 25343 14656 25407 14660
rect 25423 14716 25487 14720
rect 25423 14660 25427 14716
rect 25427 14660 25483 14716
rect 25483 14660 25487 14716
rect 25423 14656 25487 14660
rect 25503 14716 25567 14720
rect 25503 14660 25507 14716
rect 25507 14660 25563 14716
rect 25563 14660 25567 14716
rect 25503 14656 25567 14660
rect 7898 14172 7962 14176
rect 7898 14116 7902 14172
rect 7902 14116 7958 14172
rect 7958 14116 7962 14172
rect 7898 14112 7962 14116
rect 7978 14172 8042 14176
rect 7978 14116 7982 14172
rect 7982 14116 8038 14172
rect 8038 14116 8042 14172
rect 7978 14112 8042 14116
rect 8058 14172 8122 14176
rect 8058 14116 8062 14172
rect 8062 14116 8118 14172
rect 8118 14116 8122 14172
rect 8058 14112 8122 14116
rect 8138 14172 8202 14176
rect 8138 14116 8142 14172
rect 8142 14116 8198 14172
rect 8198 14116 8202 14172
rect 8138 14112 8202 14116
rect 14844 14172 14908 14176
rect 14844 14116 14848 14172
rect 14848 14116 14904 14172
rect 14904 14116 14908 14172
rect 14844 14112 14908 14116
rect 14924 14172 14988 14176
rect 14924 14116 14928 14172
rect 14928 14116 14984 14172
rect 14984 14116 14988 14172
rect 14924 14112 14988 14116
rect 15004 14172 15068 14176
rect 15004 14116 15008 14172
rect 15008 14116 15064 14172
rect 15064 14116 15068 14172
rect 15004 14112 15068 14116
rect 15084 14172 15148 14176
rect 15084 14116 15088 14172
rect 15088 14116 15144 14172
rect 15144 14116 15148 14172
rect 15084 14112 15148 14116
rect 21790 14172 21854 14176
rect 21790 14116 21794 14172
rect 21794 14116 21850 14172
rect 21850 14116 21854 14172
rect 21790 14112 21854 14116
rect 21870 14172 21934 14176
rect 21870 14116 21874 14172
rect 21874 14116 21930 14172
rect 21930 14116 21934 14172
rect 21870 14112 21934 14116
rect 21950 14172 22014 14176
rect 21950 14116 21954 14172
rect 21954 14116 22010 14172
rect 22010 14116 22014 14172
rect 21950 14112 22014 14116
rect 22030 14172 22094 14176
rect 22030 14116 22034 14172
rect 22034 14116 22090 14172
rect 22090 14116 22094 14172
rect 22030 14112 22094 14116
rect 28736 14172 28800 14176
rect 28736 14116 28740 14172
rect 28740 14116 28796 14172
rect 28796 14116 28800 14172
rect 28736 14112 28800 14116
rect 28816 14172 28880 14176
rect 28816 14116 28820 14172
rect 28820 14116 28876 14172
rect 28876 14116 28880 14172
rect 28816 14112 28880 14116
rect 28896 14172 28960 14176
rect 28896 14116 28900 14172
rect 28900 14116 28956 14172
rect 28956 14116 28960 14172
rect 28896 14112 28960 14116
rect 28976 14172 29040 14176
rect 28976 14116 28980 14172
rect 28980 14116 29036 14172
rect 29036 14116 29040 14172
rect 28976 14112 29040 14116
rect 4425 13628 4489 13632
rect 4425 13572 4429 13628
rect 4429 13572 4485 13628
rect 4485 13572 4489 13628
rect 4425 13568 4489 13572
rect 4505 13628 4569 13632
rect 4505 13572 4509 13628
rect 4509 13572 4565 13628
rect 4565 13572 4569 13628
rect 4505 13568 4569 13572
rect 4585 13628 4649 13632
rect 4585 13572 4589 13628
rect 4589 13572 4645 13628
rect 4645 13572 4649 13628
rect 4585 13568 4649 13572
rect 4665 13628 4729 13632
rect 4665 13572 4669 13628
rect 4669 13572 4725 13628
rect 4725 13572 4729 13628
rect 4665 13568 4729 13572
rect 11371 13628 11435 13632
rect 11371 13572 11375 13628
rect 11375 13572 11431 13628
rect 11431 13572 11435 13628
rect 11371 13568 11435 13572
rect 11451 13628 11515 13632
rect 11451 13572 11455 13628
rect 11455 13572 11511 13628
rect 11511 13572 11515 13628
rect 11451 13568 11515 13572
rect 11531 13628 11595 13632
rect 11531 13572 11535 13628
rect 11535 13572 11591 13628
rect 11591 13572 11595 13628
rect 11531 13568 11595 13572
rect 11611 13628 11675 13632
rect 11611 13572 11615 13628
rect 11615 13572 11671 13628
rect 11671 13572 11675 13628
rect 11611 13568 11675 13572
rect 18317 13628 18381 13632
rect 18317 13572 18321 13628
rect 18321 13572 18377 13628
rect 18377 13572 18381 13628
rect 18317 13568 18381 13572
rect 18397 13628 18461 13632
rect 18397 13572 18401 13628
rect 18401 13572 18457 13628
rect 18457 13572 18461 13628
rect 18397 13568 18461 13572
rect 18477 13628 18541 13632
rect 18477 13572 18481 13628
rect 18481 13572 18537 13628
rect 18537 13572 18541 13628
rect 18477 13568 18541 13572
rect 18557 13628 18621 13632
rect 18557 13572 18561 13628
rect 18561 13572 18617 13628
rect 18617 13572 18621 13628
rect 18557 13568 18621 13572
rect 25263 13628 25327 13632
rect 25263 13572 25267 13628
rect 25267 13572 25323 13628
rect 25323 13572 25327 13628
rect 25263 13568 25327 13572
rect 25343 13628 25407 13632
rect 25343 13572 25347 13628
rect 25347 13572 25403 13628
rect 25403 13572 25407 13628
rect 25343 13568 25407 13572
rect 25423 13628 25487 13632
rect 25423 13572 25427 13628
rect 25427 13572 25483 13628
rect 25483 13572 25487 13628
rect 25423 13568 25487 13572
rect 25503 13628 25567 13632
rect 25503 13572 25507 13628
rect 25507 13572 25563 13628
rect 25563 13572 25567 13628
rect 25503 13568 25567 13572
rect 7898 13084 7962 13088
rect 7898 13028 7902 13084
rect 7902 13028 7958 13084
rect 7958 13028 7962 13084
rect 7898 13024 7962 13028
rect 7978 13084 8042 13088
rect 7978 13028 7982 13084
rect 7982 13028 8038 13084
rect 8038 13028 8042 13084
rect 7978 13024 8042 13028
rect 8058 13084 8122 13088
rect 8058 13028 8062 13084
rect 8062 13028 8118 13084
rect 8118 13028 8122 13084
rect 8058 13024 8122 13028
rect 8138 13084 8202 13088
rect 8138 13028 8142 13084
rect 8142 13028 8198 13084
rect 8198 13028 8202 13084
rect 8138 13024 8202 13028
rect 14844 13084 14908 13088
rect 14844 13028 14848 13084
rect 14848 13028 14904 13084
rect 14904 13028 14908 13084
rect 14844 13024 14908 13028
rect 14924 13084 14988 13088
rect 14924 13028 14928 13084
rect 14928 13028 14984 13084
rect 14984 13028 14988 13084
rect 14924 13024 14988 13028
rect 15004 13084 15068 13088
rect 15004 13028 15008 13084
rect 15008 13028 15064 13084
rect 15064 13028 15068 13084
rect 15004 13024 15068 13028
rect 15084 13084 15148 13088
rect 15084 13028 15088 13084
rect 15088 13028 15144 13084
rect 15144 13028 15148 13084
rect 15084 13024 15148 13028
rect 21790 13084 21854 13088
rect 21790 13028 21794 13084
rect 21794 13028 21850 13084
rect 21850 13028 21854 13084
rect 21790 13024 21854 13028
rect 21870 13084 21934 13088
rect 21870 13028 21874 13084
rect 21874 13028 21930 13084
rect 21930 13028 21934 13084
rect 21870 13024 21934 13028
rect 21950 13084 22014 13088
rect 21950 13028 21954 13084
rect 21954 13028 22010 13084
rect 22010 13028 22014 13084
rect 21950 13024 22014 13028
rect 22030 13084 22094 13088
rect 22030 13028 22034 13084
rect 22034 13028 22090 13084
rect 22090 13028 22094 13084
rect 22030 13024 22094 13028
rect 28736 13084 28800 13088
rect 28736 13028 28740 13084
rect 28740 13028 28796 13084
rect 28796 13028 28800 13084
rect 28736 13024 28800 13028
rect 28816 13084 28880 13088
rect 28816 13028 28820 13084
rect 28820 13028 28876 13084
rect 28876 13028 28880 13084
rect 28816 13024 28880 13028
rect 28896 13084 28960 13088
rect 28896 13028 28900 13084
rect 28900 13028 28956 13084
rect 28956 13028 28960 13084
rect 28896 13024 28960 13028
rect 28976 13084 29040 13088
rect 28976 13028 28980 13084
rect 28980 13028 29036 13084
rect 29036 13028 29040 13084
rect 28976 13024 29040 13028
rect 4425 12540 4489 12544
rect 4425 12484 4429 12540
rect 4429 12484 4485 12540
rect 4485 12484 4489 12540
rect 4425 12480 4489 12484
rect 4505 12540 4569 12544
rect 4505 12484 4509 12540
rect 4509 12484 4565 12540
rect 4565 12484 4569 12540
rect 4505 12480 4569 12484
rect 4585 12540 4649 12544
rect 4585 12484 4589 12540
rect 4589 12484 4645 12540
rect 4645 12484 4649 12540
rect 4585 12480 4649 12484
rect 4665 12540 4729 12544
rect 4665 12484 4669 12540
rect 4669 12484 4725 12540
rect 4725 12484 4729 12540
rect 4665 12480 4729 12484
rect 11371 12540 11435 12544
rect 11371 12484 11375 12540
rect 11375 12484 11431 12540
rect 11431 12484 11435 12540
rect 11371 12480 11435 12484
rect 11451 12540 11515 12544
rect 11451 12484 11455 12540
rect 11455 12484 11511 12540
rect 11511 12484 11515 12540
rect 11451 12480 11515 12484
rect 11531 12540 11595 12544
rect 11531 12484 11535 12540
rect 11535 12484 11591 12540
rect 11591 12484 11595 12540
rect 11531 12480 11595 12484
rect 11611 12540 11675 12544
rect 11611 12484 11615 12540
rect 11615 12484 11671 12540
rect 11671 12484 11675 12540
rect 11611 12480 11675 12484
rect 18317 12540 18381 12544
rect 18317 12484 18321 12540
rect 18321 12484 18377 12540
rect 18377 12484 18381 12540
rect 18317 12480 18381 12484
rect 18397 12540 18461 12544
rect 18397 12484 18401 12540
rect 18401 12484 18457 12540
rect 18457 12484 18461 12540
rect 18397 12480 18461 12484
rect 18477 12540 18541 12544
rect 18477 12484 18481 12540
rect 18481 12484 18537 12540
rect 18537 12484 18541 12540
rect 18477 12480 18541 12484
rect 18557 12540 18621 12544
rect 18557 12484 18561 12540
rect 18561 12484 18617 12540
rect 18617 12484 18621 12540
rect 18557 12480 18621 12484
rect 25263 12540 25327 12544
rect 25263 12484 25267 12540
rect 25267 12484 25323 12540
rect 25323 12484 25327 12540
rect 25263 12480 25327 12484
rect 25343 12540 25407 12544
rect 25343 12484 25347 12540
rect 25347 12484 25403 12540
rect 25403 12484 25407 12540
rect 25343 12480 25407 12484
rect 25423 12540 25487 12544
rect 25423 12484 25427 12540
rect 25427 12484 25483 12540
rect 25483 12484 25487 12540
rect 25423 12480 25487 12484
rect 25503 12540 25567 12544
rect 25503 12484 25507 12540
rect 25507 12484 25563 12540
rect 25563 12484 25567 12540
rect 25503 12480 25567 12484
rect 7898 11996 7962 12000
rect 7898 11940 7902 11996
rect 7902 11940 7958 11996
rect 7958 11940 7962 11996
rect 7898 11936 7962 11940
rect 7978 11996 8042 12000
rect 7978 11940 7982 11996
rect 7982 11940 8038 11996
rect 8038 11940 8042 11996
rect 7978 11936 8042 11940
rect 8058 11996 8122 12000
rect 8058 11940 8062 11996
rect 8062 11940 8118 11996
rect 8118 11940 8122 11996
rect 8058 11936 8122 11940
rect 8138 11996 8202 12000
rect 8138 11940 8142 11996
rect 8142 11940 8198 11996
rect 8198 11940 8202 11996
rect 8138 11936 8202 11940
rect 14844 11996 14908 12000
rect 14844 11940 14848 11996
rect 14848 11940 14904 11996
rect 14904 11940 14908 11996
rect 14844 11936 14908 11940
rect 14924 11996 14988 12000
rect 14924 11940 14928 11996
rect 14928 11940 14984 11996
rect 14984 11940 14988 11996
rect 14924 11936 14988 11940
rect 15004 11996 15068 12000
rect 15004 11940 15008 11996
rect 15008 11940 15064 11996
rect 15064 11940 15068 11996
rect 15004 11936 15068 11940
rect 15084 11996 15148 12000
rect 15084 11940 15088 11996
rect 15088 11940 15144 11996
rect 15144 11940 15148 11996
rect 15084 11936 15148 11940
rect 21790 11996 21854 12000
rect 21790 11940 21794 11996
rect 21794 11940 21850 11996
rect 21850 11940 21854 11996
rect 21790 11936 21854 11940
rect 21870 11996 21934 12000
rect 21870 11940 21874 11996
rect 21874 11940 21930 11996
rect 21930 11940 21934 11996
rect 21870 11936 21934 11940
rect 21950 11996 22014 12000
rect 21950 11940 21954 11996
rect 21954 11940 22010 11996
rect 22010 11940 22014 11996
rect 21950 11936 22014 11940
rect 22030 11996 22094 12000
rect 22030 11940 22034 11996
rect 22034 11940 22090 11996
rect 22090 11940 22094 11996
rect 22030 11936 22094 11940
rect 28736 11996 28800 12000
rect 28736 11940 28740 11996
rect 28740 11940 28796 11996
rect 28796 11940 28800 11996
rect 28736 11936 28800 11940
rect 28816 11996 28880 12000
rect 28816 11940 28820 11996
rect 28820 11940 28876 11996
rect 28876 11940 28880 11996
rect 28816 11936 28880 11940
rect 28896 11996 28960 12000
rect 28896 11940 28900 11996
rect 28900 11940 28956 11996
rect 28956 11940 28960 11996
rect 28896 11936 28960 11940
rect 28976 11996 29040 12000
rect 28976 11940 28980 11996
rect 28980 11940 29036 11996
rect 29036 11940 29040 11996
rect 28976 11936 29040 11940
rect 4425 11452 4489 11456
rect 4425 11396 4429 11452
rect 4429 11396 4485 11452
rect 4485 11396 4489 11452
rect 4425 11392 4489 11396
rect 4505 11452 4569 11456
rect 4505 11396 4509 11452
rect 4509 11396 4565 11452
rect 4565 11396 4569 11452
rect 4505 11392 4569 11396
rect 4585 11452 4649 11456
rect 4585 11396 4589 11452
rect 4589 11396 4645 11452
rect 4645 11396 4649 11452
rect 4585 11392 4649 11396
rect 4665 11452 4729 11456
rect 4665 11396 4669 11452
rect 4669 11396 4725 11452
rect 4725 11396 4729 11452
rect 4665 11392 4729 11396
rect 11371 11452 11435 11456
rect 11371 11396 11375 11452
rect 11375 11396 11431 11452
rect 11431 11396 11435 11452
rect 11371 11392 11435 11396
rect 11451 11452 11515 11456
rect 11451 11396 11455 11452
rect 11455 11396 11511 11452
rect 11511 11396 11515 11452
rect 11451 11392 11515 11396
rect 11531 11452 11595 11456
rect 11531 11396 11535 11452
rect 11535 11396 11591 11452
rect 11591 11396 11595 11452
rect 11531 11392 11595 11396
rect 11611 11452 11675 11456
rect 11611 11396 11615 11452
rect 11615 11396 11671 11452
rect 11671 11396 11675 11452
rect 11611 11392 11675 11396
rect 18317 11452 18381 11456
rect 18317 11396 18321 11452
rect 18321 11396 18377 11452
rect 18377 11396 18381 11452
rect 18317 11392 18381 11396
rect 18397 11452 18461 11456
rect 18397 11396 18401 11452
rect 18401 11396 18457 11452
rect 18457 11396 18461 11452
rect 18397 11392 18461 11396
rect 18477 11452 18541 11456
rect 18477 11396 18481 11452
rect 18481 11396 18537 11452
rect 18537 11396 18541 11452
rect 18477 11392 18541 11396
rect 18557 11452 18621 11456
rect 18557 11396 18561 11452
rect 18561 11396 18617 11452
rect 18617 11396 18621 11452
rect 18557 11392 18621 11396
rect 25263 11452 25327 11456
rect 25263 11396 25267 11452
rect 25267 11396 25323 11452
rect 25323 11396 25327 11452
rect 25263 11392 25327 11396
rect 25343 11452 25407 11456
rect 25343 11396 25347 11452
rect 25347 11396 25403 11452
rect 25403 11396 25407 11452
rect 25343 11392 25407 11396
rect 25423 11452 25487 11456
rect 25423 11396 25427 11452
rect 25427 11396 25483 11452
rect 25483 11396 25487 11452
rect 25423 11392 25487 11396
rect 25503 11452 25567 11456
rect 25503 11396 25507 11452
rect 25507 11396 25563 11452
rect 25563 11396 25567 11452
rect 25503 11392 25567 11396
rect 7898 10908 7962 10912
rect 7898 10852 7902 10908
rect 7902 10852 7958 10908
rect 7958 10852 7962 10908
rect 7898 10848 7962 10852
rect 7978 10908 8042 10912
rect 7978 10852 7982 10908
rect 7982 10852 8038 10908
rect 8038 10852 8042 10908
rect 7978 10848 8042 10852
rect 8058 10908 8122 10912
rect 8058 10852 8062 10908
rect 8062 10852 8118 10908
rect 8118 10852 8122 10908
rect 8058 10848 8122 10852
rect 8138 10908 8202 10912
rect 8138 10852 8142 10908
rect 8142 10852 8198 10908
rect 8198 10852 8202 10908
rect 8138 10848 8202 10852
rect 14844 10908 14908 10912
rect 14844 10852 14848 10908
rect 14848 10852 14904 10908
rect 14904 10852 14908 10908
rect 14844 10848 14908 10852
rect 14924 10908 14988 10912
rect 14924 10852 14928 10908
rect 14928 10852 14984 10908
rect 14984 10852 14988 10908
rect 14924 10848 14988 10852
rect 15004 10908 15068 10912
rect 15004 10852 15008 10908
rect 15008 10852 15064 10908
rect 15064 10852 15068 10908
rect 15004 10848 15068 10852
rect 15084 10908 15148 10912
rect 15084 10852 15088 10908
rect 15088 10852 15144 10908
rect 15144 10852 15148 10908
rect 15084 10848 15148 10852
rect 21790 10908 21854 10912
rect 21790 10852 21794 10908
rect 21794 10852 21850 10908
rect 21850 10852 21854 10908
rect 21790 10848 21854 10852
rect 21870 10908 21934 10912
rect 21870 10852 21874 10908
rect 21874 10852 21930 10908
rect 21930 10852 21934 10908
rect 21870 10848 21934 10852
rect 21950 10908 22014 10912
rect 21950 10852 21954 10908
rect 21954 10852 22010 10908
rect 22010 10852 22014 10908
rect 21950 10848 22014 10852
rect 22030 10908 22094 10912
rect 22030 10852 22034 10908
rect 22034 10852 22090 10908
rect 22090 10852 22094 10908
rect 22030 10848 22094 10852
rect 28736 10908 28800 10912
rect 28736 10852 28740 10908
rect 28740 10852 28796 10908
rect 28796 10852 28800 10908
rect 28736 10848 28800 10852
rect 28816 10908 28880 10912
rect 28816 10852 28820 10908
rect 28820 10852 28876 10908
rect 28876 10852 28880 10908
rect 28816 10848 28880 10852
rect 28896 10908 28960 10912
rect 28896 10852 28900 10908
rect 28900 10852 28956 10908
rect 28956 10852 28960 10908
rect 28896 10848 28960 10852
rect 28976 10908 29040 10912
rect 28976 10852 28980 10908
rect 28980 10852 29036 10908
rect 29036 10852 29040 10908
rect 28976 10848 29040 10852
rect 4425 10364 4489 10368
rect 4425 10308 4429 10364
rect 4429 10308 4485 10364
rect 4485 10308 4489 10364
rect 4425 10304 4489 10308
rect 4505 10364 4569 10368
rect 4505 10308 4509 10364
rect 4509 10308 4565 10364
rect 4565 10308 4569 10364
rect 4505 10304 4569 10308
rect 4585 10364 4649 10368
rect 4585 10308 4589 10364
rect 4589 10308 4645 10364
rect 4645 10308 4649 10364
rect 4585 10304 4649 10308
rect 4665 10364 4729 10368
rect 4665 10308 4669 10364
rect 4669 10308 4725 10364
rect 4725 10308 4729 10364
rect 4665 10304 4729 10308
rect 11371 10364 11435 10368
rect 11371 10308 11375 10364
rect 11375 10308 11431 10364
rect 11431 10308 11435 10364
rect 11371 10304 11435 10308
rect 11451 10364 11515 10368
rect 11451 10308 11455 10364
rect 11455 10308 11511 10364
rect 11511 10308 11515 10364
rect 11451 10304 11515 10308
rect 11531 10364 11595 10368
rect 11531 10308 11535 10364
rect 11535 10308 11591 10364
rect 11591 10308 11595 10364
rect 11531 10304 11595 10308
rect 11611 10364 11675 10368
rect 11611 10308 11615 10364
rect 11615 10308 11671 10364
rect 11671 10308 11675 10364
rect 11611 10304 11675 10308
rect 18317 10364 18381 10368
rect 18317 10308 18321 10364
rect 18321 10308 18377 10364
rect 18377 10308 18381 10364
rect 18317 10304 18381 10308
rect 18397 10364 18461 10368
rect 18397 10308 18401 10364
rect 18401 10308 18457 10364
rect 18457 10308 18461 10364
rect 18397 10304 18461 10308
rect 18477 10364 18541 10368
rect 18477 10308 18481 10364
rect 18481 10308 18537 10364
rect 18537 10308 18541 10364
rect 18477 10304 18541 10308
rect 18557 10364 18621 10368
rect 18557 10308 18561 10364
rect 18561 10308 18617 10364
rect 18617 10308 18621 10364
rect 18557 10304 18621 10308
rect 25263 10364 25327 10368
rect 25263 10308 25267 10364
rect 25267 10308 25323 10364
rect 25323 10308 25327 10364
rect 25263 10304 25327 10308
rect 25343 10364 25407 10368
rect 25343 10308 25347 10364
rect 25347 10308 25403 10364
rect 25403 10308 25407 10364
rect 25343 10304 25407 10308
rect 25423 10364 25487 10368
rect 25423 10308 25427 10364
rect 25427 10308 25483 10364
rect 25483 10308 25487 10364
rect 25423 10304 25487 10308
rect 25503 10364 25567 10368
rect 25503 10308 25507 10364
rect 25507 10308 25563 10364
rect 25563 10308 25567 10364
rect 25503 10304 25567 10308
rect 7898 9820 7962 9824
rect 7898 9764 7902 9820
rect 7902 9764 7958 9820
rect 7958 9764 7962 9820
rect 7898 9760 7962 9764
rect 7978 9820 8042 9824
rect 7978 9764 7982 9820
rect 7982 9764 8038 9820
rect 8038 9764 8042 9820
rect 7978 9760 8042 9764
rect 8058 9820 8122 9824
rect 8058 9764 8062 9820
rect 8062 9764 8118 9820
rect 8118 9764 8122 9820
rect 8058 9760 8122 9764
rect 8138 9820 8202 9824
rect 8138 9764 8142 9820
rect 8142 9764 8198 9820
rect 8198 9764 8202 9820
rect 8138 9760 8202 9764
rect 14844 9820 14908 9824
rect 14844 9764 14848 9820
rect 14848 9764 14904 9820
rect 14904 9764 14908 9820
rect 14844 9760 14908 9764
rect 14924 9820 14988 9824
rect 14924 9764 14928 9820
rect 14928 9764 14984 9820
rect 14984 9764 14988 9820
rect 14924 9760 14988 9764
rect 15004 9820 15068 9824
rect 15004 9764 15008 9820
rect 15008 9764 15064 9820
rect 15064 9764 15068 9820
rect 15004 9760 15068 9764
rect 15084 9820 15148 9824
rect 15084 9764 15088 9820
rect 15088 9764 15144 9820
rect 15144 9764 15148 9820
rect 15084 9760 15148 9764
rect 21790 9820 21854 9824
rect 21790 9764 21794 9820
rect 21794 9764 21850 9820
rect 21850 9764 21854 9820
rect 21790 9760 21854 9764
rect 21870 9820 21934 9824
rect 21870 9764 21874 9820
rect 21874 9764 21930 9820
rect 21930 9764 21934 9820
rect 21870 9760 21934 9764
rect 21950 9820 22014 9824
rect 21950 9764 21954 9820
rect 21954 9764 22010 9820
rect 22010 9764 22014 9820
rect 21950 9760 22014 9764
rect 22030 9820 22094 9824
rect 22030 9764 22034 9820
rect 22034 9764 22090 9820
rect 22090 9764 22094 9820
rect 22030 9760 22094 9764
rect 28736 9820 28800 9824
rect 28736 9764 28740 9820
rect 28740 9764 28796 9820
rect 28796 9764 28800 9820
rect 28736 9760 28800 9764
rect 28816 9820 28880 9824
rect 28816 9764 28820 9820
rect 28820 9764 28876 9820
rect 28876 9764 28880 9820
rect 28816 9760 28880 9764
rect 28896 9820 28960 9824
rect 28896 9764 28900 9820
rect 28900 9764 28956 9820
rect 28956 9764 28960 9820
rect 28896 9760 28960 9764
rect 28976 9820 29040 9824
rect 28976 9764 28980 9820
rect 28980 9764 29036 9820
rect 29036 9764 29040 9820
rect 28976 9760 29040 9764
rect 4425 9276 4489 9280
rect 4425 9220 4429 9276
rect 4429 9220 4485 9276
rect 4485 9220 4489 9276
rect 4425 9216 4489 9220
rect 4505 9276 4569 9280
rect 4505 9220 4509 9276
rect 4509 9220 4565 9276
rect 4565 9220 4569 9276
rect 4505 9216 4569 9220
rect 4585 9276 4649 9280
rect 4585 9220 4589 9276
rect 4589 9220 4645 9276
rect 4645 9220 4649 9276
rect 4585 9216 4649 9220
rect 4665 9276 4729 9280
rect 4665 9220 4669 9276
rect 4669 9220 4725 9276
rect 4725 9220 4729 9276
rect 4665 9216 4729 9220
rect 11371 9276 11435 9280
rect 11371 9220 11375 9276
rect 11375 9220 11431 9276
rect 11431 9220 11435 9276
rect 11371 9216 11435 9220
rect 11451 9276 11515 9280
rect 11451 9220 11455 9276
rect 11455 9220 11511 9276
rect 11511 9220 11515 9276
rect 11451 9216 11515 9220
rect 11531 9276 11595 9280
rect 11531 9220 11535 9276
rect 11535 9220 11591 9276
rect 11591 9220 11595 9276
rect 11531 9216 11595 9220
rect 11611 9276 11675 9280
rect 11611 9220 11615 9276
rect 11615 9220 11671 9276
rect 11671 9220 11675 9276
rect 11611 9216 11675 9220
rect 18317 9276 18381 9280
rect 18317 9220 18321 9276
rect 18321 9220 18377 9276
rect 18377 9220 18381 9276
rect 18317 9216 18381 9220
rect 18397 9276 18461 9280
rect 18397 9220 18401 9276
rect 18401 9220 18457 9276
rect 18457 9220 18461 9276
rect 18397 9216 18461 9220
rect 18477 9276 18541 9280
rect 18477 9220 18481 9276
rect 18481 9220 18537 9276
rect 18537 9220 18541 9276
rect 18477 9216 18541 9220
rect 18557 9276 18621 9280
rect 18557 9220 18561 9276
rect 18561 9220 18617 9276
rect 18617 9220 18621 9276
rect 18557 9216 18621 9220
rect 25263 9276 25327 9280
rect 25263 9220 25267 9276
rect 25267 9220 25323 9276
rect 25323 9220 25327 9276
rect 25263 9216 25327 9220
rect 25343 9276 25407 9280
rect 25343 9220 25347 9276
rect 25347 9220 25403 9276
rect 25403 9220 25407 9276
rect 25343 9216 25407 9220
rect 25423 9276 25487 9280
rect 25423 9220 25427 9276
rect 25427 9220 25483 9276
rect 25483 9220 25487 9276
rect 25423 9216 25487 9220
rect 25503 9276 25567 9280
rect 25503 9220 25507 9276
rect 25507 9220 25563 9276
rect 25563 9220 25567 9276
rect 25503 9216 25567 9220
rect 7898 8732 7962 8736
rect 7898 8676 7902 8732
rect 7902 8676 7958 8732
rect 7958 8676 7962 8732
rect 7898 8672 7962 8676
rect 7978 8732 8042 8736
rect 7978 8676 7982 8732
rect 7982 8676 8038 8732
rect 8038 8676 8042 8732
rect 7978 8672 8042 8676
rect 8058 8732 8122 8736
rect 8058 8676 8062 8732
rect 8062 8676 8118 8732
rect 8118 8676 8122 8732
rect 8058 8672 8122 8676
rect 8138 8732 8202 8736
rect 8138 8676 8142 8732
rect 8142 8676 8198 8732
rect 8198 8676 8202 8732
rect 8138 8672 8202 8676
rect 14844 8732 14908 8736
rect 14844 8676 14848 8732
rect 14848 8676 14904 8732
rect 14904 8676 14908 8732
rect 14844 8672 14908 8676
rect 14924 8732 14988 8736
rect 14924 8676 14928 8732
rect 14928 8676 14984 8732
rect 14984 8676 14988 8732
rect 14924 8672 14988 8676
rect 15004 8732 15068 8736
rect 15004 8676 15008 8732
rect 15008 8676 15064 8732
rect 15064 8676 15068 8732
rect 15004 8672 15068 8676
rect 15084 8732 15148 8736
rect 15084 8676 15088 8732
rect 15088 8676 15144 8732
rect 15144 8676 15148 8732
rect 15084 8672 15148 8676
rect 21790 8732 21854 8736
rect 21790 8676 21794 8732
rect 21794 8676 21850 8732
rect 21850 8676 21854 8732
rect 21790 8672 21854 8676
rect 21870 8732 21934 8736
rect 21870 8676 21874 8732
rect 21874 8676 21930 8732
rect 21930 8676 21934 8732
rect 21870 8672 21934 8676
rect 21950 8732 22014 8736
rect 21950 8676 21954 8732
rect 21954 8676 22010 8732
rect 22010 8676 22014 8732
rect 21950 8672 22014 8676
rect 22030 8732 22094 8736
rect 22030 8676 22034 8732
rect 22034 8676 22090 8732
rect 22090 8676 22094 8732
rect 22030 8672 22094 8676
rect 28736 8732 28800 8736
rect 28736 8676 28740 8732
rect 28740 8676 28796 8732
rect 28796 8676 28800 8732
rect 28736 8672 28800 8676
rect 28816 8732 28880 8736
rect 28816 8676 28820 8732
rect 28820 8676 28876 8732
rect 28876 8676 28880 8732
rect 28816 8672 28880 8676
rect 28896 8732 28960 8736
rect 28896 8676 28900 8732
rect 28900 8676 28956 8732
rect 28956 8676 28960 8732
rect 28896 8672 28960 8676
rect 28976 8732 29040 8736
rect 28976 8676 28980 8732
rect 28980 8676 29036 8732
rect 29036 8676 29040 8732
rect 28976 8672 29040 8676
rect 4425 8188 4489 8192
rect 4425 8132 4429 8188
rect 4429 8132 4485 8188
rect 4485 8132 4489 8188
rect 4425 8128 4489 8132
rect 4505 8188 4569 8192
rect 4505 8132 4509 8188
rect 4509 8132 4565 8188
rect 4565 8132 4569 8188
rect 4505 8128 4569 8132
rect 4585 8188 4649 8192
rect 4585 8132 4589 8188
rect 4589 8132 4645 8188
rect 4645 8132 4649 8188
rect 4585 8128 4649 8132
rect 4665 8188 4729 8192
rect 4665 8132 4669 8188
rect 4669 8132 4725 8188
rect 4725 8132 4729 8188
rect 4665 8128 4729 8132
rect 11371 8188 11435 8192
rect 11371 8132 11375 8188
rect 11375 8132 11431 8188
rect 11431 8132 11435 8188
rect 11371 8128 11435 8132
rect 11451 8188 11515 8192
rect 11451 8132 11455 8188
rect 11455 8132 11511 8188
rect 11511 8132 11515 8188
rect 11451 8128 11515 8132
rect 11531 8188 11595 8192
rect 11531 8132 11535 8188
rect 11535 8132 11591 8188
rect 11591 8132 11595 8188
rect 11531 8128 11595 8132
rect 11611 8188 11675 8192
rect 11611 8132 11615 8188
rect 11615 8132 11671 8188
rect 11671 8132 11675 8188
rect 11611 8128 11675 8132
rect 18317 8188 18381 8192
rect 18317 8132 18321 8188
rect 18321 8132 18377 8188
rect 18377 8132 18381 8188
rect 18317 8128 18381 8132
rect 18397 8188 18461 8192
rect 18397 8132 18401 8188
rect 18401 8132 18457 8188
rect 18457 8132 18461 8188
rect 18397 8128 18461 8132
rect 18477 8188 18541 8192
rect 18477 8132 18481 8188
rect 18481 8132 18537 8188
rect 18537 8132 18541 8188
rect 18477 8128 18541 8132
rect 18557 8188 18621 8192
rect 18557 8132 18561 8188
rect 18561 8132 18617 8188
rect 18617 8132 18621 8188
rect 18557 8128 18621 8132
rect 25263 8188 25327 8192
rect 25263 8132 25267 8188
rect 25267 8132 25323 8188
rect 25323 8132 25327 8188
rect 25263 8128 25327 8132
rect 25343 8188 25407 8192
rect 25343 8132 25347 8188
rect 25347 8132 25403 8188
rect 25403 8132 25407 8188
rect 25343 8128 25407 8132
rect 25423 8188 25487 8192
rect 25423 8132 25427 8188
rect 25427 8132 25483 8188
rect 25483 8132 25487 8188
rect 25423 8128 25487 8132
rect 25503 8188 25567 8192
rect 25503 8132 25507 8188
rect 25507 8132 25563 8188
rect 25563 8132 25567 8188
rect 25503 8128 25567 8132
rect 7898 7644 7962 7648
rect 7898 7588 7902 7644
rect 7902 7588 7958 7644
rect 7958 7588 7962 7644
rect 7898 7584 7962 7588
rect 7978 7644 8042 7648
rect 7978 7588 7982 7644
rect 7982 7588 8038 7644
rect 8038 7588 8042 7644
rect 7978 7584 8042 7588
rect 8058 7644 8122 7648
rect 8058 7588 8062 7644
rect 8062 7588 8118 7644
rect 8118 7588 8122 7644
rect 8058 7584 8122 7588
rect 8138 7644 8202 7648
rect 8138 7588 8142 7644
rect 8142 7588 8198 7644
rect 8198 7588 8202 7644
rect 8138 7584 8202 7588
rect 14844 7644 14908 7648
rect 14844 7588 14848 7644
rect 14848 7588 14904 7644
rect 14904 7588 14908 7644
rect 14844 7584 14908 7588
rect 14924 7644 14988 7648
rect 14924 7588 14928 7644
rect 14928 7588 14984 7644
rect 14984 7588 14988 7644
rect 14924 7584 14988 7588
rect 15004 7644 15068 7648
rect 15004 7588 15008 7644
rect 15008 7588 15064 7644
rect 15064 7588 15068 7644
rect 15004 7584 15068 7588
rect 15084 7644 15148 7648
rect 15084 7588 15088 7644
rect 15088 7588 15144 7644
rect 15144 7588 15148 7644
rect 15084 7584 15148 7588
rect 21790 7644 21854 7648
rect 21790 7588 21794 7644
rect 21794 7588 21850 7644
rect 21850 7588 21854 7644
rect 21790 7584 21854 7588
rect 21870 7644 21934 7648
rect 21870 7588 21874 7644
rect 21874 7588 21930 7644
rect 21930 7588 21934 7644
rect 21870 7584 21934 7588
rect 21950 7644 22014 7648
rect 21950 7588 21954 7644
rect 21954 7588 22010 7644
rect 22010 7588 22014 7644
rect 21950 7584 22014 7588
rect 22030 7644 22094 7648
rect 22030 7588 22034 7644
rect 22034 7588 22090 7644
rect 22090 7588 22094 7644
rect 22030 7584 22094 7588
rect 28736 7644 28800 7648
rect 28736 7588 28740 7644
rect 28740 7588 28796 7644
rect 28796 7588 28800 7644
rect 28736 7584 28800 7588
rect 28816 7644 28880 7648
rect 28816 7588 28820 7644
rect 28820 7588 28876 7644
rect 28876 7588 28880 7644
rect 28816 7584 28880 7588
rect 28896 7644 28960 7648
rect 28896 7588 28900 7644
rect 28900 7588 28956 7644
rect 28956 7588 28960 7644
rect 28896 7584 28960 7588
rect 28976 7644 29040 7648
rect 28976 7588 28980 7644
rect 28980 7588 29036 7644
rect 29036 7588 29040 7644
rect 28976 7584 29040 7588
rect 4425 7100 4489 7104
rect 4425 7044 4429 7100
rect 4429 7044 4485 7100
rect 4485 7044 4489 7100
rect 4425 7040 4489 7044
rect 4505 7100 4569 7104
rect 4505 7044 4509 7100
rect 4509 7044 4565 7100
rect 4565 7044 4569 7100
rect 4505 7040 4569 7044
rect 4585 7100 4649 7104
rect 4585 7044 4589 7100
rect 4589 7044 4645 7100
rect 4645 7044 4649 7100
rect 4585 7040 4649 7044
rect 4665 7100 4729 7104
rect 4665 7044 4669 7100
rect 4669 7044 4725 7100
rect 4725 7044 4729 7100
rect 4665 7040 4729 7044
rect 11371 7100 11435 7104
rect 11371 7044 11375 7100
rect 11375 7044 11431 7100
rect 11431 7044 11435 7100
rect 11371 7040 11435 7044
rect 11451 7100 11515 7104
rect 11451 7044 11455 7100
rect 11455 7044 11511 7100
rect 11511 7044 11515 7100
rect 11451 7040 11515 7044
rect 11531 7100 11595 7104
rect 11531 7044 11535 7100
rect 11535 7044 11591 7100
rect 11591 7044 11595 7100
rect 11531 7040 11595 7044
rect 11611 7100 11675 7104
rect 11611 7044 11615 7100
rect 11615 7044 11671 7100
rect 11671 7044 11675 7100
rect 11611 7040 11675 7044
rect 18317 7100 18381 7104
rect 18317 7044 18321 7100
rect 18321 7044 18377 7100
rect 18377 7044 18381 7100
rect 18317 7040 18381 7044
rect 18397 7100 18461 7104
rect 18397 7044 18401 7100
rect 18401 7044 18457 7100
rect 18457 7044 18461 7100
rect 18397 7040 18461 7044
rect 18477 7100 18541 7104
rect 18477 7044 18481 7100
rect 18481 7044 18537 7100
rect 18537 7044 18541 7100
rect 18477 7040 18541 7044
rect 18557 7100 18621 7104
rect 18557 7044 18561 7100
rect 18561 7044 18617 7100
rect 18617 7044 18621 7100
rect 18557 7040 18621 7044
rect 25263 7100 25327 7104
rect 25263 7044 25267 7100
rect 25267 7044 25323 7100
rect 25323 7044 25327 7100
rect 25263 7040 25327 7044
rect 25343 7100 25407 7104
rect 25343 7044 25347 7100
rect 25347 7044 25403 7100
rect 25403 7044 25407 7100
rect 25343 7040 25407 7044
rect 25423 7100 25487 7104
rect 25423 7044 25427 7100
rect 25427 7044 25483 7100
rect 25483 7044 25487 7100
rect 25423 7040 25487 7044
rect 25503 7100 25567 7104
rect 25503 7044 25507 7100
rect 25507 7044 25563 7100
rect 25563 7044 25567 7100
rect 25503 7040 25567 7044
rect 7898 6556 7962 6560
rect 7898 6500 7902 6556
rect 7902 6500 7958 6556
rect 7958 6500 7962 6556
rect 7898 6496 7962 6500
rect 7978 6556 8042 6560
rect 7978 6500 7982 6556
rect 7982 6500 8038 6556
rect 8038 6500 8042 6556
rect 7978 6496 8042 6500
rect 8058 6556 8122 6560
rect 8058 6500 8062 6556
rect 8062 6500 8118 6556
rect 8118 6500 8122 6556
rect 8058 6496 8122 6500
rect 8138 6556 8202 6560
rect 8138 6500 8142 6556
rect 8142 6500 8198 6556
rect 8198 6500 8202 6556
rect 8138 6496 8202 6500
rect 14844 6556 14908 6560
rect 14844 6500 14848 6556
rect 14848 6500 14904 6556
rect 14904 6500 14908 6556
rect 14844 6496 14908 6500
rect 14924 6556 14988 6560
rect 14924 6500 14928 6556
rect 14928 6500 14984 6556
rect 14984 6500 14988 6556
rect 14924 6496 14988 6500
rect 15004 6556 15068 6560
rect 15004 6500 15008 6556
rect 15008 6500 15064 6556
rect 15064 6500 15068 6556
rect 15004 6496 15068 6500
rect 15084 6556 15148 6560
rect 15084 6500 15088 6556
rect 15088 6500 15144 6556
rect 15144 6500 15148 6556
rect 15084 6496 15148 6500
rect 21790 6556 21854 6560
rect 21790 6500 21794 6556
rect 21794 6500 21850 6556
rect 21850 6500 21854 6556
rect 21790 6496 21854 6500
rect 21870 6556 21934 6560
rect 21870 6500 21874 6556
rect 21874 6500 21930 6556
rect 21930 6500 21934 6556
rect 21870 6496 21934 6500
rect 21950 6556 22014 6560
rect 21950 6500 21954 6556
rect 21954 6500 22010 6556
rect 22010 6500 22014 6556
rect 21950 6496 22014 6500
rect 22030 6556 22094 6560
rect 22030 6500 22034 6556
rect 22034 6500 22090 6556
rect 22090 6500 22094 6556
rect 22030 6496 22094 6500
rect 28736 6556 28800 6560
rect 28736 6500 28740 6556
rect 28740 6500 28796 6556
rect 28796 6500 28800 6556
rect 28736 6496 28800 6500
rect 28816 6556 28880 6560
rect 28816 6500 28820 6556
rect 28820 6500 28876 6556
rect 28876 6500 28880 6556
rect 28816 6496 28880 6500
rect 28896 6556 28960 6560
rect 28896 6500 28900 6556
rect 28900 6500 28956 6556
rect 28956 6500 28960 6556
rect 28896 6496 28960 6500
rect 28976 6556 29040 6560
rect 28976 6500 28980 6556
rect 28980 6500 29036 6556
rect 29036 6500 29040 6556
rect 28976 6496 29040 6500
rect 4425 6012 4489 6016
rect 4425 5956 4429 6012
rect 4429 5956 4485 6012
rect 4485 5956 4489 6012
rect 4425 5952 4489 5956
rect 4505 6012 4569 6016
rect 4505 5956 4509 6012
rect 4509 5956 4565 6012
rect 4565 5956 4569 6012
rect 4505 5952 4569 5956
rect 4585 6012 4649 6016
rect 4585 5956 4589 6012
rect 4589 5956 4645 6012
rect 4645 5956 4649 6012
rect 4585 5952 4649 5956
rect 4665 6012 4729 6016
rect 4665 5956 4669 6012
rect 4669 5956 4725 6012
rect 4725 5956 4729 6012
rect 4665 5952 4729 5956
rect 11371 6012 11435 6016
rect 11371 5956 11375 6012
rect 11375 5956 11431 6012
rect 11431 5956 11435 6012
rect 11371 5952 11435 5956
rect 11451 6012 11515 6016
rect 11451 5956 11455 6012
rect 11455 5956 11511 6012
rect 11511 5956 11515 6012
rect 11451 5952 11515 5956
rect 11531 6012 11595 6016
rect 11531 5956 11535 6012
rect 11535 5956 11591 6012
rect 11591 5956 11595 6012
rect 11531 5952 11595 5956
rect 11611 6012 11675 6016
rect 11611 5956 11615 6012
rect 11615 5956 11671 6012
rect 11671 5956 11675 6012
rect 11611 5952 11675 5956
rect 18317 6012 18381 6016
rect 18317 5956 18321 6012
rect 18321 5956 18377 6012
rect 18377 5956 18381 6012
rect 18317 5952 18381 5956
rect 18397 6012 18461 6016
rect 18397 5956 18401 6012
rect 18401 5956 18457 6012
rect 18457 5956 18461 6012
rect 18397 5952 18461 5956
rect 18477 6012 18541 6016
rect 18477 5956 18481 6012
rect 18481 5956 18537 6012
rect 18537 5956 18541 6012
rect 18477 5952 18541 5956
rect 18557 6012 18621 6016
rect 18557 5956 18561 6012
rect 18561 5956 18617 6012
rect 18617 5956 18621 6012
rect 18557 5952 18621 5956
rect 25263 6012 25327 6016
rect 25263 5956 25267 6012
rect 25267 5956 25323 6012
rect 25323 5956 25327 6012
rect 25263 5952 25327 5956
rect 25343 6012 25407 6016
rect 25343 5956 25347 6012
rect 25347 5956 25403 6012
rect 25403 5956 25407 6012
rect 25343 5952 25407 5956
rect 25423 6012 25487 6016
rect 25423 5956 25427 6012
rect 25427 5956 25483 6012
rect 25483 5956 25487 6012
rect 25423 5952 25487 5956
rect 25503 6012 25567 6016
rect 25503 5956 25507 6012
rect 25507 5956 25563 6012
rect 25563 5956 25567 6012
rect 25503 5952 25567 5956
rect 7898 5468 7962 5472
rect 7898 5412 7902 5468
rect 7902 5412 7958 5468
rect 7958 5412 7962 5468
rect 7898 5408 7962 5412
rect 7978 5468 8042 5472
rect 7978 5412 7982 5468
rect 7982 5412 8038 5468
rect 8038 5412 8042 5468
rect 7978 5408 8042 5412
rect 8058 5468 8122 5472
rect 8058 5412 8062 5468
rect 8062 5412 8118 5468
rect 8118 5412 8122 5468
rect 8058 5408 8122 5412
rect 8138 5468 8202 5472
rect 8138 5412 8142 5468
rect 8142 5412 8198 5468
rect 8198 5412 8202 5468
rect 8138 5408 8202 5412
rect 14844 5468 14908 5472
rect 14844 5412 14848 5468
rect 14848 5412 14904 5468
rect 14904 5412 14908 5468
rect 14844 5408 14908 5412
rect 14924 5468 14988 5472
rect 14924 5412 14928 5468
rect 14928 5412 14984 5468
rect 14984 5412 14988 5468
rect 14924 5408 14988 5412
rect 15004 5468 15068 5472
rect 15004 5412 15008 5468
rect 15008 5412 15064 5468
rect 15064 5412 15068 5468
rect 15004 5408 15068 5412
rect 15084 5468 15148 5472
rect 15084 5412 15088 5468
rect 15088 5412 15144 5468
rect 15144 5412 15148 5468
rect 15084 5408 15148 5412
rect 21790 5468 21854 5472
rect 21790 5412 21794 5468
rect 21794 5412 21850 5468
rect 21850 5412 21854 5468
rect 21790 5408 21854 5412
rect 21870 5468 21934 5472
rect 21870 5412 21874 5468
rect 21874 5412 21930 5468
rect 21930 5412 21934 5468
rect 21870 5408 21934 5412
rect 21950 5468 22014 5472
rect 21950 5412 21954 5468
rect 21954 5412 22010 5468
rect 22010 5412 22014 5468
rect 21950 5408 22014 5412
rect 22030 5468 22094 5472
rect 22030 5412 22034 5468
rect 22034 5412 22090 5468
rect 22090 5412 22094 5468
rect 22030 5408 22094 5412
rect 28736 5468 28800 5472
rect 28736 5412 28740 5468
rect 28740 5412 28796 5468
rect 28796 5412 28800 5468
rect 28736 5408 28800 5412
rect 28816 5468 28880 5472
rect 28816 5412 28820 5468
rect 28820 5412 28876 5468
rect 28876 5412 28880 5468
rect 28816 5408 28880 5412
rect 28896 5468 28960 5472
rect 28896 5412 28900 5468
rect 28900 5412 28956 5468
rect 28956 5412 28960 5468
rect 28896 5408 28960 5412
rect 28976 5468 29040 5472
rect 28976 5412 28980 5468
rect 28980 5412 29036 5468
rect 29036 5412 29040 5468
rect 28976 5408 29040 5412
rect 4425 4924 4489 4928
rect 4425 4868 4429 4924
rect 4429 4868 4485 4924
rect 4485 4868 4489 4924
rect 4425 4864 4489 4868
rect 4505 4924 4569 4928
rect 4505 4868 4509 4924
rect 4509 4868 4565 4924
rect 4565 4868 4569 4924
rect 4505 4864 4569 4868
rect 4585 4924 4649 4928
rect 4585 4868 4589 4924
rect 4589 4868 4645 4924
rect 4645 4868 4649 4924
rect 4585 4864 4649 4868
rect 4665 4924 4729 4928
rect 4665 4868 4669 4924
rect 4669 4868 4725 4924
rect 4725 4868 4729 4924
rect 4665 4864 4729 4868
rect 11371 4924 11435 4928
rect 11371 4868 11375 4924
rect 11375 4868 11431 4924
rect 11431 4868 11435 4924
rect 11371 4864 11435 4868
rect 11451 4924 11515 4928
rect 11451 4868 11455 4924
rect 11455 4868 11511 4924
rect 11511 4868 11515 4924
rect 11451 4864 11515 4868
rect 11531 4924 11595 4928
rect 11531 4868 11535 4924
rect 11535 4868 11591 4924
rect 11591 4868 11595 4924
rect 11531 4864 11595 4868
rect 11611 4924 11675 4928
rect 11611 4868 11615 4924
rect 11615 4868 11671 4924
rect 11671 4868 11675 4924
rect 11611 4864 11675 4868
rect 18317 4924 18381 4928
rect 18317 4868 18321 4924
rect 18321 4868 18377 4924
rect 18377 4868 18381 4924
rect 18317 4864 18381 4868
rect 18397 4924 18461 4928
rect 18397 4868 18401 4924
rect 18401 4868 18457 4924
rect 18457 4868 18461 4924
rect 18397 4864 18461 4868
rect 18477 4924 18541 4928
rect 18477 4868 18481 4924
rect 18481 4868 18537 4924
rect 18537 4868 18541 4924
rect 18477 4864 18541 4868
rect 18557 4924 18621 4928
rect 18557 4868 18561 4924
rect 18561 4868 18617 4924
rect 18617 4868 18621 4924
rect 18557 4864 18621 4868
rect 25263 4924 25327 4928
rect 25263 4868 25267 4924
rect 25267 4868 25323 4924
rect 25323 4868 25327 4924
rect 25263 4864 25327 4868
rect 25343 4924 25407 4928
rect 25343 4868 25347 4924
rect 25347 4868 25403 4924
rect 25403 4868 25407 4924
rect 25343 4864 25407 4868
rect 25423 4924 25487 4928
rect 25423 4868 25427 4924
rect 25427 4868 25483 4924
rect 25483 4868 25487 4924
rect 25423 4864 25487 4868
rect 25503 4924 25567 4928
rect 25503 4868 25507 4924
rect 25507 4868 25563 4924
rect 25563 4868 25567 4924
rect 25503 4864 25567 4868
rect 7898 4380 7962 4384
rect 7898 4324 7902 4380
rect 7902 4324 7958 4380
rect 7958 4324 7962 4380
rect 7898 4320 7962 4324
rect 7978 4380 8042 4384
rect 7978 4324 7982 4380
rect 7982 4324 8038 4380
rect 8038 4324 8042 4380
rect 7978 4320 8042 4324
rect 8058 4380 8122 4384
rect 8058 4324 8062 4380
rect 8062 4324 8118 4380
rect 8118 4324 8122 4380
rect 8058 4320 8122 4324
rect 8138 4380 8202 4384
rect 8138 4324 8142 4380
rect 8142 4324 8198 4380
rect 8198 4324 8202 4380
rect 8138 4320 8202 4324
rect 14844 4380 14908 4384
rect 14844 4324 14848 4380
rect 14848 4324 14904 4380
rect 14904 4324 14908 4380
rect 14844 4320 14908 4324
rect 14924 4380 14988 4384
rect 14924 4324 14928 4380
rect 14928 4324 14984 4380
rect 14984 4324 14988 4380
rect 14924 4320 14988 4324
rect 15004 4380 15068 4384
rect 15004 4324 15008 4380
rect 15008 4324 15064 4380
rect 15064 4324 15068 4380
rect 15004 4320 15068 4324
rect 15084 4380 15148 4384
rect 15084 4324 15088 4380
rect 15088 4324 15144 4380
rect 15144 4324 15148 4380
rect 15084 4320 15148 4324
rect 21790 4380 21854 4384
rect 21790 4324 21794 4380
rect 21794 4324 21850 4380
rect 21850 4324 21854 4380
rect 21790 4320 21854 4324
rect 21870 4380 21934 4384
rect 21870 4324 21874 4380
rect 21874 4324 21930 4380
rect 21930 4324 21934 4380
rect 21870 4320 21934 4324
rect 21950 4380 22014 4384
rect 21950 4324 21954 4380
rect 21954 4324 22010 4380
rect 22010 4324 22014 4380
rect 21950 4320 22014 4324
rect 22030 4380 22094 4384
rect 22030 4324 22034 4380
rect 22034 4324 22090 4380
rect 22090 4324 22094 4380
rect 22030 4320 22094 4324
rect 28736 4380 28800 4384
rect 28736 4324 28740 4380
rect 28740 4324 28796 4380
rect 28796 4324 28800 4380
rect 28736 4320 28800 4324
rect 28816 4380 28880 4384
rect 28816 4324 28820 4380
rect 28820 4324 28876 4380
rect 28876 4324 28880 4380
rect 28816 4320 28880 4324
rect 28896 4380 28960 4384
rect 28896 4324 28900 4380
rect 28900 4324 28956 4380
rect 28956 4324 28960 4380
rect 28896 4320 28960 4324
rect 28976 4380 29040 4384
rect 28976 4324 28980 4380
rect 28980 4324 29036 4380
rect 29036 4324 29040 4380
rect 28976 4320 29040 4324
rect 4425 3836 4489 3840
rect 4425 3780 4429 3836
rect 4429 3780 4485 3836
rect 4485 3780 4489 3836
rect 4425 3776 4489 3780
rect 4505 3836 4569 3840
rect 4505 3780 4509 3836
rect 4509 3780 4565 3836
rect 4565 3780 4569 3836
rect 4505 3776 4569 3780
rect 4585 3836 4649 3840
rect 4585 3780 4589 3836
rect 4589 3780 4645 3836
rect 4645 3780 4649 3836
rect 4585 3776 4649 3780
rect 4665 3836 4729 3840
rect 4665 3780 4669 3836
rect 4669 3780 4725 3836
rect 4725 3780 4729 3836
rect 4665 3776 4729 3780
rect 11371 3836 11435 3840
rect 11371 3780 11375 3836
rect 11375 3780 11431 3836
rect 11431 3780 11435 3836
rect 11371 3776 11435 3780
rect 11451 3836 11515 3840
rect 11451 3780 11455 3836
rect 11455 3780 11511 3836
rect 11511 3780 11515 3836
rect 11451 3776 11515 3780
rect 11531 3836 11595 3840
rect 11531 3780 11535 3836
rect 11535 3780 11591 3836
rect 11591 3780 11595 3836
rect 11531 3776 11595 3780
rect 11611 3836 11675 3840
rect 11611 3780 11615 3836
rect 11615 3780 11671 3836
rect 11671 3780 11675 3836
rect 11611 3776 11675 3780
rect 18317 3836 18381 3840
rect 18317 3780 18321 3836
rect 18321 3780 18377 3836
rect 18377 3780 18381 3836
rect 18317 3776 18381 3780
rect 18397 3836 18461 3840
rect 18397 3780 18401 3836
rect 18401 3780 18457 3836
rect 18457 3780 18461 3836
rect 18397 3776 18461 3780
rect 18477 3836 18541 3840
rect 18477 3780 18481 3836
rect 18481 3780 18537 3836
rect 18537 3780 18541 3836
rect 18477 3776 18541 3780
rect 18557 3836 18621 3840
rect 18557 3780 18561 3836
rect 18561 3780 18617 3836
rect 18617 3780 18621 3836
rect 18557 3776 18621 3780
rect 25263 3836 25327 3840
rect 25263 3780 25267 3836
rect 25267 3780 25323 3836
rect 25323 3780 25327 3836
rect 25263 3776 25327 3780
rect 25343 3836 25407 3840
rect 25343 3780 25347 3836
rect 25347 3780 25403 3836
rect 25403 3780 25407 3836
rect 25343 3776 25407 3780
rect 25423 3836 25487 3840
rect 25423 3780 25427 3836
rect 25427 3780 25483 3836
rect 25483 3780 25487 3836
rect 25423 3776 25487 3780
rect 25503 3836 25567 3840
rect 25503 3780 25507 3836
rect 25507 3780 25563 3836
rect 25563 3780 25567 3836
rect 25503 3776 25567 3780
rect 7898 3292 7962 3296
rect 7898 3236 7902 3292
rect 7902 3236 7958 3292
rect 7958 3236 7962 3292
rect 7898 3232 7962 3236
rect 7978 3292 8042 3296
rect 7978 3236 7982 3292
rect 7982 3236 8038 3292
rect 8038 3236 8042 3292
rect 7978 3232 8042 3236
rect 8058 3292 8122 3296
rect 8058 3236 8062 3292
rect 8062 3236 8118 3292
rect 8118 3236 8122 3292
rect 8058 3232 8122 3236
rect 8138 3292 8202 3296
rect 8138 3236 8142 3292
rect 8142 3236 8198 3292
rect 8198 3236 8202 3292
rect 8138 3232 8202 3236
rect 14844 3292 14908 3296
rect 14844 3236 14848 3292
rect 14848 3236 14904 3292
rect 14904 3236 14908 3292
rect 14844 3232 14908 3236
rect 14924 3292 14988 3296
rect 14924 3236 14928 3292
rect 14928 3236 14984 3292
rect 14984 3236 14988 3292
rect 14924 3232 14988 3236
rect 15004 3292 15068 3296
rect 15004 3236 15008 3292
rect 15008 3236 15064 3292
rect 15064 3236 15068 3292
rect 15004 3232 15068 3236
rect 15084 3292 15148 3296
rect 15084 3236 15088 3292
rect 15088 3236 15144 3292
rect 15144 3236 15148 3292
rect 15084 3232 15148 3236
rect 21790 3292 21854 3296
rect 21790 3236 21794 3292
rect 21794 3236 21850 3292
rect 21850 3236 21854 3292
rect 21790 3232 21854 3236
rect 21870 3292 21934 3296
rect 21870 3236 21874 3292
rect 21874 3236 21930 3292
rect 21930 3236 21934 3292
rect 21870 3232 21934 3236
rect 21950 3292 22014 3296
rect 21950 3236 21954 3292
rect 21954 3236 22010 3292
rect 22010 3236 22014 3292
rect 21950 3232 22014 3236
rect 22030 3292 22094 3296
rect 22030 3236 22034 3292
rect 22034 3236 22090 3292
rect 22090 3236 22094 3292
rect 22030 3232 22094 3236
rect 28736 3292 28800 3296
rect 28736 3236 28740 3292
rect 28740 3236 28796 3292
rect 28796 3236 28800 3292
rect 28736 3232 28800 3236
rect 28816 3292 28880 3296
rect 28816 3236 28820 3292
rect 28820 3236 28876 3292
rect 28876 3236 28880 3292
rect 28816 3232 28880 3236
rect 28896 3292 28960 3296
rect 28896 3236 28900 3292
rect 28900 3236 28956 3292
rect 28956 3236 28960 3292
rect 28896 3232 28960 3236
rect 28976 3292 29040 3296
rect 28976 3236 28980 3292
rect 28980 3236 29036 3292
rect 29036 3236 29040 3292
rect 28976 3232 29040 3236
rect 4425 2748 4489 2752
rect 4425 2692 4429 2748
rect 4429 2692 4485 2748
rect 4485 2692 4489 2748
rect 4425 2688 4489 2692
rect 4505 2748 4569 2752
rect 4505 2692 4509 2748
rect 4509 2692 4565 2748
rect 4565 2692 4569 2748
rect 4505 2688 4569 2692
rect 4585 2748 4649 2752
rect 4585 2692 4589 2748
rect 4589 2692 4645 2748
rect 4645 2692 4649 2748
rect 4585 2688 4649 2692
rect 4665 2748 4729 2752
rect 4665 2692 4669 2748
rect 4669 2692 4725 2748
rect 4725 2692 4729 2748
rect 4665 2688 4729 2692
rect 11371 2748 11435 2752
rect 11371 2692 11375 2748
rect 11375 2692 11431 2748
rect 11431 2692 11435 2748
rect 11371 2688 11435 2692
rect 11451 2748 11515 2752
rect 11451 2692 11455 2748
rect 11455 2692 11511 2748
rect 11511 2692 11515 2748
rect 11451 2688 11515 2692
rect 11531 2748 11595 2752
rect 11531 2692 11535 2748
rect 11535 2692 11591 2748
rect 11591 2692 11595 2748
rect 11531 2688 11595 2692
rect 11611 2748 11675 2752
rect 11611 2692 11615 2748
rect 11615 2692 11671 2748
rect 11671 2692 11675 2748
rect 11611 2688 11675 2692
rect 18317 2748 18381 2752
rect 18317 2692 18321 2748
rect 18321 2692 18377 2748
rect 18377 2692 18381 2748
rect 18317 2688 18381 2692
rect 18397 2748 18461 2752
rect 18397 2692 18401 2748
rect 18401 2692 18457 2748
rect 18457 2692 18461 2748
rect 18397 2688 18461 2692
rect 18477 2748 18541 2752
rect 18477 2692 18481 2748
rect 18481 2692 18537 2748
rect 18537 2692 18541 2748
rect 18477 2688 18541 2692
rect 18557 2748 18621 2752
rect 18557 2692 18561 2748
rect 18561 2692 18617 2748
rect 18617 2692 18621 2748
rect 18557 2688 18621 2692
rect 25263 2748 25327 2752
rect 25263 2692 25267 2748
rect 25267 2692 25323 2748
rect 25323 2692 25327 2748
rect 25263 2688 25327 2692
rect 25343 2748 25407 2752
rect 25343 2692 25347 2748
rect 25347 2692 25403 2748
rect 25403 2692 25407 2748
rect 25343 2688 25407 2692
rect 25423 2748 25487 2752
rect 25423 2692 25427 2748
rect 25427 2692 25483 2748
rect 25483 2692 25487 2748
rect 25423 2688 25487 2692
rect 25503 2748 25567 2752
rect 25503 2692 25507 2748
rect 25507 2692 25563 2748
rect 25563 2692 25567 2748
rect 25503 2688 25567 2692
rect 7898 2204 7962 2208
rect 7898 2148 7902 2204
rect 7902 2148 7958 2204
rect 7958 2148 7962 2204
rect 7898 2144 7962 2148
rect 7978 2204 8042 2208
rect 7978 2148 7982 2204
rect 7982 2148 8038 2204
rect 8038 2148 8042 2204
rect 7978 2144 8042 2148
rect 8058 2204 8122 2208
rect 8058 2148 8062 2204
rect 8062 2148 8118 2204
rect 8118 2148 8122 2204
rect 8058 2144 8122 2148
rect 8138 2204 8202 2208
rect 8138 2148 8142 2204
rect 8142 2148 8198 2204
rect 8198 2148 8202 2204
rect 8138 2144 8202 2148
rect 14844 2204 14908 2208
rect 14844 2148 14848 2204
rect 14848 2148 14904 2204
rect 14904 2148 14908 2204
rect 14844 2144 14908 2148
rect 14924 2204 14988 2208
rect 14924 2148 14928 2204
rect 14928 2148 14984 2204
rect 14984 2148 14988 2204
rect 14924 2144 14988 2148
rect 15004 2204 15068 2208
rect 15004 2148 15008 2204
rect 15008 2148 15064 2204
rect 15064 2148 15068 2204
rect 15004 2144 15068 2148
rect 15084 2204 15148 2208
rect 15084 2148 15088 2204
rect 15088 2148 15144 2204
rect 15144 2148 15148 2204
rect 15084 2144 15148 2148
rect 21790 2204 21854 2208
rect 21790 2148 21794 2204
rect 21794 2148 21850 2204
rect 21850 2148 21854 2204
rect 21790 2144 21854 2148
rect 21870 2204 21934 2208
rect 21870 2148 21874 2204
rect 21874 2148 21930 2204
rect 21930 2148 21934 2204
rect 21870 2144 21934 2148
rect 21950 2204 22014 2208
rect 21950 2148 21954 2204
rect 21954 2148 22010 2204
rect 22010 2148 22014 2204
rect 21950 2144 22014 2148
rect 22030 2204 22094 2208
rect 22030 2148 22034 2204
rect 22034 2148 22090 2204
rect 22090 2148 22094 2204
rect 22030 2144 22094 2148
rect 28736 2204 28800 2208
rect 28736 2148 28740 2204
rect 28740 2148 28796 2204
rect 28796 2148 28800 2204
rect 28736 2144 28800 2148
rect 28816 2204 28880 2208
rect 28816 2148 28820 2204
rect 28820 2148 28876 2204
rect 28876 2148 28880 2204
rect 28816 2144 28880 2148
rect 28896 2204 28960 2208
rect 28896 2148 28900 2204
rect 28900 2148 28956 2204
rect 28956 2148 28960 2204
rect 28896 2144 28960 2148
rect 28976 2204 29040 2208
rect 28976 2148 28980 2204
rect 28980 2148 29036 2204
rect 29036 2148 29040 2204
rect 28976 2144 29040 2148
<< metal4 >>
rect 4417 47360 4737 47376
rect 4417 47296 4425 47360
rect 4489 47296 4505 47360
rect 4569 47296 4585 47360
rect 4649 47296 4665 47360
rect 4729 47296 4737 47360
rect 4417 46272 4737 47296
rect 4417 46208 4425 46272
rect 4489 46208 4505 46272
rect 4569 46208 4585 46272
rect 4649 46208 4665 46272
rect 4729 46208 4737 46272
rect 4417 45184 4737 46208
rect 4417 45120 4425 45184
rect 4489 45120 4505 45184
rect 4569 45120 4585 45184
rect 4649 45120 4665 45184
rect 4729 45120 4737 45184
rect 4417 44096 4737 45120
rect 4417 44032 4425 44096
rect 4489 44032 4505 44096
rect 4569 44032 4585 44096
rect 4649 44032 4665 44096
rect 4729 44032 4737 44096
rect 4417 43008 4737 44032
rect 4417 42944 4425 43008
rect 4489 42944 4505 43008
rect 4569 42944 4585 43008
rect 4649 42944 4665 43008
rect 4729 42944 4737 43008
rect 4417 41920 4737 42944
rect 4417 41856 4425 41920
rect 4489 41856 4505 41920
rect 4569 41856 4585 41920
rect 4649 41856 4665 41920
rect 4729 41856 4737 41920
rect 4417 40832 4737 41856
rect 4417 40768 4425 40832
rect 4489 40768 4505 40832
rect 4569 40768 4585 40832
rect 4649 40768 4665 40832
rect 4729 40768 4737 40832
rect 4417 39744 4737 40768
rect 4417 39680 4425 39744
rect 4489 39680 4505 39744
rect 4569 39680 4585 39744
rect 4649 39680 4665 39744
rect 4729 39680 4737 39744
rect 4417 38656 4737 39680
rect 4417 38592 4425 38656
rect 4489 38592 4505 38656
rect 4569 38592 4585 38656
rect 4649 38592 4665 38656
rect 4729 38592 4737 38656
rect 4417 37568 4737 38592
rect 4417 37504 4425 37568
rect 4489 37504 4505 37568
rect 4569 37504 4585 37568
rect 4649 37504 4665 37568
rect 4729 37504 4737 37568
rect 4417 36480 4737 37504
rect 4417 36416 4425 36480
rect 4489 36416 4505 36480
rect 4569 36416 4585 36480
rect 4649 36416 4665 36480
rect 4729 36416 4737 36480
rect 4417 35392 4737 36416
rect 4417 35328 4425 35392
rect 4489 35328 4505 35392
rect 4569 35328 4585 35392
rect 4649 35328 4665 35392
rect 4729 35328 4737 35392
rect 4417 34304 4737 35328
rect 4417 34240 4425 34304
rect 4489 34240 4505 34304
rect 4569 34240 4585 34304
rect 4649 34240 4665 34304
rect 4729 34240 4737 34304
rect 4417 33216 4737 34240
rect 4417 33152 4425 33216
rect 4489 33152 4505 33216
rect 4569 33152 4585 33216
rect 4649 33152 4665 33216
rect 4729 33152 4737 33216
rect 4417 32128 4737 33152
rect 4417 32064 4425 32128
rect 4489 32064 4505 32128
rect 4569 32064 4585 32128
rect 4649 32064 4665 32128
rect 4729 32064 4737 32128
rect 4417 31040 4737 32064
rect 4417 30976 4425 31040
rect 4489 30976 4505 31040
rect 4569 30976 4585 31040
rect 4649 30976 4665 31040
rect 4729 30976 4737 31040
rect 4417 29952 4737 30976
rect 4417 29888 4425 29952
rect 4489 29888 4505 29952
rect 4569 29888 4585 29952
rect 4649 29888 4665 29952
rect 4729 29888 4737 29952
rect 4417 28864 4737 29888
rect 4417 28800 4425 28864
rect 4489 28800 4505 28864
rect 4569 28800 4585 28864
rect 4649 28800 4665 28864
rect 4729 28800 4737 28864
rect 4417 27776 4737 28800
rect 4417 27712 4425 27776
rect 4489 27712 4505 27776
rect 4569 27712 4585 27776
rect 4649 27712 4665 27776
rect 4729 27712 4737 27776
rect 4417 26688 4737 27712
rect 4417 26624 4425 26688
rect 4489 26624 4505 26688
rect 4569 26624 4585 26688
rect 4649 26624 4665 26688
rect 4729 26624 4737 26688
rect 4417 25600 4737 26624
rect 4417 25536 4425 25600
rect 4489 25536 4505 25600
rect 4569 25536 4585 25600
rect 4649 25536 4665 25600
rect 4729 25536 4737 25600
rect 4417 24512 4737 25536
rect 4417 24448 4425 24512
rect 4489 24448 4505 24512
rect 4569 24448 4585 24512
rect 4649 24448 4665 24512
rect 4729 24448 4737 24512
rect 4417 23424 4737 24448
rect 4417 23360 4425 23424
rect 4489 23360 4505 23424
rect 4569 23360 4585 23424
rect 4649 23360 4665 23424
rect 4729 23360 4737 23424
rect 4417 22336 4737 23360
rect 4417 22272 4425 22336
rect 4489 22272 4505 22336
rect 4569 22272 4585 22336
rect 4649 22272 4665 22336
rect 4729 22272 4737 22336
rect 4417 21248 4737 22272
rect 4417 21184 4425 21248
rect 4489 21184 4505 21248
rect 4569 21184 4585 21248
rect 4649 21184 4665 21248
rect 4729 21184 4737 21248
rect 4417 20160 4737 21184
rect 4417 20096 4425 20160
rect 4489 20096 4505 20160
rect 4569 20096 4585 20160
rect 4649 20096 4665 20160
rect 4729 20096 4737 20160
rect 4417 19072 4737 20096
rect 4417 19008 4425 19072
rect 4489 19008 4505 19072
rect 4569 19008 4585 19072
rect 4649 19008 4665 19072
rect 4729 19008 4737 19072
rect 4417 17984 4737 19008
rect 4417 17920 4425 17984
rect 4489 17920 4505 17984
rect 4569 17920 4585 17984
rect 4649 17920 4665 17984
rect 4729 17920 4737 17984
rect 4417 16896 4737 17920
rect 4417 16832 4425 16896
rect 4489 16832 4505 16896
rect 4569 16832 4585 16896
rect 4649 16832 4665 16896
rect 4729 16832 4737 16896
rect 4417 15808 4737 16832
rect 4417 15744 4425 15808
rect 4489 15744 4505 15808
rect 4569 15744 4585 15808
rect 4649 15744 4665 15808
rect 4729 15744 4737 15808
rect 4417 14720 4737 15744
rect 4417 14656 4425 14720
rect 4489 14656 4505 14720
rect 4569 14656 4585 14720
rect 4649 14656 4665 14720
rect 4729 14656 4737 14720
rect 4417 13632 4737 14656
rect 4417 13568 4425 13632
rect 4489 13568 4505 13632
rect 4569 13568 4585 13632
rect 4649 13568 4665 13632
rect 4729 13568 4737 13632
rect 4417 12544 4737 13568
rect 4417 12480 4425 12544
rect 4489 12480 4505 12544
rect 4569 12480 4585 12544
rect 4649 12480 4665 12544
rect 4729 12480 4737 12544
rect 4417 11456 4737 12480
rect 4417 11392 4425 11456
rect 4489 11392 4505 11456
rect 4569 11392 4585 11456
rect 4649 11392 4665 11456
rect 4729 11392 4737 11456
rect 4417 10368 4737 11392
rect 4417 10304 4425 10368
rect 4489 10304 4505 10368
rect 4569 10304 4585 10368
rect 4649 10304 4665 10368
rect 4729 10304 4737 10368
rect 4417 9280 4737 10304
rect 4417 9216 4425 9280
rect 4489 9216 4505 9280
rect 4569 9216 4585 9280
rect 4649 9216 4665 9280
rect 4729 9216 4737 9280
rect 4417 8192 4737 9216
rect 4417 8128 4425 8192
rect 4489 8128 4505 8192
rect 4569 8128 4585 8192
rect 4649 8128 4665 8192
rect 4729 8128 4737 8192
rect 4417 7104 4737 8128
rect 4417 7040 4425 7104
rect 4489 7040 4505 7104
rect 4569 7040 4585 7104
rect 4649 7040 4665 7104
rect 4729 7040 4737 7104
rect 4417 6016 4737 7040
rect 4417 5952 4425 6016
rect 4489 5952 4505 6016
rect 4569 5952 4585 6016
rect 4649 5952 4665 6016
rect 4729 5952 4737 6016
rect 4417 4928 4737 5952
rect 4417 4864 4425 4928
rect 4489 4864 4505 4928
rect 4569 4864 4585 4928
rect 4649 4864 4665 4928
rect 4729 4864 4737 4928
rect 4417 3840 4737 4864
rect 4417 3776 4425 3840
rect 4489 3776 4505 3840
rect 4569 3776 4585 3840
rect 4649 3776 4665 3840
rect 4729 3776 4737 3840
rect 4417 2752 4737 3776
rect 4417 2688 4425 2752
rect 4489 2688 4505 2752
rect 4569 2688 4585 2752
rect 4649 2688 4665 2752
rect 4729 2688 4737 2752
rect 4417 2128 4737 2688
rect 7890 46816 8210 47376
rect 7890 46752 7898 46816
rect 7962 46752 7978 46816
rect 8042 46752 8058 46816
rect 8122 46752 8138 46816
rect 8202 46752 8210 46816
rect 7890 45728 8210 46752
rect 7890 45664 7898 45728
rect 7962 45664 7978 45728
rect 8042 45664 8058 45728
rect 8122 45664 8138 45728
rect 8202 45664 8210 45728
rect 7890 44640 8210 45664
rect 7890 44576 7898 44640
rect 7962 44576 7978 44640
rect 8042 44576 8058 44640
rect 8122 44576 8138 44640
rect 8202 44576 8210 44640
rect 7890 43552 8210 44576
rect 7890 43488 7898 43552
rect 7962 43488 7978 43552
rect 8042 43488 8058 43552
rect 8122 43488 8138 43552
rect 8202 43488 8210 43552
rect 7890 42464 8210 43488
rect 7890 42400 7898 42464
rect 7962 42400 7978 42464
rect 8042 42400 8058 42464
rect 8122 42400 8138 42464
rect 8202 42400 8210 42464
rect 7890 41376 8210 42400
rect 7890 41312 7898 41376
rect 7962 41312 7978 41376
rect 8042 41312 8058 41376
rect 8122 41312 8138 41376
rect 8202 41312 8210 41376
rect 7890 40288 8210 41312
rect 7890 40224 7898 40288
rect 7962 40224 7978 40288
rect 8042 40224 8058 40288
rect 8122 40224 8138 40288
rect 8202 40224 8210 40288
rect 7890 39200 8210 40224
rect 7890 39136 7898 39200
rect 7962 39136 7978 39200
rect 8042 39136 8058 39200
rect 8122 39136 8138 39200
rect 8202 39136 8210 39200
rect 7890 38112 8210 39136
rect 7890 38048 7898 38112
rect 7962 38048 7978 38112
rect 8042 38048 8058 38112
rect 8122 38048 8138 38112
rect 8202 38048 8210 38112
rect 7890 37024 8210 38048
rect 7890 36960 7898 37024
rect 7962 36960 7978 37024
rect 8042 36960 8058 37024
rect 8122 36960 8138 37024
rect 8202 36960 8210 37024
rect 7890 35936 8210 36960
rect 7890 35872 7898 35936
rect 7962 35872 7978 35936
rect 8042 35872 8058 35936
rect 8122 35872 8138 35936
rect 8202 35872 8210 35936
rect 7890 34848 8210 35872
rect 7890 34784 7898 34848
rect 7962 34784 7978 34848
rect 8042 34784 8058 34848
rect 8122 34784 8138 34848
rect 8202 34784 8210 34848
rect 7890 33760 8210 34784
rect 7890 33696 7898 33760
rect 7962 33696 7978 33760
rect 8042 33696 8058 33760
rect 8122 33696 8138 33760
rect 8202 33696 8210 33760
rect 7890 32672 8210 33696
rect 7890 32608 7898 32672
rect 7962 32608 7978 32672
rect 8042 32608 8058 32672
rect 8122 32608 8138 32672
rect 8202 32608 8210 32672
rect 7890 31584 8210 32608
rect 7890 31520 7898 31584
rect 7962 31520 7978 31584
rect 8042 31520 8058 31584
rect 8122 31520 8138 31584
rect 8202 31520 8210 31584
rect 7890 30496 8210 31520
rect 7890 30432 7898 30496
rect 7962 30432 7978 30496
rect 8042 30432 8058 30496
rect 8122 30432 8138 30496
rect 8202 30432 8210 30496
rect 7890 29408 8210 30432
rect 7890 29344 7898 29408
rect 7962 29344 7978 29408
rect 8042 29344 8058 29408
rect 8122 29344 8138 29408
rect 8202 29344 8210 29408
rect 7890 28320 8210 29344
rect 7890 28256 7898 28320
rect 7962 28256 7978 28320
rect 8042 28256 8058 28320
rect 8122 28256 8138 28320
rect 8202 28256 8210 28320
rect 7890 27232 8210 28256
rect 7890 27168 7898 27232
rect 7962 27168 7978 27232
rect 8042 27168 8058 27232
rect 8122 27168 8138 27232
rect 8202 27168 8210 27232
rect 7890 26144 8210 27168
rect 7890 26080 7898 26144
rect 7962 26080 7978 26144
rect 8042 26080 8058 26144
rect 8122 26080 8138 26144
rect 8202 26080 8210 26144
rect 7890 25056 8210 26080
rect 7890 24992 7898 25056
rect 7962 24992 7978 25056
rect 8042 24992 8058 25056
rect 8122 24992 8138 25056
rect 8202 24992 8210 25056
rect 7890 23968 8210 24992
rect 7890 23904 7898 23968
rect 7962 23904 7978 23968
rect 8042 23904 8058 23968
rect 8122 23904 8138 23968
rect 8202 23904 8210 23968
rect 7890 22880 8210 23904
rect 7890 22816 7898 22880
rect 7962 22816 7978 22880
rect 8042 22816 8058 22880
rect 8122 22816 8138 22880
rect 8202 22816 8210 22880
rect 7890 21792 8210 22816
rect 7890 21728 7898 21792
rect 7962 21728 7978 21792
rect 8042 21728 8058 21792
rect 8122 21728 8138 21792
rect 8202 21728 8210 21792
rect 7890 20704 8210 21728
rect 7890 20640 7898 20704
rect 7962 20640 7978 20704
rect 8042 20640 8058 20704
rect 8122 20640 8138 20704
rect 8202 20640 8210 20704
rect 7890 19616 8210 20640
rect 7890 19552 7898 19616
rect 7962 19552 7978 19616
rect 8042 19552 8058 19616
rect 8122 19552 8138 19616
rect 8202 19552 8210 19616
rect 7890 18528 8210 19552
rect 7890 18464 7898 18528
rect 7962 18464 7978 18528
rect 8042 18464 8058 18528
rect 8122 18464 8138 18528
rect 8202 18464 8210 18528
rect 7890 17440 8210 18464
rect 7890 17376 7898 17440
rect 7962 17376 7978 17440
rect 8042 17376 8058 17440
rect 8122 17376 8138 17440
rect 8202 17376 8210 17440
rect 7890 16352 8210 17376
rect 7890 16288 7898 16352
rect 7962 16288 7978 16352
rect 8042 16288 8058 16352
rect 8122 16288 8138 16352
rect 8202 16288 8210 16352
rect 7890 15264 8210 16288
rect 7890 15200 7898 15264
rect 7962 15200 7978 15264
rect 8042 15200 8058 15264
rect 8122 15200 8138 15264
rect 8202 15200 8210 15264
rect 7890 14176 8210 15200
rect 7890 14112 7898 14176
rect 7962 14112 7978 14176
rect 8042 14112 8058 14176
rect 8122 14112 8138 14176
rect 8202 14112 8210 14176
rect 7890 13088 8210 14112
rect 7890 13024 7898 13088
rect 7962 13024 7978 13088
rect 8042 13024 8058 13088
rect 8122 13024 8138 13088
rect 8202 13024 8210 13088
rect 7890 12000 8210 13024
rect 7890 11936 7898 12000
rect 7962 11936 7978 12000
rect 8042 11936 8058 12000
rect 8122 11936 8138 12000
rect 8202 11936 8210 12000
rect 7890 10912 8210 11936
rect 7890 10848 7898 10912
rect 7962 10848 7978 10912
rect 8042 10848 8058 10912
rect 8122 10848 8138 10912
rect 8202 10848 8210 10912
rect 7890 9824 8210 10848
rect 7890 9760 7898 9824
rect 7962 9760 7978 9824
rect 8042 9760 8058 9824
rect 8122 9760 8138 9824
rect 8202 9760 8210 9824
rect 7890 8736 8210 9760
rect 7890 8672 7898 8736
rect 7962 8672 7978 8736
rect 8042 8672 8058 8736
rect 8122 8672 8138 8736
rect 8202 8672 8210 8736
rect 7890 7648 8210 8672
rect 7890 7584 7898 7648
rect 7962 7584 7978 7648
rect 8042 7584 8058 7648
rect 8122 7584 8138 7648
rect 8202 7584 8210 7648
rect 7890 6560 8210 7584
rect 7890 6496 7898 6560
rect 7962 6496 7978 6560
rect 8042 6496 8058 6560
rect 8122 6496 8138 6560
rect 8202 6496 8210 6560
rect 7890 5472 8210 6496
rect 7890 5408 7898 5472
rect 7962 5408 7978 5472
rect 8042 5408 8058 5472
rect 8122 5408 8138 5472
rect 8202 5408 8210 5472
rect 7890 4384 8210 5408
rect 7890 4320 7898 4384
rect 7962 4320 7978 4384
rect 8042 4320 8058 4384
rect 8122 4320 8138 4384
rect 8202 4320 8210 4384
rect 7890 3296 8210 4320
rect 7890 3232 7898 3296
rect 7962 3232 7978 3296
rect 8042 3232 8058 3296
rect 8122 3232 8138 3296
rect 8202 3232 8210 3296
rect 7890 2208 8210 3232
rect 7890 2144 7898 2208
rect 7962 2144 7978 2208
rect 8042 2144 8058 2208
rect 8122 2144 8138 2208
rect 8202 2144 8210 2208
rect 7890 2128 8210 2144
rect 11363 47360 11683 47376
rect 11363 47296 11371 47360
rect 11435 47296 11451 47360
rect 11515 47296 11531 47360
rect 11595 47296 11611 47360
rect 11675 47296 11683 47360
rect 11363 46272 11683 47296
rect 11363 46208 11371 46272
rect 11435 46208 11451 46272
rect 11515 46208 11531 46272
rect 11595 46208 11611 46272
rect 11675 46208 11683 46272
rect 11363 45184 11683 46208
rect 11363 45120 11371 45184
rect 11435 45120 11451 45184
rect 11515 45120 11531 45184
rect 11595 45120 11611 45184
rect 11675 45120 11683 45184
rect 11363 44096 11683 45120
rect 11363 44032 11371 44096
rect 11435 44032 11451 44096
rect 11515 44032 11531 44096
rect 11595 44032 11611 44096
rect 11675 44032 11683 44096
rect 11363 43008 11683 44032
rect 11363 42944 11371 43008
rect 11435 42944 11451 43008
rect 11515 42944 11531 43008
rect 11595 42944 11611 43008
rect 11675 42944 11683 43008
rect 11363 41920 11683 42944
rect 11363 41856 11371 41920
rect 11435 41856 11451 41920
rect 11515 41856 11531 41920
rect 11595 41856 11611 41920
rect 11675 41856 11683 41920
rect 11363 40832 11683 41856
rect 11363 40768 11371 40832
rect 11435 40768 11451 40832
rect 11515 40768 11531 40832
rect 11595 40768 11611 40832
rect 11675 40768 11683 40832
rect 11363 39744 11683 40768
rect 11363 39680 11371 39744
rect 11435 39680 11451 39744
rect 11515 39680 11531 39744
rect 11595 39680 11611 39744
rect 11675 39680 11683 39744
rect 11363 38656 11683 39680
rect 11363 38592 11371 38656
rect 11435 38592 11451 38656
rect 11515 38592 11531 38656
rect 11595 38592 11611 38656
rect 11675 38592 11683 38656
rect 11363 37568 11683 38592
rect 11363 37504 11371 37568
rect 11435 37504 11451 37568
rect 11515 37504 11531 37568
rect 11595 37504 11611 37568
rect 11675 37504 11683 37568
rect 11363 36480 11683 37504
rect 11363 36416 11371 36480
rect 11435 36416 11451 36480
rect 11515 36416 11531 36480
rect 11595 36416 11611 36480
rect 11675 36416 11683 36480
rect 11363 35392 11683 36416
rect 11363 35328 11371 35392
rect 11435 35328 11451 35392
rect 11515 35328 11531 35392
rect 11595 35328 11611 35392
rect 11675 35328 11683 35392
rect 11363 34304 11683 35328
rect 11363 34240 11371 34304
rect 11435 34240 11451 34304
rect 11515 34240 11531 34304
rect 11595 34240 11611 34304
rect 11675 34240 11683 34304
rect 11363 33216 11683 34240
rect 11363 33152 11371 33216
rect 11435 33152 11451 33216
rect 11515 33152 11531 33216
rect 11595 33152 11611 33216
rect 11675 33152 11683 33216
rect 11363 32128 11683 33152
rect 11363 32064 11371 32128
rect 11435 32064 11451 32128
rect 11515 32064 11531 32128
rect 11595 32064 11611 32128
rect 11675 32064 11683 32128
rect 11363 31040 11683 32064
rect 11363 30976 11371 31040
rect 11435 30976 11451 31040
rect 11515 30976 11531 31040
rect 11595 30976 11611 31040
rect 11675 30976 11683 31040
rect 11363 29952 11683 30976
rect 11363 29888 11371 29952
rect 11435 29888 11451 29952
rect 11515 29888 11531 29952
rect 11595 29888 11611 29952
rect 11675 29888 11683 29952
rect 11363 28864 11683 29888
rect 11363 28800 11371 28864
rect 11435 28800 11451 28864
rect 11515 28800 11531 28864
rect 11595 28800 11611 28864
rect 11675 28800 11683 28864
rect 11363 27776 11683 28800
rect 11363 27712 11371 27776
rect 11435 27712 11451 27776
rect 11515 27712 11531 27776
rect 11595 27712 11611 27776
rect 11675 27712 11683 27776
rect 11363 26688 11683 27712
rect 11363 26624 11371 26688
rect 11435 26624 11451 26688
rect 11515 26624 11531 26688
rect 11595 26624 11611 26688
rect 11675 26624 11683 26688
rect 11363 25600 11683 26624
rect 11363 25536 11371 25600
rect 11435 25536 11451 25600
rect 11515 25536 11531 25600
rect 11595 25536 11611 25600
rect 11675 25536 11683 25600
rect 11363 24512 11683 25536
rect 11363 24448 11371 24512
rect 11435 24448 11451 24512
rect 11515 24448 11531 24512
rect 11595 24448 11611 24512
rect 11675 24448 11683 24512
rect 11363 23424 11683 24448
rect 11363 23360 11371 23424
rect 11435 23360 11451 23424
rect 11515 23360 11531 23424
rect 11595 23360 11611 23424
rect 11675 23360 11683 23424
rect 11363 22336 11683 23360
rect 11363 22272 11371 22336
rect 11435 22272 11451 22336
rect 11515 22272 11531 22336
rect 11595 22272 11611 22336
rect 11675 22272 11683 22336
rect 11363 21248 11683 22272
rect 11363 21184 11371 21248
rect 11435 21184 11451 21248
rect 11515 21184 11531 21248
rect 11595 21184 11611 21248
rect 11675 21184 11683 21248
rect 11363 20160 11683 21184
rect 11363 20096 11371 20160
rect 11435 20096 11451 20160
rect 11515 20096 11531 20160
rect 11595 20096 11611 20160
rect 11675 20096 11683 20160
rect 11363 19072 11683 20096
rect 11363 19008 11371 19072
rect 11435 19008 11451 19072
rect 11515 19008 11531 19072
rect 11595 19008 11611 19072
rect 11675 19008 11683 19072
rect 11363 17984 11683 19008
rect 11363 17920 11371 17984
rect 11435 17920 11451 17984
rect 11515 17920 11531 17984
rect 11595 17920 11611 17984
rect 11675 17920 11683 17984
rect 11363 16896 11683 17920
rect 11363 16832 11371 16896
rect 11435 16832 11451 16896
rect 11515 16832 11531 16896
rect 11595 16832 11611 16896
rect 11675 16832 11683 16896
rect 11363 15808 11683 16832
rect 11363 15744 11371 15808
rect 11435 15744 11451 15808
rect 11515 15744 11531 15808
rect 11595 15744 11611 15808
rect 11675 15744 11683 15808
rect 11363 14720 11683 15744
rect 11363 14656 11371 14720
rect 11435 14656 11451 14720
rect 11515 14656 11531 14720
rect 11595 14656 11611 14720
rect 11675 14656 11683 14720
rect 11363 13632 11683 14656
rect 11363 13568 11371 13632
rect 11435 13568 11451 13632
rect 11515 13568 11531 13632
rect 11595 13568 11611 13632
rect 11675 13568 11683 13632
rect 11363 12544 11683 13568
rect 11363 12480 11371 12544
rect 11435 12480 11451 12544
rect 11515 12480 11531 12544
rect 11595 12480 11611 12544
rect 11675 12480 11683 12544
rect 11363 11456 11683 12480
rect 11363 11392 11371 11456
rect 11435 11392 11451 11456
rect 11515 11392 11531 11456
rect 11595 11392 11611 11456
rect 11675 11392 11683 11456
rect 11363 10368 11683 11392
rect 11363 10304 11371 10368
rect 11435 10304 11451 10368
rect 11515 10304 11531 10368
rect 11595 10304 11611 10368
rect 11675 10304 11683 10368
rect 11363 9280 11683 10304
rect 11363 9216 11371 9280
rect 11435 9216 11451 9280
rect 11515 9216 11531 9280
rect 11595 9216 11611 9280
rect 11675 9216 11683 9280
rect 11363 8192 11683 9216
rect 11363 8128 11371 8192
rect 11435 8128 11451 8192
rect 11515 8128 11531 8192
rect 11595 8128 11611 8192
rect 11675 8128 11683 8192
rect 11363 7104 11683 8128
rect 11363 7040 11371 7104
rect 11435 7040 11451 7104
rect 11515 7040 11531 7104
rect 11595 7040 11611 7104
rect 11675 7040 11683 7104
rect 11363 6016 11683 7040
rect 11363 5952 11371 6016
rect 11435 5952 11451 6016
rect 11515 5952 11531 6016
rect 11595 5952 11611 6016
rect 11675 5952 11683 6016
rect 11363 4928 11683 5952
rect 11363 4864 11371 4928
rect 11435 4864 11451 4928
rect 11515 4864 11531 4928
rect 11595 4864 11611 4928
rect 11675 4864 11683 4928
rect 11363 3840 11683 4864
rect 11363 3776 11371 3840
rect 11435 3776 11451 3840
rect 11515 3776 11531 3840
rect 11595 3776 11611 3840
rect 11675 3776 11683 3840
rect 11363 2752 11683 3776
rect 11363 2688 11371 2752
rect 11435 2688 11451 2752
rect 11515 2688 11531 2752
rect 11595 2688 11611 2752
rect 11675 2688 11683 2752
rect 11363 2128 11683 2688
rect 14836 46816 15156 47376
rect 14836 46752 14844 46816
rect 14908 46752 14924 46816
rect 14988 46752 15004 46816
rect 15068 46752 15084 46816
rect 15148 46752 15156 46816
rect 14836 45728 15156 46752
rect 14836 45664 14844 45728
rect 14908 45664 14924 45728
rect 14988 45664 15004 45728
rect 15068 45664 15084 45728
rect 15148 45664 15156 45728
rect 14836 44640 15156 45664
rect 14836 44576 14844 44640
rect 14908 44576 14924 44640
rect 14988 44576 15004 44640
rect 15068 44576 15084 44640
rect 15148 44576 15156 44640
rect 14836 43552 15156 44576
rect 14836 43488 14844 43552
rect 14908 43488 14924 43552
rect 14988 43488 15004 43552
rect 15068 43488 15084 43552
rect 15148 43488 15156 43552
rect 14836 42464 15156 43488
rect 14836 42400 14844 42464
rect 14908 42400 14924 42464
rect 14988 42400 15004 42464
rect 15068 42400 15084 42464
rect 15148 42400 15156 42464
rect 14836 41376 15156 42400
rect 14836 41312 14844 41376
rect 14908 41312 14924 41376
rect 14988 41312 15004 41376
rect 15068 41312 15084 41376
rect 15148 41312 15156 41376
rect 14836 40288 15156 41312
rect 14836 40224 14844 40288
rect 14908 40224 14924 40288
rect 14988 40224 15004 40288
rect 15068 40224 15084 40288
rect 15148 40224 15156 40288
rect 14836 39200 15156 40224
rect 14836 39136 14844 39200
rect 14908 39136 14924 39200
rect 14988 39136 15004 39200
rect 15068 39136 15084 39200
rect 15148 39136 15156 39200
rect 14836 38112 15156 39136
rect 14836 38048 14844 38112
rect 14908 38048 14924 38112
rect 14988 38048 15004 38112
rect 15068 38048 15084 38112
rect 15148 38048 15156 38112
rect 14836 37024 15156 38048
rect 14836 36960 14844 37024
rect 14908 36960 14924 37024
rect 14988 36960 15004 37024
rect 15068 36960 15084 37024
rect 15148 36960 15156 37024
rect 14836 35936 15156 36960
rect 14836 35872 14844 35936
rect 14908 35872 14924 35936
rect 14988 35872 15004 35936
rect 15068 35872 15084 35936
rect 15148 35872 15156 35936
rect 14836 34848 15156 35872
rect 14836 34784 14844 34848
rect 14908 34784 14924 34848
rect 14988 34784 15004 34848
rect 15068 34784 15084 34848
rect 15148 34784 15156 34848
rect 14836 33760 15156 34784
rect 14836 33696 14844 33760
rect 14908 33696 14924 33760
rect 14988 33696 15004 33760
rect 15068 33696 15084 33760
rect 15148 33696 15156 33760
rect 14836 32672 15156 33696
rect 14836 32608 14844 32672
rect 14908 32608 14924 32672
rect 14988 32608 15004 32672
rect 15068 32608 15084 32672
rect 15148 32608 15156 32672
rect 14836 31584 15156 32608
rect 14836 31520 14844 31584
rect 14908 31520 14924 31584
rect 14988 31520 15004 31584
rect 15068 31520 15084 31584
rect 15148 31520 15156 31584
rect 14836 30496 15156 31520
rect 14836 30432 14844 30496
rect 14908 30432 14924 30496
rect 14988 30432 15004 30496
rect 15068 30432 15084 30496
rect 15148 30432 15156 30496
rect 14836 29408 15156 30432
rect 14836 29344 14844 29408
rect 14908 29344 14924 29408
rect 14988 29344 15004 29408
rect 15068 29344 15084 29408
rect 15148 29344 15156 29408
rect 14836 28320 15156 29344
rect 14836 28256 14844 28320
rect 14908 28256 14924 28320
rect 14988 28256 15004 28320
rect 15068 28256 15084 28320
rect 15148 28256 15156 28320
rect 14836 27232 15156 28256
rect 14836 27168 14844 27232
rect 14908 27168 14924 27232
rect 14988 27168 15004 27232
rect 15068 27168 15084 27232
rect 15148 27168 15156 27232
rect 14836 26144 15156 27168
rect 14836 26080 14844 26144
rect 14908 26080 14924 26144
rect 14988 26080 15004 26144
rect 15068 26080 15084 26144
rect 15148 26080 15156 26144
rect 14836 25056 15156 26080
rect 14836 24992 14844 25056
rect 14908 24992 14924 25056
rect 14988 24992 15004 25056
rect 15068 24992 15084 25056
rect 15148 24992 15156 25056
rect 14836 23968 15156 24992
rect 14836 23904 14844 23968
rect 14908 23904 14924 23968
rect 14988 23904 15004 23968
rect 15068 23904 15084 23968
rect 15148 23904 15156 23968
rect 14836 22880 15156 23904
rect 14836 22816 14844 22880
rect 14908 22816 14924 22880
rect 14988 22816 15004 22880
rect 15068 22816 15084 22880
rect 15148 22816 15156 22880
rect 14836 21792 15156 22816
rect 14836 21728 14844 21792
rect 14908 21728 14924 21792
rect 14988 21728 15004 21792
rect 15068 21728 15084 21792
rect 15148 21728 15156 21792
rect 14836 20704 15156 21728
rect 14836 20640 14844 20704
rect 14908 20640 14924 20704
rect 14988 20640 15004 20704
rect 15068 20640 15084 20704
rect 15148 20640 15156 20704
rect 14836 19616 15156 20640
rect 14836 19552 14844 19616
rect 14908 19552 14924 19616
rect 14988 19552 15004 19616
rect 15068 19552 15084 19616
rect 15148 19552 15156 19616
rect 14836 18528 15156 19552
rect 14836 18464 14844 18528
rect 14908 18464 14924 18528
rect 14988 18464 15004 18528
rect 15068 18464 15084 18528
rect 15148 18464 15156 18528
rect 14836 17440 15156 18464
rect 14836 17376 14844 17440
rect 14908 17376 14924 17440
rect 14988 17376 15004 17440
rect 15068 17376 15084 17440
rect 15148 17376 15156 17440
rect 14836 16352 15156 17376
rect 14836 16288 14844 16352
rect 14908 16288 14924 16352
rect 14988 16288 15004 16352
rect 15068 16288 15084 16352
rect 15148 16288 15156 16352
rect 14836 15264 15156 16288
rect 14836 15200 14844 15264
rect 14908 15200 14924 15264
rect 14988 15200 15004 15264
rect 15068 15200 15084 15264
rect 15148 15200 15156 15264
rect 14836 14176 15156 15200
rect 14836 14112 14844 14176
rect 14908 14112 14924 14176
rect 14988 14112 15004 14176
rect 15068 14112 15084 14176
rect 15148 14112 15156 14176
rect 14836 13088 15156 14112
rect 14836 13024 14844 13088
rect 14908 13024 14924 13088
rect 14988 13024 15004 13088
rect 15068 13024 15084 13088
rect 15148 13024 15156 13088
rect 14836 12000 15156 13024
rect 14836 11936 14844 12000
rect 14908 11936 14924 12000
rect 14988 11936 15004 12000
rect 15068 11936 15084 12000
rect 15148 11936 15156 12000
rect 14836 10912 15156 11936
rect 14836 10848 14844 10912
rect 14908 10848 14924 10912
rect 14988 10848 15004 10912
rect 15068 10848 15084 10912
rect 15148 10848 15156 10912
rect 14836 9824 15156 10848
rect 14836 9760 14844 9824
rect 14908 9760 14924 9824
rect 14988 9760 15004 9824
rect 15068 9760 15084 9824
rect 15148 9760 15156 9824
rect 14836 8736 15156 9760
rect 14836 8672 14844 8736
rect 14908 8672 14924 8736
rect 14988 8672 15004 8736
rect 15068 8672 15084 8736
rect 15148 8672 15156 8736
rect 14836 7648 15156 8672
rect 14836 7584 14844 7648
rect 14908 7584 14924 7648
rect 14988 7584 15004 7648
rect 15068 7584 15084 7648
rect 15148 7584 15156 7648
rect 14836 6560 15156 7584
rect 14836 6496 14844 6560
rect 14908 6496 14924 6560
rect 14988 6496 15004 6560
rect 15068 6496 15084 6560
rect 15148 6496 15156 6560
rect 14836 5472 15156 6496
rect 14836 5408 14844 5472
rect 14908 5408 14924 5472
rect 14988 5408 15004 5472
rect 15068 5408 15084 5472
rect 15148 5408 15156 5472
rect 14836 4384 15156 5408
rect 14836 4320 14844 4384
rect 14908 4320 14924 4384
rect 14988 4320 15004 4384
rect 15068 4320 15084 4384
rect 15148 4320 15156 4384
rect 14836 3296 15156 4320
rect 14836 3232 14844 3296
rect 14908 3232 14924 3296
rect 14988 3232 15004 3296
rect 15068 3232 15084 3296
rect 15148 3232 15156 3296
rect 14836 2208 15156 3232
rect 14836 2144 14844 2208
rect 14908 2144 14924 2208
rect 14988 2144 15004 2208
rect 15068 2144 15084 2208
rect 15148 2144 15156 2208
rect 14836 2128 15156 2144
rect 18309 47360 18629 47376
rect 18309 47296 18317 47360
rect 18381 47296 18397 47360
rect 18461 47296 18477 47360
rect 18541 47296 18557 47360
rect 18621 47296 18629 47360
rect 18309 46272 18629 47296
rect 18309 46208 18317 46272
rect 18381 46208 18397 46272
rect 18461 46208 18477 46272
rect 18541 46208 18557 46272
rect 18621 46208 18629 46272
rect 18309 45184 18629 46208
rect 18309 45120 18317 45184
rect 18381 45120 18397 45184
rect 18461 45120 18477 45184
rect 18541 45120 18557 45184
rect 18621 45120 18629 45184
rect 18309 44096 18629 45120
rect 18309 44032 18317 44096
rect 18381 44032 18397 44096
rect 18461 44032 18477 44096
rect 18541 44032 18557 44096
rect 18621 44032 18629 44096
rect 18309 43008 18629 44032
rect 18309 42944 18317 43008
rect 18381 42944 18397 43008
rect 18461 42944 18477 43008
rect 18541 42944 18557 43008
rect 18621 42944 18629 43008
rect 18309 41920 18629 42944
rect 21782 46816 22102 47376
rect 21782 46752 21790 46816
rect 21854 46752 21870 46816
rect 21934 46752 21950 46816
rect 22014 46752 22030 46816
rect 22094 46752 22102 46816
rect 21782 45728 22102 46752
rect 21782 45664 21790 45728
rect 21854 45664 21870 45728
rect 21934 45664 21950 45728
rect 22014 45664 22030 45728
rect 22094 45664 22102 45728
rect 21782 44640 22102 45664
rect 21782 44576 21790 44640
rect 21854 44576 21870 44640
rect 21934 44576 21950 44640
rect 22014 44576 22030 44640
rect 22094 44576 22102 44640
rect 21782 43552 22102 44576
rect 21782 43488 21790 43552
rect 21854 43488 21870 43552
rect 21934 43488 21950 43552
rect 22014 43488 22030 43552
rect 22094 43488 22102 43552
rect 19563 42940 19629 42941
rect 19563 42876 19564 42940
rect 19628 42876 19629 42940
rect 19563 42875 19629 42876
rect 18309 41856 18317 41920
rect 18381 41856 18397 41920
rect 18461 41856 18477 41920
rect 18541 41856 18557 41920
rect 18621 41856 18629 41920
rect 18309 40832 18629 41856
rect 18309 40768 18317 40832
rect 18381 40768 18397 40832
rect 18461 40768 18477 40832
rect 18541 40768 18557 40832
rect 18621 40768 18629 40832
rect 18309 39744 18629 40768
rect 18309 39680 18317 39744
rect 18381 39680 18397 39744
rect 18461 39680 18477 39744
rect 18541 39680 18557 39744
rect 18621 39680 18629 39744
rect 18309 38656 18629 39680
rect 18309 38592 18317 38656
rect 18381 38592 18397 38656
rect 18461 38592 18477 38656
rect 18541 38592 18557 38656
rect 18621 38592 18629 38656
rect 18309 37568 18629 38592
rect 18309 37504 18317 37568
rect 18381 37504 18397 37568
rect 18461 37504 18477 37568
rect 18541 37504 18557 37568
rect 18621 37504 18629 37568
rect 18309 36480 18629 37504
rect 18309 36416 18317 36480
rect 18381 36416 18397 36480
rect 18461 36416 18477 36480
rect 18541 36416 18557 36480
rect 18621 36416 18629 36480
rect 18309 35392 18629 36416
rect 18309 35328 18317 35392
rect 18381 35328 18397 35392
rect 18461 35328 18477 35392
rect 18541 35328 18557 35392
rect 18621 35328 18629 35392
rect 18309 34304 18629 35328
rect 18309 34240 18317 34304
rect 18381 34240 18397 34304
rect 18461 34240 18477 34304
rect 18541 34240 18557 34304
rect 18621 34240 18629 34304
rect 18309 33216 18629 34240
rect 18309 33152 18317 33216
rect 18381 33152 18397 33216
rect 18461 33152 18477 33216
rect 18541 33152 18557 33216
rect 18621 33152 18629 33216
rect 18309 32128 18629 33152
rect 18309 32064 18317 32128
rect 18381 32064 18397 32128
rect 18461 32064 18477 32128
rect 18541 32064 18557 32128
rect 18621 32064 18629 32128
rect 18309 31040 18629 32064
rect 18309 30976 18317 31040
rect 18381 30976 18397 31040
rect 18461 30976 18477 31040
rect 18541 30976 18557 31040
rect 18621 30976 18629 31040
rect 18309 29952 18629 30976
rect 18309 29888 18317 29952
rect 18381 29888 18397 29952
rect 18461 29888 18477 29952
rect 18541 29888 18557 29952
rect 18621 29888 18629 29952
rect 18309 28864 18629 29888
rect 18309 28800 18317 28864
rect 18381 28800 18397 28864
rect 18461 28800 18477 28864
rect 18541 28800 18557 28864
rect 18621 28800 18629 28864
rect 18309 27776 18629 28800
rect 18309 27712 18317 27776
rect 18381 27712 18397 27776
rect 18461 27712 18477 27776
rect 18541 27712 18557 27776
rect 18621 27712 18629 27776
rect 18309 26688 18629 27712
rect 18309 26624 18317 26688
rect 18381 26624 18397 26688
rect 18461 26624 18477 26688
rect 18541 26624 18557 26688
rect 18621 26624 18629 26688
rect 18309 25600 18629 26624
rect 18309 25536 18317 25600
rect 18381 25536 18397 25600
rect 18461 25536 18477 25600
rect 18541 25536 18557 25600
rect 18621 25536 18629 25600
rect 18309 24512 18629 25536
rect 19566 24717 19626 42875
rect 21782 42464 22102 43488
rect 21782 42400 21790 42464
rect 21854 42400 21870 42464
rect 21934 42400 21950 42464
rect 22014 42400 22030 42464
rect 22094 42400 22102 42464
rect 21782 41376 22102 42400
rect 21782 41312 21790 41376
rect 21854 41312 21870 41376
rect 21934 41312 21950 41376
rect 22014 41312 22030 41376
rect 22094 41312 22102 41376
rect 21782 40288 22102 41312
rect 21782 40224 21790 40288
rect 21854 40224 21870 40288
rect 21934 40224 21950 40288
rect 22014 40224 22030 40288
rect 22094 40224 22102 40288
rect 21782 39200 22102 40224
rect 21782 39136 21790 39200
rect 21854 39136 21870 39200
rect 21934 39136 21950 39200
rect 22014 39136 22030 39200
rect 22094 39136 22102 39200
rect 21782 38112 22102 39136
rect 21782 38048 21790 38112
rect 21854 38048 21870 38112
rect 21934 38048 21950 38112
rect 22014 38048 22030 38112
rect 22094 38048 22102 38112
rect 21782 37024 22102 38048
rect 21782 36960 21790 37024
rect 21854 36960 21870 37024
rect 21934 36960 21950 37024
rect 22014 36960 22030 37024
rect 22094 36960 22102 37024
rect 21782 35936 22102 36960
rect 21782 35872 21790 35936
rect 21854 35872 21870 35936
rect 21934 35872 21950 35936
rect 22014 35872 22030 35936
rect 22094 35872 22102 35936
rect 21782 34848 22102 35872
rect 21782 34784 21790 34848
rect 21854 34784 21870 34848
rect 21934 34784 21950 34848
rect 22014 34784 22030 34848
rect 22094 34784 22102 34848
rect 21782 33760 22102 34784
rect 21782 33696 21790 33760
rect 21854 33696 21870 33760
rect 21934 33696 21950 33760
rect 22014 33696 22030 33760
rect 22094 33696 22102 33760
rect 21782 32672 22102 33696
rect 21782 32608 21790 32672
rect 21854 32608 21870 32672
rect 21934 32608 21950 32672
rect 22014 32608 22030 32672
rect 22094 32608 22102 32672
rect 21782 31584 22102 32608
rect 21782 31520 21790 31584
rect 21854 31520 21870 31584
rect 21934 31520 21950 31584
rect 22014 31520 22030 31584
rect 22094 31520 22102 31584
rect 21782 30496 22102 31520
rect 21782 30432 21790 30496
rect 21854 30432 21870 30496
rect 21934 30432 21950 30496
rect 22014 30432 22030 30496
rect 22094 30432 22102 30496
rect 21782 29408 22102 30432
rect 21782 29344 21790 29408
rect 21854 29344 21870 29408
rect 21934 29344 21950 29408
rect 22014 29344 22030 29408
rect 22094 29344 22102 29408
rect 21782 28320 22102 29344
rect 21782 28256 21790 28320
rect 21854 28256 21870 28320
rect 21934 28256 21950 28320
rect 22014 28256 22030 28320
rect 22094 28256 22102 28320
rect 21782 27232 22102 28256
rect 21782 27168 21790 27232
rect 21854 27168 21870 27232
rect 21934 27168 21950 27232
rect 22014 27168 22030 27232
rect 22094 27168 22102 27232
rect 21782 26144 22102 27168
rect 21782 26080 21790 26144
rect 21854 26080 21870 26144
rect 21934 26080 21950 26144
rect 22014 26080 22030 26144
rect 22094 26080 22102 26144
rect 21782 25056 22102 26080
rect 21782 24992 21790 25056
rect 21854 24992 21870 25056
rect 21934 24992 21950 25056
rect 22014 24992 22030 25056
rect 22094 24992 22102 25056
rect 19563 24716 19629 24717
rect 19563 24652 19564 24716
rect 19628 24652 19629 24716
rect 19563 24651 19629 24652
rect 18309 24448 18317 24512
rect 18381 24448 18397 24512
rect 18461 24448 18477 24512
rect 18541 24448 18557 24512
rect 18621 24448 18629 24512
rect 18309 23424 18629 24448
rect 18309 23360 18317 23424
rect 18381 23360 18397 23424
rect 18461 23360 18477 23424
rect 18541 23360 18557 23424
rect 18621 23360 18629 23424
rect 18309 22336 18629 23360
rect 18309 22272 18317 22336
rect 18381 22272 18397 22336
rect 18461 22272 18477 22336
rect 18541 22272 18557 22336
rect 18621 22272 18629 22336
rect 18309 21248 18629 22272
rect 18309 21184 18317 21248
rect 18381 21184 18397 21248
rect 18461 21184 18477 21248
rect 18541 21184 18557 21248
rect 18621 21184 18629 21248
rect 18309 20160 18629 21184
rect 18309 20096 18317 20160
rect 18381 20096 18397 20160
rect 18461 20096 18477 20160
rect 18541 20096 18557 20160
rect 18621 20096 18629 20160
rect 18309 19072 18629 20096
rect 18309 19008 18317 19072
rect 18381 19008 18397 19072
rect 18461 19008 18477 19072
rect 18541 19008 18557 19072
rect 18621 19008 18629 19072
rect 18309 17984 18629 19008
rect 18309 17920 18317 17984
rect 18381 17920 18397 17984
rect 18461 17920 18477 17984
rect 18541 17920 18557 17984
rect 18621 17920 18629 17984
rect 18309 16896 18629 17920
rect 18309 16832 18317 16896
rect 18381 16832 18397 16896
rect 18461 16832 18477 16896
rect 18541 16832 18557 16896
rect 18621 16832 18629 16896
rect 18309 15808 18629 16832
rect 18309 15744 18317 15808
rect 18381 15744 18397 15808
rect 18461 15744 18477 15808
rect 18541 15744 18557 15808
rect 18621 15744 18629 15808
rect 18309 14720 18629 15744
rect 18309 14656 18317 14720
rect 18381 14656 18397 14720
rect 18461 14656 18477 14720
rect 18541 14656 18557 14720
rect 18621 14656 18629 14720
rect 18309 13632 18629 14656
rect 18309 13568 18317 13632
rect 18381 13568 18397 13632
rect 18461 13568 18477 13632
rect 18541 13568 18557 13632
rect 18621 13568 18629 13632
rect 18309 12544 18629 13568
rect 18309 12480 18317 12544
rect 18381 12480 18397 12544
rect 18461 12480 18477 12544
rect 18541 12480 18557 12544
rect 18621 12480 18629 12544
rect 18309 11456 18629 12480
rect 18309 11392 18317 11456
rect 18381 11392 18397 11456
rect 18461 11392 18477 11456
rect 18541 11392 18557 11456
rect 18621 11392 18629 11456
rect 18309 10368 18629 11392
rect 18309 10304 18317 10368
rect 18381 10304 18397 10368
rect 18461 10304 18477 10368
rect 18541 10304 18557 10368
rect 18621 10304 18629 10368
rect 18309 9280 18629 10304
rect 18309 9216 18317 9280
rect 18381 9216 18397 9280
rect 18461 9216 18477 9280
rect 18541 9216 18557 9280
rect 18621 9216 18629 9280
rect 18309 8192 18629 9216
rect 18309 8128 18317 8192
rect 18381 8128 18397 8192
rect 18461 8128 18477 8192
rect 18541 8128 18557 8192
rect 18621 8128 18629 8192
rect 18309 7104 18629 8128
rect 18309 7040 18317 7104
rect 18381 7040 18397 7104
rect 18461 7040 18477 7104
rect 18541 7040 18557 7104
rect 18621 7040 18629 7104
rect 18309 6016 18629 7040
rect 18309 5952 18317 6016
rect 18381 5952 18397 6016
rect 18461 5952 18477 6016
rect 18541 5952 18557 6016
rect 18621 5952 18629 6016
rect 18309 4928 18629 5952
rect 18309 4864 18317 4928
rect 18381 4864 18397 4928
rect 18461 4864 18477 4928
rect 18541 4864 18557 4928
rect 18621 4864 18629 4928
rect 18309 3840 18629 4864
rect 18309 3776 18317 3840
rect 18381 3776 18397 3840
rect 18461 3776 18477 3840
rect 18541 3776 18557 3840
rect 18621 3776 18629 3840
rect 18309 2752 18629 3776
rect 18309 2688 18317 2752
rect 18381 2688 18397 2752
rect 18461 2688 18477 2752
rect 18541 2688 18557 2752
rect 18621 2688 18629 2752
rect 18309 2128 18629 2688
rect 21782 23968 22102 24992
rect 21782 23904 21790 23968
rect 21854 23904 21870 23968
rect 21934 23904 21950 23968
rect 22014 23904 22030 23968
rect 22094 23904 22102 23968
rect 21782 22880 22102 23904
rect 21782 22816 21790 22880
rect 21854 22816 21870 22880
rect 21934 22816 21950 22880
rect 22014 22816 22030 22880
rect 22094 22816 22102 22880
rect 21782 21792 22102 22816
rect 21782 21728 21790 21792
rect 21854 21728 21870 21792
rect 21934 21728 21950 21792
rect 22014 21728 22030 21792
rect 22094 21728 22102 21792
rect 21782 20704 22102 21728
rect 21782 20640 21790 20704
rect 21854 20640 21870 20704
rect 21934 20640 21950 20704
rect 22014 20640 22030 20704
rect 22094 20640 22102 20704
rect 21782 19616 22102 20640
rect 21782 19552 21790 19616
rect 21854 19552 21870 19616
rect 21934 19552 21950 19616
rect 22014 19552 22030 19616
rect 22094 19552 22102 19616
rect 21782 18528 22102 19552
rect 21782 18464 21790 18528
rect 21854 18464 21870 18528
rect 21934 18464 21950 18528
rect 22014 18464 22030 18528
rect 22094 18464 22102 18528
rect 21782 17440 22102 18464
rect 21782 17376 21790 17440
rect 21854 17376 21870 17440
rect 21934 17376 21950 17440
rect 22014 17376 22030 17440
rect 22094 17376 22102 17440
rect 21782 16352 22102 17376
rect 21782 16288 21790 16352
rect 21854 16288 21870 16352
rect 21934 16288 21950 16352
rect 22014 16288 22030 16352
rect 22094 16288 22102 16352
rect 21782 15264 22102 16288
rect 21782 15200 21790 15264
rect 21854 15200 21870 15264
rect 21934 15200 21950 15264
rect 22014 15200 22030 15264
rect 22094 15200 22102 15264
rect 21782 14176 22102 15200
rect 21782 14112 21790 14176
rect 21854 14112 21870 14176
rect 21934 14112 21950 14176
rect 22014 14112 22030 14176
rect 22094 14112 22102 14176
rect 21782 13088 22102 14112
rect 21782 13024 21790 13088
rect 21854 13024 21870 13088
rect 21934 13024 21950 13088
rect 22014 13024 22030 13088
rect 22094 13024 22102 13088
rect 21782 12000 22102 13024
rect 21782 11936 21790 12000
rect 21854 11936 21870 12000
rect 21934 11936 21950 12000
rect 22014 11936 22030 12000
rect 22094 11936 22102 12000
rect 21782 10912 22102 11936
rect 21782 10848 21790 10912
rect 21854 10848 21870 10912
rect 21934 10848 21950 10912
rect 22014 10848 22030 10912
rect 22094 10848 22102 10912
rect 21782 9824 22102 10848
rect 21782 9760 21790 9824
rect 21854 9760 21870 9824
rect 21934 9760 21950 9824
rect 22014 9760 22030 9824
rect 22094 9760 22102 9824
rect 21782 8736 22102 9760
rect 21782 8672 21790 8736
rect 21854 8672 21870 8736
rect 21934 8672 21950 8736
rect 22014 8672 22030 8736
rect 22094 8672 22102 8736
rect 21782 7648 22102 8672
rect 21782 7584 21790 7648
rect 21854 7584 21870 7648
rect 21934 7584 21950 7648
rect 22014 7584 22030 7648
rect 22094 7584 22102 7648
rect 21782 6560 22102 7584
rect 21782 6496 21790 6560
rect 21854 6496 21870 6560
rect 21934 6496 21950 6560
rect 22014 6496 22030 6560
rect 22094 6496 22102 6560
rect 21782 5472 22102 6496
rect 21782 5408 21790 5472
rect 21854 5408 21870 5472
rect 21934 5408 21950 5472
rect 22014 5408 22030 5472
rect 22094 5408 22102 5472
rect 21782 4384 22102 5408
rect 21782 4320 21790 4384
rect 21854 4320 21870 4384
rect 21934 4320 21950 4384
rect 22014 4320 22030 4384
rect 22094 4320 22102 4384
rect 21782 3296 22102 4320
rect 21782 3232 21790 3296
rect 21854 3232 21870 3296
rect 21934 3232 21950 3296
rect 22014 3232 22030 3296
rect 22094 3232 22102 3296
rect 21782 2208 22102 3232
rect 21782 2144 21790 2208
rect 21854 2144 21870 2208
rect 21934 2144 21950 2208
rect 22014 2144 22030 2208
rect 22094 2144 22102 2208
rect 21782 2128 22102 2144
rect 25255 47360 25575 47376
rect 25255 47296 25263 47360
rect 25327 47296 25343 47360
rect 25407 47296 25423 47360
rect 25487 47296 25503 47360
rect 25567 47296 25575 47360
rect 25255 46272 25575 47296
rect 25255 46208 25263 46272
rect 25327 46208 25343 46272
rect 25407 46208 25423 46272
rect 25487 46208 25503 46272
rect 25567 46208 25575 46272
rect 25255 45184 25575 46208
rect 25255 45120 25263 45184
rect 25327 45120 25343 45184
rect 25407 45120 25423 45184
rect 25487 45120 25503 45184
rect 25567 45120 25575 45184
rect 25255 44096 25575 45120
rect 25255 44032 25263 44096
rect 25327 44032 25343 44096
rect 25407 44032 25423 44096
rect 25487 44032 25503 44096
rect 25567 44032 25575 44096
rect 25255 43008 25575 44032
rect 25255 42944 25263 43008
rect 25327 42944 25343 43008
rect 25407 42944 25423 43008
rect 25487 42944 25503 43008
rect 25567 42944 25575 43008
rect 25255 41920 25575 42944
rect 25255 41856 25263 41920
rect 25327 41856 25343 41920
rect 25407 41856 25423 41920
rect 25487 41856 25503 41920
rect 25567 41856 25575 41920
rect 25255 40832 25575 41856
rect 25255 40768 25263 40832
rect 25327 40768 25343 40832
rect 25407 40768 25423 40832
rect 25487 40768 25503 40832
rect 25567 40768 25575 40832
rect 25255 39744 25575 40768
rect 25255 39680 25263 39744
rect 25327 39680 25343 39744
rect 25407 39680 25423 39744
rect 25487 39680 25503 39744
rect 25567 39680 25575 39744
rect 25255 38656 25575 39680
rect 25255 38592 25263 38656
rect 25327 38592 25343 38656
rect 25407 38592 25423 38656
rect 25487 38592 25503 38656
rect 25567 38592 25575 38656
rect 25255 37568 25575 38592
rect 25255 37504 25263 37568
rect 25327 37504 25343 37568
rect 25407 37504 25423 37568
rect 25487 37504 25503 37568
rect 25567 37504 25575 37568
rect 25255 36480 25575 37504
rect 25255 36416 25263 36480
rect 25327 36416 25343 36480
rect 25407 36416 25423 36480
rect 25487 36416 25503 36480
rect 25567 36416 25575 36480
rect 25255 35392 25575 36416
rect 25255 35328 25263 35392
rect 25327 35328 25343 35392
rect 25407 35328 25423 35392
rect 25487 35328 25503 35392
rect 25567 35328 25575 35392
rect 25255 34304 25575 35328
rect 25255 34240 25263 34304
rect 25327 34240 25343 34304
rect 25407 34240 25423 34304
rect 25487 34240 25503 34304
rect 25567 34240 25575 34304
rect 25255 33216 25575 34240
rect 25255 33152 25263 33216
rect 25327 33152 25343 33216
rect 25407 33152 25423 33216
rect 25487 33152 25503 33216
rect 25567 33152 25575 33216
rect 25255 32128 25575 33152
rect 25255 32064 25263 32128
rect 25327 32064 25343 32128
rect 25407 32064 25423 32128
rect 25487 32064 25503 32128
rect 25567 32064 25575 32128
rect 25255 31040 25575 32064
rect 25255 30976 25263 31040
rect 25327 30976 25343 31040
rect 25407 30976 25423 31040
rect 25487 30976 25503 31040
rect 25567 30976 25575 31040
rect 25255 29952 25575 30976
rect 25255 29888 25263 29952
rect 25327 29888 25343 29952
rect 25407 29888 25423 29952
rect 25487 29888 25503 29952
rect 25567 29888 25575 29952
rect 25255 28864 25575 29888
rect 25255 28800 25263 28864
rect 25327 28800 25343 28864
rect 25407 28800 25423 28864
rect 25487 28800 25503 28864
rect 25567 28800 25575 28864
rect 25255 27776 25575 28800
rect 25255 27712 25263 27776
rect 25327 27712 25343 27776
rect 25407 27712 25423 27776
rect 25487 27712 25503 27776
rect 25567 27712 25575 27776
rect 25255 26688 25575 27712
rect 25255 26624 25263 26688
rect 25327 26624 25343 26688
rect 25407 26624 25423 26688
rect 25487 26624 25503 26688
rect 25567 26624 25575 26688
rect 25255 25600 25575 26624
rect 25255 25536 25263 25600
rect 25327 25536 25343 25600
rect 25407 25536 25423 25600
rect 25487 25536 25503 25600
rect 25567 25536 25575 25600
rect 25255 24512 25575 25536
rect 25255 24448 25263 24512
rect 25327 24448 25343 24512
rect 25407 24448 25423 24512
rect 25487 24448 25503 24512
rect 25567 24448 25575 24512
rect 25255 23424 25575 24448
rect 25255 23360 25263 23424
rect 25327 23360 25343 23424
rect 25407 23360 25423 23424
rect 25487 23360 25503 23424
rect 25567 23360 25575 23424
rect 25255 22336 25575 23360
rect 25255 22272 25263 22336
rect 25327 22272 25343 22336
rect 25407 22272 25423 22336
rect 25487 22272 25503 22336
rect 25567 22272 25575 22336
rect 25255 21248 25575 22272
rect 25255 21184 25263 21248
rect 25327 21184 25343 21248
rect 25407 21184 25423 21248
rect 25487 21184 25503 21248
rect 25567 21184 25575 21248
rect 25255 20160 25575 21184
rect 25255 20096 25263 20160
rect 25327 20096 25343 20160
rect 25407 20096 25423 20160
rect 25487 20096 25503 20160
rect 25567 20096 25575 20160
rect 25255 19072 25575 20096
rect 25255 19008 25263 19072
rect 25327 19008 25343 19072
rect 25407 19008 25423 19072
rect 25487 19008 25503 19072
rect 25567 19008 25575 19072
rect 25255 17984 25575 19008
rect 25255 17920 25263 17984
rect 25327 17920 25343 17984
rect 25407 17920 25423 17984
rect 25487 17920 25503 17984
rect 25567 17920 25575 17984
rect 25255 16896 25575 17920
rect 25255 16832 25263 16896
rect 25327 16832 25343 16896
rect 25407 16832 25423 16896
rect 25487 16832 25503 16896
rect 25567 16832 25575 16896
rect 25255 15808 25575 16832
rect 25255 15744 25263 15808
rect 25327 15744 25343 15808
rect 25407 15744 25423 15808
rect 25487 15744 25503 15808
rect 25567 15744 25575 15808
rect 25255 14720 25575 15744
rect 25255 14656 25263 14720
rect 25327 14656 25343 14720
rect 25407 14656 25423 14720
rect 25487 14656 25503 14720
rect 25567 14656 25575 14720
rect 25255 13632 25575 14656
rect 25255 13568 25263 13632
rect 25327 13568 25343 13632
rect 25407 13568 25423 13632
rect 25487 13568 25503 13632
rect 25567 13568 25575 13632
rect 25255 12544 25575 13568
rect 25255 12480 25263 12544
rect 25327 12480 25343 12544
rect 25407 12480 25423 12544
rect 25487 12480 25503 12544
rect 25567 12480 25575 12544
rect 25255 11456 25575 12480
rect 25255 11392 25263 11456
rect 25327 11392 25343 11456
rect 25407 11392 25423 11456
rect 25487 11392 25503 11456
rect 25567 11392 25575 11456
rect 25255 10368 25575 11392
rect 25255 10304 25263 10368
rect 25327 10304 25343 10368
rect 25407 10304 25423 10368
rect 25487 10304 25503 10368
rect 25567 10304 25575 10368
rect 25255 9280 25575 10304
rect 25255 9216 25263 9280
rect 25327 9216 25343 9280
rect 25407 9216 25423 9280
rect 25487 9216 25503 9280
rect 25567 9216 25575 9280
rect 25255 8192 25575 9216
rect 25255 8128 25263 8192
rect 25327 8128 25343 8192
rect 25407 8128 25423 8192
rect 25487 8128 25503 8192
rect 25567 8128 25575 8192
rect 25255 7104 25575 8128
rect 25255 7040 25263 7104
rect 25327 7040 25343 7104
rect 25407 7040 25423 7104
rect 25487 7040 25503 7104
rect 25567 7040 25575 7104
rect 25255 6016 25575 7040
rect 25255 5952 25263 6016
rect 25327 5952 25343 6016
rect 25407 5952 25423 6016
rect 25487 5952 25503 6016
rect 25567 5952 25575 6016
rect 25255 4928 25575 5952
rect 25255 4864 25263 4928
rect 25327 4864 25343 4928
rect 25407 4864 25423 4928
rect 25487 4864 25503 4928
rect 25567 4864 25575 4928
rect 25255 3840 25575 4864
rect 25255 3776 25263 3840
rect 25327 3776 25343 3840
rect 25407 3776 25423 3840
rect 25487 3776 25503 3840
rect 25567 3776 25575 3840
rect 25255 2752 25575 3776
rect 25255 2688 25263 2752
rect 25327 2688 25343 2752
rect 25407 2688 25423 2752
rect 25487 2688 25503 2752
rect 25567 2688 25575 2752
rect 25255 2128 25575 2688
rect 28728 46816 29048 47376
rect 28728 46752 28736 46816
rect 28800 46752 28816 46816
rect 28880 46752 28896 46816
rect 28960 46752 28976 46816
rect 29040 46752 29048 46816
rect 28728 45728 29048 46752
rect 28728 45664 28736 45728
rect 28800 45664 28816 45728
rect 28880 45664 28896 45728
rect 28960 45664 28976 45728
rect 29040 45664 29048 45728
rect 28728 44640 29048 45664
rect 28728 44576 28736 44640
rect 28800 44576 28816 44640
rect 28880 44576 28896 44640
rect 28960 44576 28976 44640
rect 29040 44576 29048 44640
rect 28728 43552 29048 44576
rect 28728 43488 28736 43552
rect 28800 43488 28816 43552
rect 28880 43488 28896 43552
rect 28960 43488 28976 43552
rect 29040 43488 29048 43552
rect 28728 42464 29048 43488
rect 28728 42400 28736 42464
rect 28800 42400 28816 42464
rect 28880 42400 28896 42464
rect 28960 42400 28976 42464
rect 29040 42400 29048 42464
rect 28728 41376 29048 42400
rect 28728 41312 28736 41376
rect 28800 41312 28816 41376
rect 28880 41312 28896 41376
rect 28960 41312 28976 41376
rect 29040 41312 29048 41376
rect 28728 40288 29048 41312
rect 28728 40224 28736 40288
rect 28800 40224 28816 40288
rect 28880 40224 28896 40288
rect 28960 40224 28976 40288
rect 29040 40224 29048 40288
rect 28728 39200 29048 40224
rect 28728 39136 28736 39200
rect 28800 39136 28816 39200
rect 28880 39136 28896 39200
rect 28960 39136 28976 39200
rect 29040 39136 29048 39200
rect 28728 38112 29048 39136
rect 28728 38048 28736 38112
rect 28800 38048 28816 38112
rect 28880 38048 28896 38112
rect 28960 38048 28976 38112
rect 29040 38048 29048 38112
rect 28728 37024 29048 38048
rect 28728 36960 28736 37024
rect 28800 36960 28816 37024
rect 28880 36960 28896 37024
rect 28960 36960 28976 37024
rect 29040 36960 29048 37024
rect 28728 35936 29048 36960
rect 28728 35872 28736 35936
rect 28800 35872 28816 35936
rect 28880 35872 28896 35936
rect 28960 35872 28976 35936
rect 29040 35872 29048 35936
rect 28728 34848 29048 35872
rect 28728 34784 28736 34848
rect 28800 34784 28816 34848
rect 28880 34784 28896 34848
rect 28960 34784 28976 34848
rect 29040 34784 29048 34848
rect 28728 33760 29048 34784
rect 28728 33696 28736 33760
rect 28800 33696 28816 33760
rect 28880 33696 28896 33760
rect 28960 33696 28976 33760
rect 29040 33696 29048 33760
rect 28728 32672 29048 33696
rect 28728 32608 28736 32672
rect 28800 32608 28816 32672
rect 28880 32608 28896 32672
rect 28960 32608 28976 32672
rect 29040 32608 29048 32672
rect 28728 31584 29048 32608
rect 28728 31520 28736 31584
rect 28800 31520 28816 31584
rect 28880 31520 28896 31584
rect 28960 31520 28976 31584
rect 29040 31520 29048 31584
rect 28728 30496 29048 31520
rect 28728 30432 28736 30496
rect 28800 30432 28816 30496
rect 28880 30432 28896 30496
rect 28960 30432 28976 30496
rect 29040 30432 29048 30496
rect 28728 29408 29048 30432
rect 28728 29344 28736 29408
rect 28800 29344 28816 29408
rect 28880 29344 28896 29408
rect 28960 29344 28976 29408
rect 29040 29344 29048 29408
rect 28728 28320 29048 29344
rect 28728 28256 28736 28320
rect 28800 28256 28816 28320
rect 28880 28256 28896 28320
rect 28960 28256 28976 28320
rect 29040 28256 29048 28320
rect 28728 27232 29048 28256
rect 28728 27168 28736 27232
rect 28800 27168 28816 27232
rect 28880 27168 28896 27232
rect 28960 27168 28976 27232
rect 29040 27168 29048 27232
rect 28728 26144 29048 27168
rect 28728 26080 28736 26144
rect 28800 26080 28816 26144
rect 28880 26080 28896 26144
rect 28960 26080 28976 26144
rect 29040 26080 29048 26144
rect 28728 25056 29048 26080
rect 28728 24992 28736 25056
rect 28800 24992 28816 25056
rect 28880 24992 28896 25056
rect 28960 24992 28976 25056
rect 29040 24992 29048 25056
rect 28728 23968 29048 24992
rect 28728 23904 28736 23968
rect 28800 23904 28816 23968
rect 28880 23904 28896 23968
rect 28960 23904 28976 23968
rect 29040 23904 29048 23968
rect 28728 22880 29048 23904
rect 28728 22816 28736 22880
rect 28800 22816 28816 22880
rect 28880 22816 28896 22880
rect 28960 22816 28976 22880
rect 29040 22816 29048 22880
rect 28728 21792 29048 22816
rect 28728 21728 28736 21792
rect 28800 21728 28816 21792
rect 28880 21728 28896 21792
rect 28960 21728 28976 21792
rect 29040 21728 29048 21792
rect 28728 20704 29048 21728
rect 28728 20640 28736 20704
rect 28800 20640 28816 20704
rect 28880 20640 28896 20704
rect 28960 20640 28976 20704
rect 29040 20640 29048 20704
rect 28728 19616 29048 20640
rect 28728 19552 28736 19616
rect 28800 19552 28816 19616
rect 28880 19552 28896 19616
rect 28960 19552 28976 19616
rect 29040 19552 29048 19616
rect 28728 18528 29048 19552
rect 28728 18464 28736 18528
rect 28800 18464 28816 18528
rect 28880 18464 28896 18528
rect 28960 18464 28976 18528
rect 29040 18464 29048 18528
rect 28728 17440 29048 18464
rect 28728 17376 28736 17440
rect 28800 17376 28816 17440
rect 28880 17376 28896 17440
rect 28960 17376 28976 17440
rect 29040 17376 29048 17440
rect 28728 16352 29048 17376
rect 28728 16288 28736 16352
rect 28800 16288 28816 16352
rect 28880 16288 28896 16352
rect 28960 16288 28976 16352
rect 29040 16288 29048 16352
rect 28728 15264 29048 16288
rect 28728 15200 28736 15264
rect 28800 15200 28816 15264
rect 28880 15200 28896 15264
rect 28960 15200 28976 15264
rect 29040 15200 29048 15264
rect 28728 14176 29048 15200
rect 28728 14112 28736 14176
rect 28800 14112 28816 14176
rect 28880 14112 28896 14176
rect 28960 14112 28976 14176
rect 29040 14112 29048 14176
rect 28728 13088 29048 14112
rect 28728 13024 28736 13088
rect 28800 13024 28816 13088
rect 28880 13024 28896 13088
rect 28960 13024 28976 13088
rect 29040 13024 29048 13088
rect 28728 12000 29048 13024
rect 28728 11936 28736 12000
rect 28800 11936 28816 12000
rect 28880 11936 28896 12000
rect 28960 11936 28976 12000
rect 29040 11936 29048 12000
rect 28728 10912 29048 11936
rect 28728 10848 28736 10912
rect 28800 10848 28816 10912
rect 28880 10848 28896 10912
rect 28960 10848 28976 10912
rect 29040 10848 29048 10912
rect 28728 9824 29048 10848
rect 28728 9760 28736 9824
rect 28800 9760 28816 9824
rect 28880 9760 28896 9824
rect 28960 9760 28976 9824
rect 29040 9760 29048 9824
rect 28728 8736 29048 9760
rect 28728 8672 28736 8736
rect 28800 8672 28816 8736
rect 28880 8672 28896 8736
rect 28960 8672 28976 8736
rect 29040 8672 29048 8736
rect 28728 7648 29048 8672
rect 28728 7584 28736 7648
rect 28800 7584 28816 7648
rect 28880 7584 28896 7648
rect 28960 7584 28976 7648
rect 29040 7584 29048 7648
rect 28728 6560 29048 7584
rect 28728 6496 28736 6560
rect 28800 6496 28816 6560
rect 28880 6496 28896 6560
rect 28960 6496 28976 6560
rect 29040 6496 29048 6560
rect 28728 5472 29048 6496
rect 28728 5408 28736 5472
rect 28800 5408 28816 5472
rect 28880 5408 28896 5472
rect 28960 5408 28976 5472
rect 29040 5408 29048 5472
rect 28728 4384 29048 5408
rect 28728 4320 28736 4384
rect 28800 4320 28816 4384
rect 28880 4320 28896 4384
rect 28960 4320 28976 4384
rect 29040 4320 29048 4384
rect 28728 3296 29048 4320
rect 28728 3232 28736 3296
rect 28800 3232 28816 3296
rect 28880 3232 28896 3296
rect 28960 3232 28976 3296
rect 29040 3232 29048 3296
rect 28728 2208 29048 3232
rect 28728 2144 28736 2208
rect 28800 2144 28816 2208
rect 28880 2144 28896 2208
rect 28960 2144 28976 2208
rect 29040 2144 29048 2208
rect 28728 2128 29048 2144
use sky130_fd_sc_hd__decap_4  FILLER_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 1380 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 1748 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11
timestamp 1667941163
transform 1 0 2116 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15
timestamp 1667941163
transform 1 0 2484 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19
timestamp 1667941163
transform 1 0 2852 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 3496 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29
timestamp 1667941163
transform 1 0 3772 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52
timestamp 1667941163
transform 1 0 5888 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69
timestamp 1667941163
transform 1 0 7452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_81 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_85
timestamp 1667941163
transform 1 0 8924 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97
timestamp 1667941163
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_109
timestamp 1667941163
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113
timestamp 1667941163
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_125
timestamp 1667941163
transform 1 0 12604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_137
timestamp 1667941163
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_141
timestamp 1667941163
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_153
timestamp 1667941163
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_165
timestamp 1667941163
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_169
timestamp 1667941163
transform 1 0 16652 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_175
timestamp 1667941163
transform 1 0 17204 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_182
timestamp 1667941163
transform 1 0 17848 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_194
timestamp 1667941163
transform 1 0 18952 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_197
timestamp 1667941163
transform 1 0 19228 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_220
timestamp 1667941163
transform 1 0 21344 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_225
timestamp 1667941163
transform 1 0 21804 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_237
timestamp 1667941163
transform 1 0 22908 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_249
timestamp 1667941163
transform 1 0 24012 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_253
timestamp 1667941163
transform 1 0 24380 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_265 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 25484 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_273
timestamp 1667941163
transform 1 0 26220 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_278
timestamp 1667941163
transform 1 0 26680 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_281
timestamp 1667941163
transform 1 0 26956 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_292 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 27968 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_298
timestamp 1667941163
transform 1 0 28520 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_3
timestamp 1667941163
transform 1 0 1380 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_28
timestamp 1667941163
transform 1 0 3680 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_32
timestamp 1667941163
transform 1 0 4048 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_54
timestamp 1667941163
transform 1 0 6072 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_1_57
timestamp 1667941163
transform 1 0 6348 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_84
timestamp 1667941163
transform 1 0 8832 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_1_109
timestamp 1667941163
transform 1 0 11132 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_1_113
timestamp 1667941163
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_125
timestamp 1667941163
transform 1 0 12604 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_130
timestamp 1667941163
transform 1 0 13064 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_138
timestamp 1667941163
transform 1 0 13800 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_1_161
timestamp 1667941163
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 1667941163
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_169
timestamp 1667941163
transform 1 0 16652 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_192
timestamp 1667941163
transform 1 0 18768 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_217
timestamp 1667941163
transform 1 0 21068 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_223
timestamp 1667941163
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_225
timestamp 1667941163
transform 1 0 21804 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_237
timestamp 1667941163
transform 1 0 22908 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_249
timestamp 1667941163
transform 1 0 24012 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_278
timestamp 1667941163
transform 1 0 26680 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_281
timestamp 1667941163
transform 1 0 26956 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_286
timestamp 1667941163
transform 1 0 27416 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_290
timestamp 1667941163
transform 1 0 27784 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_294
timestamp 1667941163
transform 1 0 28152 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_298
timestamp 1667941163
transform 1 0 28520 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_3
timestamp 1667941163
transform 1 0 1380 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_26
timestamp 1667941163
transform 1 0 3496 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_29
timestamp 1667941163
transform 1 0 3772 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_36
timestamp 1667941163
transform 1 0 4416 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_42
timestamp 1667941163
transform 1 0 4968 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_46
timestamp 1667941163
transform 1 0 5336 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_71
timestamp 1667941163
transform 1 0 7636 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_78
timestamp 1667941163
transform 1 0 8280 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_2_85
timestamp 1667941163
transform 1 0 8924 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_90
timestamp 1667941163
transform 1 0 9384 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_97
timestamp 1667941163
transform 1 0 10028 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_122
timestamp 1667941163
transform 1 0 12328 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_131
timestamp 1667941163
transform 1 0 13156 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_138
timestamp 1667941163
transform 1 0 13800 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_141
timestamp 1667941163
transform 1 0 14076 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_146
timestamp 1667941163
transform 1 0 14536 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_158
timestamp 1667941163
transform 1 0 15640 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_165
timestamp 1667941163
transform 1 0 16284 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_172
timestamp 1667941163
transform 1 0 16928 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_181
timestamp 1667941163
transform 1 0 17756 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_188
timestamp 1667941163
transform 1 0 18400 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_197
timestamp 1667941163
transform 1 0 19228 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_2_202
timestamp 1667941163
transform 1 0 19688 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_208
timestamp 1667941163
transform 1 0 20240 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_230
timestamp 1667941163
transform 1 0 22264 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_242
timestamp 1667941163
transform 1 0 23368 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_250
timestamp 1667941163
transform 1 0 24104 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_253
timestamp 1667941163
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_265
timestamp 1667941163
transform 1 0 25484 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_272
timestamp 1667941163
transform 1 0 26128 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_297
timestamp 1667941163
transform 1 0 28428 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_3
timestamp 1667941163
transform 1 0 1380 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_10
timestamp 1667941163
transform 1 0 2024 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_17
timestamp 1667941163
transform 1 0 2668 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_24
timestamp 1667941163
transform 1 0 3312 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_49
timestamp 1667941163
transform 1 0 5612 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1667941163
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_57
timestamp 1667941163
transform 1 0 6348 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_62
timestamp 1667941163
transform 1 0 6808 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_70
timestamp 1667941163
transform 1 0 7544 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_75
timestamp 1667941163
transform 1 0 8004 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_87
timestamp 1667941163
transform 1 0 9108 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_3_99
timestamp 1667941163
transform 1 0 10212 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp 1667941163
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1667941163
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_113
timestamp 1667941163
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_125
timestamp 1667941163
transform 1 0 12604 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_148
timestamp 1667941163
transform 1 0 14720 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_160
timestamp 1667941163
transform 1 0 15824 0 -1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_3_169
timestamp 1667941163
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_181
timestamp 1667941163
transform 1 0 17756 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_189
timestamp 1667941163
transform 1 0 18492 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_194
timestamp 1667941163
transform 1 0 18952 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_206
timestamp 1667941163
transform 1 0 20056 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_213
timestamp 1667941163
transform 1 0 20700 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_220
timestamp 1667941163
transform 1 0 21344 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_225
timestamp 1667941163
transform 1 0 21804 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_3_232
timestamp 1667941163
transform 1 0 22448 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_244
timestamp 1667941163
transform 1 0 23552 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_256
timestamp 1667941163
transform 1 0 24656 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_268
timestamp 1667941163
transform 1 0 25760 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_281
timestamp 1667941163
transform 1 0 26956 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_3_292
timestamp 1667941163
transform 1 0 27968 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_298
timestamp 1667941163
transform 1 0 28520 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_3
timestamp 1667941163
transform 1 0 1380 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_8
timestamp 1667941163
transform 1 0 1840 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_15
timestamp 1667941163
transform 1 0 2484 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_19
timestamp 1667941163
transform 1 0 2852 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_23
timestamp 1667941163
transform 1 0 3220 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1667941163
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_29
timestamp 1667941163
transform 1 0 3772 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_34
timestamp 1667941163
transform 1 0 4232 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_41
timestamp 1667941163
transform 1 0 4876 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_66
timestamp 1667941163
transform 1 0 7176 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_78
timestamp 1667941163
transform 1 0 8280 0 1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1667941163
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_97
timestamp 1667941163
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_109
timestamp 1667941163
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_121
timestamp 1667941163
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp 1667941163
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1667941163
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_141
timestamp 1667941163
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_153
timestamp 1667941163
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_165
timestamp 1667941163
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_177
timestamp 1667941163
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_189
timestamp 1667941163
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 1667941163
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_197
timestamp 1667941163
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_209
timestamp 1667941163
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_221
timestamp 1667941163
transform 1 0 21436 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_227
timestamp 1667941163
transform 1 0 21988 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_249
timestamp 1667941163
transform 1 0 24012 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_253
timestamp 1667941163
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_265
timestamp 1667941163
transform 1 0 25484 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_273
timestamp 1667941163
transform 1 0 26220 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_297
timestamp 1667941163
transform 1 0 28428 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_3
timestamp 1667941163
transform 1 0 1380 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_9
timestamp 1667941163
transform 1 0 1932 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_16
timestamp 1667941163
transform 1 0 2576 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_41
timestamp 1667941163
transform 1 0 4876 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_45
timestamp 1667941163
transform 1 0 5244 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_49
timestamp 1667941163
transform 1 0 5612 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1667941163
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1667941163
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1667941163
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_81
timestamp 1667941163
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_93
timestamp 1667941163
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 1667941163
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1667941163
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_113
timestamp 1667941163
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_125
timestamp 1667941163
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_137
timestamp 1667941163
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_149
timestamp 1667941163
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp 1667941163
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1667941163
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_169
timestamp 1667941163
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_181
timestamp 1667941163
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_193
timestamp 1667941163
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_205
timestamp 1667941163
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_217
timestamp 1667941163
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_223
timestamp 1667941163
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_225
timestamp 1667941163
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_237
timestamp 1667941163
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_249
timestamp 1667941163
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_261
timestamp 1667941163
transform 1 0 25116 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_5_273
timestamp 1667941163
transform 1 0 26220 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_5_277
timestamp 1667941163
transform 1 0 26588 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_281
timestamp 1667941163
transform 1 0 26956 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_286
timestamp 1667941163
transform 1 0 27416 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_290
timestamp 1667941163
transform 1 0 27784 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_294
timestamp 1667941163
transform 1 0 28152 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_298
timestamp 1667941163
transform 1 0 28520 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_3
timestamp 1667941163
transform 1 0 1380 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_26
timestamp 1667941163
transform 1 0 3496 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_29
timestamp 1667941163
transform 1 0 3772 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_37
timestamp 1667941163
transform 1 0 4508 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_42
timestamp 1667941163
transform 1 0 4968 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_54
timestamp 1667941163
transform 1 0 6072 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_66
timestamp 1667941163
transform 1 0 7176 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_78
timestamp 1667941163
transform 1 0 8280 0 1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1667941163
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_97
timestamp 1667941163
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_109
timestamp 1667941163
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_121
timestamp 1667941163
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1667941163
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1667941163
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_141
timestamp 1667941163
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_153
timestamp 1667941163
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_165
timestamp 1667941163
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_177
timestamp 1667941163
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_189
timestamp 1667941163
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1667941163
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_197
timestamp 1667941163
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_209
timestamp 1667941163
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_221
timestamp 1667941163
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_233
timestamp 1667941163
transform 1 0 22540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_245
timestamp 1667941163
transform 1 0 23644 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp 1667941163
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_253
timestamp 1667941163
transform 1 0 24380 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_261
timestamp 1667941163
transform 1 0 25116 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_271
timestamp 1667941163
transform 1 0 26036 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_6_296
timestamp 1667941163
transform 1 0 28336 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_3
timestamp 1667941163
transform 1 0 1380 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_9
timestamp 1667941163
transform 1 0 1932 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_16
timestamp 1667941163
transform 1 0 2576 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_41
timestamp 1667941163
transform 1 0 4876 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_7_53
timestamp 1667941163
transform 1 0 5980 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1667941163
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_69
timestamp 1667941163
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_81
timestamp 1667941163
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_93
timestamp 1667941163
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 1667941163
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1667941163
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_113
timestamp 1667941163
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_125
timestamp 1667941163
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_137
timestamp 1667941163
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_149
timestamp 1667941163
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_161
timestamp 1667941163
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1667941163
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_169
timestamp 1667941163
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_181
timestamp 1667941163
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_193
timestamp 1667941163
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_205
timestamp 1667941163
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_217
timestamp 1667941163
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp 1667941163
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_225
timestamp 1667941163
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_237
timestamp 1667941163
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_249
timestamp 1667941163
transform 1 0 24012 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_278
timestamp 1667941163
transform 1 0 26680 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_281
timestamp 1667941163
transform 1 0 26956 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_285
timestamp 1667941163
transform 1 0 27324 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_289
timestamp 1667941163
transform 1 0 27692 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_297
timestamp 1667941163
transform 1 0 28428 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_3
timestamp 1667941163
transform 1 0 1380 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_26
timestamp 1667941163
transform 1 0 3496 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1667941163
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_41
timestamp 1667941163
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_53
timestamp 1667941163
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_65
timestamp 1667941163
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1667941163
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1667941163
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_85
timestamp 1667941163
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_97
timestamp 1667941163
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_109
timestamp 1667941163
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_121
timestamp 1667941163
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_133
timestamp 1667941163
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1667941163
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_141
timestamp 1667941163
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_153
timestamp 1667941163
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_165
timestamp 1667941163
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_177
timestamp 1667941163
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_189
timestamp 1667941163
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1667941163
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_197
timestamp 1667941163
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_209
timestamp 1667941163
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_221
timestamp 1667941163
transform 1 0 21436 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_233
timestamp 1667941163
transform 1 0 22540 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_8_245
timestamp 1667941163
transform 1 0 23644 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_250
timestamp 1667941163
transform 1 0 24104 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_253
timestamp 1667941163
transform 1 0 24380 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_276
timestamp 1667941163
transform 1 0 26496 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_291
timestamp 1667941163
transform 1 0 27876 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_9_3
timestamp 1667941163
transform 1 0 1380 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_9
timestamp 1667941163
transform 1 0 1932 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_13
timestamp 1667941163
transform 1 0 2300 0 -1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_9_24
timestamp 1667941163
transform 1 0 3312 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_36
timestamp 1667941163
transform 1 0 4416 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_48
timestamp 1667941163
transform 1 0 5520 0 -1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 1667941163
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_69
timestamp 1667941163
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_81
timestamp 1667941163
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_93
timestamp 1667941163
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_105
timestamp 1667941163
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1667941163
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_113
timestamp 1667941163
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_125
timestamp 1667941163
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_137
timestamp 1667941163
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_149
timestamp 1667941163
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_161
timestamp 1667941163
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1667941163
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_169
timestamp 1667941163
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_181
timestamp 1667941163
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_193
timestamp 1667941163
transform 1 0 18860 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_205
timestamp 1667941163
transform 1 0 19964 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_217
timestamp 1667941163
transform 1 0 21068 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_223
timestamp 1667941163
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_225
timestamp 1667941163
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_237
timestamp 1667941163
transform 1 0 22908 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_249
timestamp 1667941163
transform 1 0 24012 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_278
timestamp 1667941163
transform 1 0 26680 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_9_281
timestamp 1667941163
transform 1 0 26956 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_287
timestamp 1667941163
transform 1 0 27508 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_291
timestamp 1667941163
transform 1 0 27876 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_10_3
timestamp 1667941163
transform 1 0 1380 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_9
timestamp 1667941163
transform 1 0 1932 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_13
timestamp 1667941163
transform 1 0 2300 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_10_25
timestamp 1667941163
transform 1 0 3404 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_29
timestamp 1667941163
transform 1 0 3772 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_52
timestamp 1667941163
transform 1 0 5888 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_64
timestamp 1667941163
transform 1 0 6992 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_76
timestamp 1667941163
transform 1 0 8096 0 1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_10_85
timestamp 1667941163
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_97
timestamp 1667941163
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_109
timestamp 1667941163
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_121
timestamp 1667941163
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_133
timestamp 1667941163
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1667941163
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_141
timestamp 1667941163
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_153
timestamp 1667941163
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_165
timestamp 1667941163
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_177
timestamp 1667941163
transform 1 0 17388 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_189
timestamp 1667941163
transform 1 0 18492 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_195
timestamp 1667941163
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_197
timestamp 1667941163
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_209
timestamp 1667941163
transform 1 0 20332 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_221
timestamp 1667941163
transform 1 0 21436 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_233
timestamp 1667941163
transform 1 0 22540 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_245
timestamp 1667941163
transform 1 0 23644 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_251
timestamp 1667941163
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_253
timestamp 1667941163
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_265
timestamp 1667941163
transform 1 0 25484 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_273
timestamp 1667941163
transform 1 0 26220 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_297
timestamp 1667941163
transform 1 0 28428 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_3
timestamp 1667941163
transform 1 0 1380 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_27
timestamp 1667941163
transform 1 0 3588 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_34
timestamp 1667941163
transform 1 0 4232 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_11_41
timestamp 1667941163
transform 1 0 4876 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_11_53
timestamp 1667941163
transform 1 0 5980 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_11_57
timestamp 1667941163
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_69
timestamp 1667941163
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_81
timestamp 1667941163
transform 1 0 8556 0 -1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_11_92
timestamp 1667941163
transform 1 0 9568 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_104
timestamp 1667941163
transform 1 0 10672 0 -1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_11_113
timestamp 1667941163
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_125
timestamp 1667941163
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_137
timestamp 1667941163
transform 1 0 13708 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_149
timestamp 1667941163
transform 1 0 14812 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_161
timestamp 1667941163
transform 1 0 15916 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp 1667941163
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_169
timestamp 1667941163
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_181
timestamp 1667941163
transform 1 0 17756 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_193
timestamp 1667941163
transform 1 0 18860 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_205
timestamp 1667941163
transform 1 0 19964 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_217
timestamp 1667941163
transform 1 0 21068 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_223
timestamp 1667941163
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_225
timestamp 1667941163
transform 1 0 21804 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_237
timestamp 1667941163
transform 1 0 22908 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_249
timestamp 1667941163
transform 1 0 24012 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_261
timestamp 1667941163
transform 1 0 25116 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_273
timestamp 1667941163
transform 1 0 26220 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_278
timestamp 1667941163
transform 1 0 26680 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_281
timestamp 1667941163
transform 1 0 26956 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_11_292
timestamp 1667941163
transform 1 0 27968 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_298
timestamp 1667941163
transform 1 0 28520 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_3
timestamp 1667941163
transform 1 0 1380 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_26
timestamp 1667941163
transform 1 0 3496 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_29
timestamp 1667941163
transform 1 0 3772 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_34
timestamp 1667941163
transform 1 0 4232 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_46
timestamp 1667941163
transform 1 0 5336 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_58
timestamp 1667941163
transform 1 0 6440 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_70
timestamp 1667941163
transform 1 0 7544 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_82
timestamp 1667941163
transform 1 0 8648 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_85
timestamp 1667941163
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_97
timestamp 1667941163
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_109
timestamp 1667941163
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_121
timestamp 1667941163
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_133
timestamp 1667941163
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1667941163
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_141
timestamp 1667941163
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_153
timestamp 1667941163
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_165
timestamp 1667941163
transform 1 0 16284 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_177
timestamp 1667941163
transform 1 0 17388 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_189
timestamp 1667941163
transform 1 0 18492 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_195
timestamp 1667941163
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_197
timestamp 1667941163
transform 1 0 19228 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_209
timestamp 1667941163
transform 1 0 20332 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_221
timestamp 1667941163
transform 1 0 21436 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_233
timestamp 1667941163
transform 1 0 22540 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_245
timestamp 1667941163
transform 1 0 23644 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_251
timestamp 1667941163
transform 1 0 24196 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_253
timestamp 1667941163
transform 1 0 24380 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_265
timestamp 1667941163
transform 1 0 25484 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_287
timestamp 1667941163
transform 1 0 27508 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_294
timestamp 1667941163
transform 1 0 28152 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_298
timestamp 1667941163
transform 1 0 28520 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_13_3
timestamp 1667941163
transform 1 0 1380 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_9
timestamp 1667941163
transform 1 0 1932 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_16
timestamp 1667941163
transform 1 0 2576 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_20
timestamp 1667941163
transform 1 0 2944 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_42
timestamp 1667941163
transform 1 0 4968 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_54
timestamp 1667941163
transform 1 0 6072 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_57
timestamp 1667941163
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_69
timestamp 1667941163
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_81
timestamp 1667941163
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_93
timestamp 1667941163
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_105
timestamp 1667941163
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1667941163
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_113
timestamp 1667941163
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_125
timestamp 1667941163
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_137
timestamp 1667941163
transform 1 0 13708 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_149
timestamp 1667941163
transform 1 0 14812 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_161
timestamp 1667941163
transform 1 0 15916 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 1667941163
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_169
timestamp 1667941163
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_181
timestamp 1667941163
transform 1 0 17756 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_193
timestamp 1667941163
transform 1 0 18860 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_205
timestamp 1667941163
transform 1 0 19964 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_217
timestamp 1667941163
transform 1 0 21068 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_223
timestamp 1667941163
transform 1 0 21620 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_225
timestamp 1667941163
transform 1 0 21804 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_237
timestamp 1667941163
transform 1 0 22908 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_249
timestamp 1667941163
transform 1 0 24012 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_261
timestamp 1667941163
transform 1 0 25116 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_267
timestamp 1667941163
transform 1 0 25668 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_271
timestamp 1667941163
transform 1 0 26036 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_279
timestamp 1667941163
transform 1 0 26772 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_281
timestamp 1667941163
transform 1 0 26956 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_287
timestamp 1667941163
transform 1 0 27508 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_291
timestamp 1667941163
transform 1 0 27876 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_14_3
timestamp 1667941163
transform 1 0 1380 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_10
timestamp 1667941163
transform 1 0 2024 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_18
timestamp 1667941163
transform 1 0 2760 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_24
timestamp 1667941163
transform 1 0 3312 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_14_29
timestamp 1667941163
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_41
timestamp 1667941163
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_53
timestamp 1667941163
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_65
timestamp 1667941163
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp 1667941163
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1667941163
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_85
timestamp 1667941163
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_97
timestamp 1667941163
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_109
timestamp 1667941163
transform 1 0 11132 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_121
timestamp 1667941163
transform 1 0 12236 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_133
timestamp 1667941163
transform 1 0 13340 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1667941163
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_141
timestamp 1667941163
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_153
timestamp 1667941163
transform 1 0 15180 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_165
timestamp 1667941163
transform 1 0 16284 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_177
timestamp 1667941163
transform 1 0 17388 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_189
timestamp 1667941163
transform 1 0 18492 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_195
timestamp 1667941163
transform 1 0 19044 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_197
timestamp 1667941163
transform 1 0 19228 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_209
timestamp 1667941163
transform 1 0 20332 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_221
timestamp 1667941163
transform 1 0 21436 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_233
timestamp 1667941163
transform 1 0 22540 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_245
timestamp 1667941163
transform 1 0 23644 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_251
timestamp 1667941163
transform 1 0 24196 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_253
timestamp 1667941163
transform 1 0 24380 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_265
timestamp 1667941163
transform 1 0 25484 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_273
timestamp 1667941163
transform 1 0 26220 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_297
timestamp 1667941163
transform 1 0 28428 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3
timestamp 1667941163
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_15
timestamp 1667941163
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_27
timestamp 1667941163
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_39
timestamp 1667941163
transform 1 0 4692 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_51
timestamp 1667941163
transform 1 0 5796 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1667941163
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_57
timestamp 1667941163
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_69
timestamp 1667941163
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_81
timestamp 1667941163
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_93
timestamp 1667941163
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_105
timestamp 1667941163
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1667941163
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_113
timestamp 1667941163
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_125
timestamp 1667941163
transform 1 0 12604 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_137
timestamp 1667941163
transform 1 0 13708 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_149
timestamp 1667941163
transform 1 0 14812 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_161
timestamp 1667941163
transform 1 0 15916 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_167
timestamp 1667941163
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_169
timestamp 1667941163
transform 1 0 16652 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_181
timestamp 1667941163
transform 1 0 17756 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_193
timestamp 1667941163
transform 1 0 18860 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_205
timestamp 1667941163
transform 1 0 19964 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_15_218
timestamp 1667941163
transform 1 0 21160 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_15_225
timestamp 1667941163
transform 1 0 21804 0 -1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_15_236
timestamp 1667941163
transform 1 0 22816 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_248
timestamp 1667941163
transform 1 0 23920 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_260
timestamp 1667941163
transform 1 0 25024 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_15_272
timestamp 1667941163
transform 1 0 26128 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_278
timestamp 1667941163
transform 1 0 26680 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_281
timestamp 1667941163
transform 1 0 26956 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_286
timestamp 1667941163
transform 1 0 27416 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_290
timestamp 1667941163
transform 1 0 27784 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_294
timestamp 1667941163
transform 1 0 28152 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_298
timestamp 1667941163
transform 1 0 28520 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_16_3
timestamp 1667941163
transform 1 0 1380 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_9
timestamp 1667941163
transform 1 0 1932 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_16
timestamp 1667941163
transform 1 0 2576 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_29
timestamp 1667941163
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_41
timestamp 1667941163
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_53
timestamp 1667941163
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_65
timestamp 1667941163
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp 1667941163
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1667941163
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_85
timestamp 1667941163
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_97
timestamp 1667941163
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_109
timestamp 1667941163
transform 1 0 11132 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_121
timestamp 1667941163
transform 1 0 12236 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_133
timestamp 1667941163
transform 1 0 13340 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 1667941163
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_141
timestamp 1667941163
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_153
timestamp 1667941163
transform 1 0 15180 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_165
timestamp 1667941163
transform 1 0 16284 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_177
timestamp 1667941163
transform 1 0 17388 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_189
timestamp 1667941163
transform 1 0 18492 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_195
timestamp 1667941163
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_16_197
timestamp 1667941163
transform 1 0 19228 0 1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_16_205
timestamp 1667941163
transform 1 0 19964 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_226
timestamp 1667941163
transform 1 0 21896 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_233
timestamp 1667941163
transform 1 0 22540 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_245
timestamp 1667941163
transform 1 0 23644 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_251
timestamp 1667941163
transform 1 0 24196 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_253
timestamp 1667941163
transform 1 0 24380 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_262
timestamp 1667941163
transform 1 0 25208 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_274
timestamp 1667941163
transform 1 0 26312 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_297
timestamp 1667941163
transform 1 0 28428 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_3
timestamp 1667941163
transform 1 0 1380 0 -1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_17_27
timestamp 1667941163
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_39
timestamp 1667941163
transform 1 0 4692 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_51
timestamp 1667941163
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1667941163
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_57
timestamp 1667941163
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_69
timestamp 1667941163
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_81
timestamp 1667941163
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_93
timestamp 1667941163
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_105
timestamp 1667941163
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1667941163
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_113
timestamp 1667941163
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_125
timestamp 1667941163
transform 1 0 12604 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_137
timestamp 1667941163
transform 1 0 13708 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_149
timestamp 1667941163
transform 1 0 14812 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_161
timestamp 1667941163
transform 1 0 15916 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_167
timestamp 1667941163
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_169
timestamp 1667941163
transform 1 0 16652 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_181
timestamp 1667941163
transform 1 0 17756 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_193
timestamp 1667941163
transform 1 0 18860 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_17_204
timestamp 1667941163
transform 1 0 19872 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_17_219
timestamp 1667941163
transform 1 0 21252 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_223
timestamp 1667941163
transform 1 0 21620 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_225
timestamp 1667941163
transform 1 0 21804 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_235
timestamp 1667941163
transform 1 0 22724 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_247
timestamp 1667941163
transform 1 0 23828 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_258
timestamp 1667941163
transform 1 0 24840 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_265
timestamp 1667941163
transform 1 0 25484 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_17_277
timestamp 1667941163
transform 1 0 26588 0 -1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_17_281
timestamp 1667941163
transform 1 0 26956 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_293
timestamp 1667941163
transform 1 0 28060 0 -1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3
timestamp 1667941163
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_15
timestamp 1667941163
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1667941163
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_29
timestamp 1667941163
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_41
timestamp 1667941163
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_53
timestamp 1667941163
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_65
timestamp 1667941163
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_77
timestamp 1667941163
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1667941163
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_85
timestamp 1667941163
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_97
timestamp 1667941163
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_109
timestamp 1667941163
transform 1 0 11132 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_121
timestamp 1667941163
transform 1 0 12236 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_133
timestamp 1667941163
transform 1 0 13340 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_139
timestamp 1667941163
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_141
timestamp 1667941163
transform 1 0 14076 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_153
timestamp 1667941163
transform 1 0 15180 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_165
timestamp 1667941163
transform 1 0 16284 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_177
timestamp 1667941163
transform 1 0 17388 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_189
timestamp 1667941163
transform 1 0 18492 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_195
timestamp 1667941163
transform 1 0 19044 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_197
timestamp 1667941163
transform 1 0 19228 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_18_202
timestamp 1667941163
transform 1 0 19688 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_208
timestamp 1667941163
transform 1 0 20240 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_218
timestamp 1667941163
transform 1 0 21160 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_225
timestamp 1667941163
transform 1 0 21804 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_237
timestamp 1667941163
transform 1 0 22908 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_248
timestamp 1667941163
transform 1 0 23920 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_253
timestamp 1667941163
transform 1 0 24380 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_263
timestamp 1667941163
transform 1 0 25300 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_271
timestamp 1667941163
transform 1 0 26036 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_275
timestamp 1667941163
transform 1 0 26404 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_297
timestamp 1667941163
transform 1 0 28428 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_19_3
timestamp 1667941163
transform 1 0 1380 0 -1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_19_12
timestamp 1667941163
transform 1 0 2208 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_24
timestamp 1667941163
transform 1 0 3312 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_36
timestamp 1667941163
transform 1 0 4416 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_48
timestamp 1667941163
transform 1 0 5520 0 -1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_19_57
timestamp 1667941163
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_69
timestamp 1667941163
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_81
timestamp 1667941163
transform 1 0 8556 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_93
timestamp 1667941163
transform 1 0 9660 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_105
timestamp 1667941163
transform 1 0 10764 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1667941163
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_113
timestamp 1667941163
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_125
timestamp 1667941163
transform 1 0 12604 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_137
timestamp 1667941163
transform 1 0 13708 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_149
timestamp 1667941163
transform 1 0 14812 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_161
timestamp 1667941163
transform 1 0 15916 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_167
timestamp 1667941163
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_169
timestamp 1667941163
transform 1 0 16652 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_181
timestamp 1667941163
transform 1 0 17756 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_193
timestamp 1667941163
transform 1 0 18860 0 -1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_19_202
timestamp 1667941163
transform 1 0 19688 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_214
timestamp 1667941163
transform 1 0 20792 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_222
timestamp 1667941163
transform 1 0 21528 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_225
timestamp 1667941163
transform 1 0 21804 0 -1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_19_236
timestamp 1667941163
transform 1 0 22816 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_248
timestamp 1667941163
transform 1 0 23920 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_258
timestamp 1667941163
transform 1 0 24840 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_270
timestamp 1667941163
transform 1 0 25944 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_278
timestamp 1667941163
transform 1 0 26680 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_281
timestamp 1667941163
transform 1 0 26956 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_287
timestamp 1667941163
transform 1 0 27508 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_294
timestamp 1667941163
transform 1 0 28152 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_298
timestamp 1667941163
transform 1 0 28520 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_3
timestamp 1667941163
transform 1 0 1380 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_26
timestamp 1667941163
transform 1 0 3496 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_29
timestamp 1667941163
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_41
timestamp 1667941163
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_53
timestamp 1667941163
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_65
timestamp 1667941163
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_77
timestamp 1667941163
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1667941163
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_85
timestamp 1667941163
transform 1 0 8924 0 1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_20_96
timestamp 1667941163
transform 1 0 9936 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_108
timestamp 1667941163
transform 1 0 11040 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_120
timestamp 1667941163
transform 1 0 12144 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_132
timestamp 1667941163
transform 1 0 13248 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_141
timestamp 1667941163
transform 1 0 14076 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_146
timestamp 1667941163
transform 1 0 14536 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_153
timestamp 1667941163
transform 1 0 15180 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_20_165
timestamp 1667941163
transform 1 0 16284 0 1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_20_173
timestamp 1667941163
transform 1 0 17020 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_185
timestamp 1667941163
transform 1 0 18124 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_193
timestamp 1667941163
transform 1 0 18860 0 1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_20_197
timestamp 1667941163
transform 1 0 19228 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_209
timestamp 1667941163
transform 1 0 20332 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_221
timestamp 1667941163
transform 1 0 21436 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_233
timestamp 1667941163
transform 1 0 22540 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_245
timestamp 1667941163
transform 1 0 23644 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_251
timestamp 1667941163
transform 1 0 24196 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_253
timestamp 1667941163
transform 1 0 24380 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_265
timestamp 1667941163
transform 1 0 25484 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_273
timestamp 1667941163
transform 1 0 26220 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_297
timestamp 1667941163
transform 1 0 28428 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_3
timestamp 1667941163
transform 1 0 1380 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_9
timestamp 1667941163
transform 1 0 1932 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_16
timestamp 1667941163
transform 1 0 2576 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_28
timestamp 1667941163
transform 1 0 3680 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_40
timestamp 1667941163
transform 1 0 4784 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_52
timestamp 1667941163
transform 1 0 5888 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_57
timestamp 1667941163
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_69
timestamp 1667941163
transform 1 0 7452 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_77
timestamp 1667941163
transform 1 0 8188 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_99
timestamp 1667941163
transform 1 0 10212 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_110
timestamp 1667941163
transform 1 0 11224 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_113
timestamp 1667941163
transform 1 0 11500 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_136
timestamp 1667941163
transform 1 0 13616 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_142
timestamp 1667941163
transform 1 0 14168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_150
timestamp 1667941163
transform 1 0 14904 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_159
timestamp 1667941163
transform 1 0 15732 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_166
timestamp 1667941163
transform 1 0 16376 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_169
timestamp 1667941163
transform 1 0 16652 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_180
timestamp 1667941163
transform 1 0 17664 0 -1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_21_202
timestamp 1667941163
transform 1 0 19688 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_214
timestamp 1667941163
transform 1 0 20792 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_222
timestamp 1667941163
transform 1 0 21528 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_225
timestamp 1667941163
transform 1 0 21804 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_243
timestamp 1667941163
transform 1 0 23460 0 -1 14144
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_21_267
timestamp 1667941163
transform 1 0 25668 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_21_279
timestamp 1667941163
transform 1 0 26772 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_281
timestamp 1667941163
transform 1 0 26956 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_286
timestamp 1667941163
transform 1 0 27416 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_297
timestamp 1667941163
transform 1 0 28428 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_3
timestamp 1667941163
transform 1 0 1380 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_26
timestamp 1667941163
transform 1 0 3496 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_29
timestamp 1667941163
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_41
timestamp 1667941163
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_53
timestamp 1667941163
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_65
timestamp 1667941163
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_77
timestamp 1667941163
transform 1 0 8188 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_82
timestamp 1667941163
transform 1 0 8648 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_22_85
timestamp 1667941163
transform 1 0 8924 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_91
timestamp 1667941163
transform 1 0 9476 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_113
timestamp 1667941163
transform 1 0 11500 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_22_124
timestamp 1667941163
transform 1 0 12512 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_134
timestamp 1667941163
transform 1 0 13432 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_22_141
timestamp 1667941163
transform 1 0 14076 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_151
timestamp 1667941163
transform 1 0 14996 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_155
timestamp 1667941163
transform 1 0 15364 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_162
timestamp 1667941163
transform 1 0 16008 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_170
timestamp 1667941163
transform 1 0 16744 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_187
timestamp 1667941163
transform 1 0 18308 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_194
timestamp 1667941163
transform 1 0 18952 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_197
timestamp 1667941163
transform 1 0 19228 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_215
timestamp 1667941163
transform 1 0 20884 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_22_235
timestamp 1667941163
transform 1 0 22724 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_247
timestamp 1667941163
transform 1 0 23828 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_251
timestamp 1667941163
transform 1 0 24196 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_253
timestamp 1667941163
transform 1 0 24380 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_272
timestamp 1667941163
transform 1 0 26128 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_297
timestamp 1667941163
transform 1 0 28428 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_3
timestamp 1667941163
transform 1 0 1380 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_7
timestamp 1667941163
transform 1 0 1748 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_11
timestamp 1667941163
transform 1 0 2116 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_23
timestamp 1667941163
transform 1 0 3220 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_35
timestamp 1667941163
transform 1 0 4324 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_47
timestamp 1667941163
transform 1 0 5428 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1667941163
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_57
timestamp 1667941163
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_69
timestamp 1667941163
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_81
timestamp 1667941163
transform 1 0 8556 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_93
timestamp 1667941163
transform 1 0 9660 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_105
timestamp 1667941163
transform 1 0 10764 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp 1667941163
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_113
timestamp 1667941163
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_125
timestamp 1667941163
transform 1 0 12604 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_131
timestamp 1667941163
transform 1 0 13156 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_137
timestamp 1667941163
transform 1 0 13708 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_141
timestamp 1667941163
transform 1 0 14076 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_146
timestamp 1667941163
transform 1 0 14536 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_154
timestamp 1667941163
transform 1 0 15272 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_166
timestamp 1667941163
transform 1 0 16376 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_169
timestamp 1667941163
transform 1 0 16652 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_174
timestamp 1667941163
transform 1 0 17112 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_186
timestamp 1667941163
transform 1 0 18216 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_194
timestamp 1667941163
transform 1 0 18952 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_211
timestamp 1667941163
transform 1 0 20516 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_223
timestamp 1667941163
transform 1 0 21620 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_23_225
timestamp 1667941163
transform 1 0 21804 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_231
timestamp 1667941163
transform 1 0 22356 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_248
timestamp 1667941163
transform 1 0 23920 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_260
timestamp 1667941163
transform 1 0 25024 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_272
timestamp 1667941163
transform 1 0 26128 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_281
timestamp 1667941163
transform 1 0 26956 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_287
timestamp 1667941163
transform 1 0 27508 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_294
timestamp 1667941163
transform 1 0 28152 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_298
timestamp 1667941163
transform 1 0 28520 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_24_3
timestamp 1667941163
transform 1 0 1380 0 1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_24_9
timestamp 1667941163
transform 1 0 1932 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_21
timestamp 1667941163
transform 1 0 3036 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1667941163
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_29
timestamp 1667941163
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_41
timestamp 1667941163
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_53
timestamp 1667941163
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_65
timestamp 1667941163
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_77
timestamp 1667941163
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1667941163
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_85
timestamp 1667941163
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_97
timestamp 1667941163
transform 1 0 10028 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_109
timestamp 1667941163
transform 1 0 11132 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_121
timestamp 1667941163
transform 1 0 12236 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_24_133
timestamp 1667941163
transform 1 0 13340 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_138
timestamp 1667941163
transform 1 0 13800 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_141
timestamp 1667941163
transform 1 0 14076 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_148
timestamp 1667941163
transform 1 0 14720 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_156
timestamp 1667941163
transform 1 0 15456 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_163
timestamp 1667941163
transform 1 0 16100 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_175
timestamp 1667941163
transform 1 0 17204 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_187
timestamp 1667941163
transform 1 0 18308 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_195
timestamp 1667941163
transform 1 0 19044 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_197
timestamp 1667941163
transform 1 0 19228 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_205
timestamp 1667941163
transform 1 0 19964 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_215
timestamp 1667941163
transform 1 0 20884 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_24_228
timestamp 1667941163
transform 1 0 22080 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_240
timestamp 1667941163
transform 1 0 23184 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_253
timestamp 1667941163
transform 1 0 24380 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_261
timestamp 1667941163
transform 1 0 25116 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_272
timestamp 1667941163
transform 1 0 26128 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_297
timestamp 1667941163
transform 1 0 28428 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_3
timestamp 1667941163
transform 1 0 1380 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_25_27
timestamp 1667941163
transform 1 0 3588 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_39
timestamp 1667941163
transform 1 0 4692 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_51
timestamp 1667941163
transform 1 0 5796 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_55
timestamp 1667941163
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_57
timestamp 1667941163
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_69
timestamp 1667941163
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_81
timestamp 1667941163
transform 1 0 8556 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_93
timestamp 1667941163
transform 1 0 9660 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_105
timestamp 1667941163
transform 1 0 10764 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp 1667941163
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_113
timestamp 1667941163
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_125
timestamp 1667941163
transform 1 0 12604 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_137
timestamp 1667941163
transform 1 0 13708 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_25_145
timestamp 1667941163
transform 1 0 14444 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_157
timestamp 1667941163
transform 1 0 15548 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_164
timestamp 1667941163
transform 1 0 16192 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_25_169
timestamp 1667941163
transform 1 0 16652 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_181
timestamp 1667941163
transform 1 0 17756 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_193
timestamp 1667941163
transform 1 0 18860 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_214
timestamp 1667941163
transform 1 0 20792 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_222
timestamp 1667941163
transform 1 0 21528 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_225
timestamp 1667941163
transform 1 0 21804 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_236
timestamp 1667941163
transform 1 0 22816 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_248
timestamp 1667941163
transform 1 0 23920 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_254
timestamp 1667941163
transform 1 0 24472 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_258
timestamp 1667941163
transform 1 0 24840 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_278
timestamp 1667941163
transform 1 0 26680 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_281
timestamp 1667941163
transform 1 0 26956 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_285
timestamp 1667941163
transform 1 0 27324 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_289
timestamp 1667941163
transform 1 0 27692 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_25_296
timestamp 1667941163
transform 1 0 28336 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_26_3
timestamp 1667941163
transform 1 0 1380 0 1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_26_12
timestamp 1667941163
transform 1 0 2208 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_24
timestamp 1667941163
transform 1 0 3312 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_26_29
timestamp 1667941163
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_41
timestamp 1667941163
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_53
timestamp 1667941163
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_65
timestamp 1667941163
transform 1 0 7084 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_77
timestamp 1667941163
transform 1 0 8188 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 1667941163
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_85
timestamp 1667941163
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_97
timestamp 1667941163
transform 1 0 10028 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_109
timestamp 1667941163
transform 1 0 11132 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_121
timestamp 1667941163
transform 1 0 12236 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_26_129
timestamp 1667941163
transform 1 0 12972 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_138
timestamp 1667941163
transform 1 0 13800 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_141
timestamp 1667941163
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_153
timestamp 1667941163
transform 1 0 15180 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_165
timestamp 1667941163
transform 1 0 16284 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_26_187
timestamp 1667941163
transform 1 0 18308 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_194
timestamp 1667941163
transform 1 0 18952 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_197
timestamp 1667941163
transform 1 0 19228 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_203
timestamp 1667941163
transform 1 0 19780 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_211
timestamp 1667941163
transform 1 0 20516 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_222
timestamp 1667941163
transform 1 0 21528 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_242
timestamp 1667941163
transform 1 0 23368 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_26_249
timestamp 1667941163
transform 1 0 24012 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_253
timestamp 1667941163
transform 1 0 24380 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_259
timestamp 1667941163
transform 1 0 24932 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_263
timestamp 1667941163
transform 1 0 25300 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_269
timestamp 1667941163
transform 1 0 25852 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_26_281
timestamp 1667941163
transform 1 0 26956 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_286
timestamp 1667941163
transform 1 0 27416 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_293
timestamp 1667941163
transform 1 0 28060 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_27_3
timestamp 1667941163
transform 1 0 1380 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_7
timestamp 1667941163
transform 1 0 1748 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_11
timestamp 1667941163
transform 1 0 2116 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_23
timestamp 1667941163
transform 1 0 3220 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_35
timestamp 1667941163
transform 1 0 4324 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_47
timestamp 1667941163
transform 1 0 5428 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_55
timestamp 1667941163
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_57
timestamp 1667941163
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_69
timestamp 1667941163
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_81
timestamp 1667941163
transform 1 0 8556 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_93
timestamp 1667941163
transform 1 0 9660 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_105
timestamp 1667941163
transform 1 0 10764 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_111
timestamp 1667941163
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_113
timestamp 1667941163
transform 1 0 11500 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_125
timestamp 1667941163
transform 1 0 12604 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_137
timestamp 1667941163
transform 1 0 13708 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_149
timestamp 1667941163
transform 1 0 14812 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_157
timestamp 1667941163
transform 1 0 15548 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_165
timestamp 1667941163
transform 1 0 16284 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_169
timestamp 1667941163
transform 1 0 16652 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_27_174
timestamp 1667941163
transform 1 0 17112 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_180
timestamp 1667941163
transform 1 0 17664 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_184
timestamp 1667941163
transform 1 0 18032 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_196
timestamp 1667941163
transform 1 0 19136 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_27_205
timestamp 1667941163
transform 1 0 19964 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_217
timestamp 1667941163
transform 1 0 21068 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_223
timestamp 1667941163
transform 1 0 21620 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_225
timestamp 1667941163
transform 1 0 21804 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_232
timestamp 1667941163
transform 1 0 22448 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_239
timestamp 1667941163
transform 1 0 23092 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_243
timestamp 1667941163
transform 1 0 23460 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_261
timestamp 1667941163
transform 1 0 25116 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_271
timestamp 1667941163
transform 1 0 26036 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_278
timestamp 1667941163
transform 1 0 26680 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_281
timestamp 1667941163
transform 1 0 26956 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_27_292
timestamp 1667941163
transform 1 0 27968 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_298
timestamp 1667941163
transform 1 0 28520 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_3
timestamp 1667941163
transform 1 0 1380 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_26
timestamp 1667941163
transform 1 0 3496 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_29
timestamp 1667941163
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_41
timestamp 1667941163
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_53
timestamp 1667941163
transform 1 0 5980 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_65
timestamp 1667941163
transform 1 0 7084 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_77
timestamp 1667941163
transform 1 0 8188 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_83
timestamp 1667941163
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_85
timestamp 1667941163
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_97
timestamp 1667941163
transform 1 0 10028 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_109
timestamp 1667941163
transform 1 0 11132 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_121
timestamp 1667941163
transform 1 0 12236 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_133
timestamp 1667941163
transform 1 0 13340 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_139
timestamp 1667941163
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_141
timestamp 1667941163
transform 1 0 14076 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_28_153
timestamp 1667941163
transform 1 0 15180 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_28_164
timestamp 1667941163
transform 1 0 16192 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_170
timestamp 1667941163
transform 1 0 16744 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_178
timestamp 1667941163
transform 1 0 17480 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_28_193
timestamp 1667941163
transform 1 0 18860 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_197
timestamp 1667941163
transform 1 0 19228 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_203
timestamp 1667941163
transform 1 0 19780 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_215
timestamp 1667941163
transform 1 0 20884 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_227
timestamp 1667941163
transform 1 0 21988 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_235
timestamp 1667941163
transform 1 0 22724 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_244
timestamp 1667941163
transform 1 0 23552 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_253
timestamp 1667941163
transform 1 0 24380 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_272
timestamp 1667941163
transform 1 0 26128 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_297
timestamp 1667941163
transform 1 0 28428 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_3
timestamp 1667941163
transform 1 0 1380 0 -1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_29_9
timestamp 1667941163
transform 1 0 1932 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_21
timestamp 1667941163
transform 1 0 3036 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_33
timestamp 1667941163
transform 1 0 4140 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_45
timestamp 1667941163
transform 1 0 5244 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_53
timestamp 1667941163
transform 1 0 5980 0 -1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_29_57
timestamp 1667941163
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_69
timestamp 1667941163
transform 1 0 7452 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_81
timestamp 1667941163
transform 1 0 8556 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_93
timestamp 1667941163
transform 1 0 9660 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_105
timestamp 1667941163
transform 1 0 10764 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_111
timestamp 1667941163
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_113
timestamp 1667941163
transform 1 0 11500 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_125
timestamp 1667941163
transform 1 0 12604 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_137
timestamp 1667941163
transform 1 0 13708 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_149
timestamp 1667941163
transform 1 0 14812 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_157
timestamp 1667941163
transform 1 0 15548 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_163
timestamp 1667941163
transform 1 0 16100 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_167
timestamp 1667941163
transform 1 0 16468 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_169
timestamp 1667941163
transform 1 0 16652 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_29_180
timestamp 1667941163
transform 1 0 17664 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_29_206
timestamp 1667941163
transform 1 0 20056 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_29_219
timestamp 1667941163
transform 1 0 21252 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_223
timestamp 1667941163
transform 1 0 21620 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_225
timestamp 1667941163
transform 1 0 21804 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_233
timestamp 1667941163
transform 1 0 22540 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_238
timestamp 1667941163
transform 1 0 23000 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_29_262
timestamp 1667941163
transform 1 0 25208 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_274
timestamp 1667941163
transform 1 0 26312 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_29_281
timestamp 1667941163
transform 1 0 26956 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_288
timestamp 1667941163
transform 1 0 27600 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_295
timestamp 1667941163
transform 1 0 28244 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_3
timestamp 1667941163
transform 1 0 1380 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_8
timestamp 1667941163
transform 1 0 1840 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_20
timestamp 1667941163
transform 1 0 2944 0 1 18496
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_30_29
timestamp 1667941163
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_41
timestamp 1667941163
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_53
timestamp 1667941163
transform 1 0 5980 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_65
timestamp 1667941163
transform 1 0 7084 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_77
timestamp 1667941163
transform 1 0 8188 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_83
timestamp 1667941163
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_85
timestamp 1667941163
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_97
timestamp 1667941163
transform 1 0 10028 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_109
timestamp 1667941163
transform 1 0 11132 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_121
timestamp 1667941163
transform 1 0 12236 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_133
timestamp 1667941163
transform 1 0 13340 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_139
timestamp 1667941163
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_141
timestamp 1667941163
transform 1 0 14076 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_153
timestamp 1667941163
transform 1 0 15180 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_165
timestamp 1667941163
transform 1 0 16284 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_30_178
timestamp 1667941163
transform 1 0 17480 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_185
timestamp 1667941163
transform 1 0 18124 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_192
timestamp 1667941163
transform 1 0 18768 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_197
timestamp 1667941163
transform 1 0 19228 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_30_202
timestamp 1667941163
transform 1 0 19688 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_30_231
timestamp 1667941163
transform 1 0 22356 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_239
timestamp 1667941163
transform 1 0 23092 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_247
timestamp 1667941163
transform 1 0 23828 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_251
timestamp 1667941163
transform 1 0 24196 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_253
timestamp 1667941163
transform 1 0 24380 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_259
timestamp 1667941163
transform 1 0 24932 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_30_271
timestamp 1667941163
transform 1 0 26036 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_290
timestamp 1667941163
transform 1 0 27784 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_297
timestamp 1667941163
transform 1 0 28428 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_3
timestamp 1667941163
transform 1 0 1380 0 -1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_31_9
timestamp 1667941163
transform 1 0 1932 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_21
timestamp 1667941163
transform 1 0 3036 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_33
timestamp 1667941163
transform 1 0 4140 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_45
timestamp 1667941163
transform 1 0 5244 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_53
timestamp 1667941163
transform 1 0 5980 0 -1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_31_57
timestamp 1667941163
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_69
timestamp 1667941163
transform 1 0 7452 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_81
timestamp 1667941163
transform 1 0 8556 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_93
timestamp 1667941163
transform 1 0 9660 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_105
timestamp 1667941163
transform 1 0 10764 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_111
timestamp 1667941163
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_113
timestamp 1667941163
transform 1 0 11500 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_125
timestamp 1667941163
transform 1 0 12604 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_137
timestamp 1667941163
transform 1 0 13708 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_149
timestamp 1667941163
transform 1 0 14812 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_161
timestamp 1667941163
transform 1 0 15916 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_166
timestamp 1667941163
transform 1 0 16376 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_169
timestamp 1667941163
transform 1 0 16652 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_31_175
timestamp 1667941163
transform 1 0 17204 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_181
timestamp 1667941163
transform 1 0 17756 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_187
timestamp 1667941163
transform 1 0 18308 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_198
timestamp 1667941163
transform 1 0 19320 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_208
timestamp 1667941163
transform 1 0 20240 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_215
timestamp 1667941163
transform 1 0 20884 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_222
timestamp 1667941163
transform 1 0 21528 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_225
timestamp 1667941163
transform 1 0 21804 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_244
timestamp 1667941163
transform 1 0 23552 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_31_256
timestamp 1667941163
transform 1 0 24656 0 -1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_31_267
timestamp 1667941163
transform 1 0 25668 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_31_279
timestamp 1667941163
transform 1 0 26772 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_31_281
timestamp 1667941163
transform 1 0 26956 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_287
timestamp 1667941163
transform 1 0 27508 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_294
timestamp 1667941163
transform 1 0 28152 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_298
timestamp 1667941163
transform 1 0 28520 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_3
timestamp 1667941163
transform 1 0 1380 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_26
timestamp 1667941163
transform 1 0 3496 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_29
timestamp 1667941163
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_41
timestamp 1667941163
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_53
timestamp 1667941163
transform 1 0 5980 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_65
timestamp 1667941163
transform 1 0 7084 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_77
timestamp 1667941163
transform 1 0 8188 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_83
timestamp 1667941163
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_85
timestamp 1667941163
transform 1 0 8924 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_97
timestamp 1667941163
transform 1 0 10028 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_109
timestamp 1667941163
transform 1 0 11132 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_121
timestamp 1667941163
transform 1 0 12236 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_133
timestamp 1667941163
transform 1 0 13340 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_139
timestamp 1667941163
transform 1 0 13892 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_141
timestamp 1667941163
transform 1 0 14076 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_162
timestamp 1667941163
transform 1 0 16008 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_174
timestamp 1667941163
transform 1 0 17112 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_186
timestamp 1667941163
transform 1 0 18216 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_194
timestamp 1667941163
transform 1 0 18952 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_197
timestamp 1667941163
transform 1 0 19228 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_209
timestamp 1667941163
transform 1 0 20332 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_229
timestamp 1667941163
transform 1 0 22172 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_241
timestamp 1667941163
transform 1 0 23276 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_32_249
timestamp 1667941163
transform 1 0 24012 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_253
timestamp 1667941163
transform 1 0 24380 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_263
timestamp 1667941163
transform 1 0 25300 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_275
timestamp 1667941163
transform 1 0 26404 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_297
timestamp 1667941163
transform 1 0 28428 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_3
timestamp 1667941163
transform 1 0 1380 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_10
timestamp 1667941163
transform 1 0 2024 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_22
timestamp 1667941163
transform 1 0 3128 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_34
timestamp 1667941163
transform 1 0 4232 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_46
timestamp 1667941163
transform 1 0 5336 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_54
timestamp 1667941163
transform 1 0 6072 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_57
timestamp 1667941163
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_69
timestamp 1667941163
transform 1 0 7452 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_81
timestamp 1667941163
transform 1 0 8556 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_93
timestamp 1667941163
transform 1 0 9660 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_105
timestamp 1667941163
transform 1 0 10764 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_111
timestamp 1667941163
transform 1 0 11316 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_113
timestamp 1667941163
transform 1 0 11500 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_125
timestamp 1667941163
transform 1 0 12604 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_137
timestamp 1667941163
transform 1 0 13708 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_149
timestamp 1667941163
transform 1 0 14812 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_155
timestamp 1667941163
transform 1 0 15364 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_161
timestamp 1667941163
transform 1 0 15916 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_167
timestamp 1667941163
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_169
timestamp 1667941163
transform 1 0 16652 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_187
timestamp 1667941163
transform 1 0 18308 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_195
timestamp 1667941163
transform 1 0 19044 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_213
timestamp 1667941163
transform 1 0 20700 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_33_221
timestamp 1667941163
transform 1 0 21436 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_33_225
timestamp 1667941163
transform 1 0 21804 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_237
timestamp 1667941163
transform 1 0 22908 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_249
timestamp 1667941163
transform 1 0 24012 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_33_261
timestamp 1667941163
transform 1 0 25116 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_278
timestamp 1667941163
transform 1 0 26680 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_281
timestamp 1667941163
transform 1 0 26956 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_287
timestamp 1667941163
transform 1 0 27508 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_294
timestamp 1667941163
transform 1 0 28152 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_298
timestamp 1667941163
transform 1 0 28520 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_3
timestamp 1667941163
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_15
timestamp 1667941163
transform 1 0 2484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 1667941163
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_29
timestamp 1667941163
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_41
timestamp 1667941163
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_53
timestamp 1667941163
transform 1 0 5980 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_65
timestamp 1667941163
transform 1 0 7084 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_77
timestamp 1667941163
transform 1 0 8188 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_83
timestamp 1667941163
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_85
timestamp 1667941163
transform 1 0 8924 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_97
timestamp 1667941163
transform 1 0 10028 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_109
timestamp 1667941163
transform 1 0 11132 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_121
timestamp 1667941163
transform 1 0 12236 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_133
timestamp 1667941163
transform 1 0 13340 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_139
timestamp 1667941163
transform 1 0 13892 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_141
timestamp 1667941163
transform 1 0 14076 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_153
timestamp 1667941163
transform 1 0 15180 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_161
timestamp 1667941163
transform 1 0 15916 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_165
timestamp 1667941163
transform 1 0 16284 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_177
timestamp 1667941163
transform 1 0 17388 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_34_189
timestamp 1667941163
transform 1 0 18492 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_194
timestamp 1667941163
transform 1 0 18952 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_197
timestamp 1667941163
transform 1 0 19228 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_204
timestamp 1667941163
transform 1 0 19872 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_217
timestamp 1667941163
transform 1 0 21068 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_225
timestamp 1667941163
transform 1 0 21804 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_34_243
timestamp 1667941163
transform 1 0 23460 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_251
timestamp 1667941163
transform 1 0 24196 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_253
timestamp 1667941163
transform 1 0 24380 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_265
timestamp 1667941163
transform 1 0 25484 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_34_273
timestamp 1667941163
transform 1 0 26220 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_34_297
timestamp 1667941163
transform 1 0 28428 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_3
timestamp 1667941163
transform 1 0 1380 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_15
timestamp 1667941163
transform 1 0 2484 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_27
timestamp 1667941163
transform 1 0 3588 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_39
timestamp 1667941163
transform 1 0 4692 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_51
timestamp 1667941163
transform 1 0 5796 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_55
timestamp 1667941163
transform 1 0 6164 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_57
timestamp 1667941163
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_69
timestamp 1667941163
transform 1 0 7452 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_81
timestamp 1667941163
transform 1 0 8556 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_93
timestamp 1667941163
transform 1 0 9660 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_105
timestamp 1667941163
transform 1 0 10764 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_111
timestamp 1667941163
transform 1 0 11316 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_113
timestamp 1667941163
transform 1 0 11500 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_125
timestamp 1667941163
transform 1 0 12604 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_137
timestamp 1667941163
transform 1 0 13708 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_149
timestamp 1667941163
transform 1 0 14812 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_161
timestamp 1667941163
transform 1 0 15916 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_167
timestamp 1667941163
transform 1 0 16468 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_169
timestamp 1667941163
transform 1 0 16652 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_187
timestamp 1667941163
transform 1 0 18308 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_205
timestamp 1667941163
transform 1 0 19964 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_35_216
timestamp 1667941163
transform 1 0 20976 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_35_225
timestamp 1667941163
transform 1 0 21804 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_229
timestamp 1667941163
transform 1 0 22172 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_238
timestamp 1667941163
transform 1 0 23000 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_244
timestamp 1667941163
transform 1 0 23552 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_252
timestamp 1667941163
transform 1 0 24288 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_258
timestamp 1667941163
transform 1 0 24840 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_266
timestamp 1667941163
transform 1 0 25576 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_35_278
timestamp 1667941163
transform 1 0 26680 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_281
timestamp 1667941163
transform 1 0 26956 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_286
timestamp 1667941163
transform 1 0 27416 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_293
timestamp 1667941163
transform 1 0 28060 0 -1 21760
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_36_3
timestamp 1667941163
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_15
timestamp 1667941163
transform 1 0 2484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 1667941163
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_29
timestamp 1667941163
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_41
timestamp 1667941163
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_53
timestamp 1667941163
transform 1 0 5980 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_65
timestamp 1667941163
transform 1 0 7084 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_77
timestamp 1667941163
transform 1 0 8188 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_83
timestamp 1667941163
transform 1 0 8740 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_85
timestamp 1667941163
transform 1 0 8924 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_97
timestamp 1667941163
transform 1 0 10028 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_109
timestamp 1667941163
transform 1 0 11132 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_121
timestamp 1667941163
transform 1 0 12236 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_133
timestamp 1667941163
transform 1 0 13340 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_139
timestamp 1667941163
transform 1 0 13892 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_141
timestamp 1667941163
transform 1 0 14076 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_153
timestamp 1667941163
transform 1 0 15180 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_161
timestamp 1667941163
transform 1 0 15916 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_165
timestamp 1667941163
transform 1 0 16284 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_177
timestamp 1667941163
transform 1 0 17388 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_189
timestamp 1667941163
transform 1 0 18492 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_195
timestamp 1667941163
transform 1 0 19044 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_197
timestamp 1667941163
transform 1 0 19228 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_205
timestamp 1667941163
transform 1 0 19964 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_209
timestamp 1667941163
transform 1 0 20332 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_226
timestamp 1667941163
transform 1 0 21896 0 1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_36_234
timestamp 1667941163
transform 1 0 22632 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_246
timestamp 1667941163
transform 1 0 23736 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_250
timestamp 1667941163
transform 1 0 24104 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_253
timestamp 1667941163
transform 1 0 24380 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_36_263
timestamp 1667941163
transform 1 0 25300 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_275
timestamp 1667941163
transform 1 0 26404 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_297
timestamp 1667941163
transform 1 0 28428 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_3
timestamp 1667941163
transform 1 0 1380 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_15
timestamp 1667941163
transform 1 0 2484 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_27
timestamp 1667941163
transform 1 0 3588 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_39
timestamp 1667941163
transform 1 0 4692 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_51
timestamp 1667941163
transform 1 0 5796 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_55
timestamp 1667941163
transform 1 0 6164 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_57
timestamp 1667941163
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_69
timestamp 1667941163
transform 1 0 7452 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_81
timestamp 1667941163
transform 1 0 8556 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_93
timestamp 1667941163
transform 1 0 9660 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_105
timestamp 1667941163
transform 1 0 10764 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_111
timestamp 1667941163
transform 1 0 11316 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_113
timestamp 1667941163
transform 1 0 11500 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_125
timestamp 1667941163
transform 1 0 12604 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_137
timestamp 1667941163
transform 1 0 13708 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_149
timestamp 1667941163
transform 1 0 14812 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_161
timestamp 1667941163
transform 1 0 15916 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_167
timestamp 1667941163
transform 1 0 16468 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_169
timestamp 1667941163
transform 1 0 16652 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_37_179
timestamp 1667941163
transform 1 0 17572 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_187
timestamp 1667941163
transform 1 0 18308 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_197
timestamp 1667941163
transform 1 0 19228 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_204
timestamp 1667941163
transform 1 0 19872 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_212
timestamp 1667941163
transform 1 0 20608 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_222
timestamp 1667941163
transform 1 0 21528 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_37_225
timestamp 1667941163
transform 1 0 21804 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_233
timestamp 1667941163
transform 1 0 22540 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_37_238
timestamp 1667941163
transform 1 0 23000 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_244
timestamp 1667941163
transform 1 0 23552 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_253
timestamp 1667941163
transform 1 0 24380 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_278
timestamp 1667941163
transform 1 0 26680 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_281
timestamp 1667941163
transform 1 0 26956 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_286
timestamp 1667941163
transform 1 0 27416 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_290
timestamp 1667941163
transform 1 0 27784 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_294
timestamp 1667941163
transform 1 0 28152 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_298
timestamp 1667941163
transform 1 0 28520 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_3
timestamp 1667941163
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_15
timestamp 1667941163
transform 1 0 2484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 1667941163
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_29
timestamp 1667941163
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_41
timestamp 1667941163
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_53
timestamp 1667941163
transform 1 0 5980 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_65
timestamp 1667941163
transform 1 0 7084 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_77
timestamp 1667941163
transform 1 0 8188 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_83
timestamp 1667941163
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_85
timestamp 1667941163
transform 1 0 8924 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_97
timestamp 1667941163
transform 1 0 10028 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_109
timestamp 1667941163
transform 1 0 11132 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_121
timestamp 1667941163
transform 1 0 12236 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_133
timestamp 1667941163
transform 1 0 13340 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_139
timestamp 1667941163
transform 1 0 13892 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_141
timestamp 1667941163
transform 1 0 14076 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_153
timestamp 1667941163
transform 1 0 15180 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_157
timestamp 1667941163
transform 1 0 15548 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_161
timestamp 1667941163
transform 1 0 15916 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_170
timestamp 1667941163
transform 1 0 16744 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_174
timestamp 1667941163
transform 1 0 17112 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_183
timestamp 1667941163
transform 1 0 17940 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_190
timestamp 1667941163
transform 1 0 18584 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_38_197
timestamp 1667941163
transform 1 0 19228 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_38_204
timestamp 1667941163
transform 1 0 19872 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_210
timestamp 1667941163
transform 1 0 20424 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_216
timestamp 1667941163
transform 1 0 20976 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_228
timestamp 1667941163
transform 1 0 22080 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_38_240
timestamp 1667941163
transform 1 0 23184 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_38_247
timestamp 1667941163
transform 1 0 23828 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_251
timestamp 1667941163
transform 1 0 24196 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_38_253
timestamp 1667941163
transform 1 0 24380 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_38_266
timestamp 1667941163
transform 1 0 25576 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_274
timestamp 1667941163
transform 1 0 26312 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_297
timestamp 1667941163
transform 1 0 28428 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_39_3
timestamp 1667941163
transform 1 0 1380 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_15
timestamp 1667941163
transform 1 0 2484 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_27
timestamp 1667941163
transform 1 0 3588 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_39
timestamp 1667941163
transform 1 0 4692 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_51
timestamp 1667941163
transform 1 0 5796 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_55
timestamp 1667941163
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_57
timestamp 1667941163
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_69
timestamp 1667941163
transform 1 0 7452 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_81
timestamp 1667941163
transform 1 0 8556 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_93
timestamp 1667941163
transform 1 0 9660 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_105
timestamp 1667941163
transform 1 0 10764 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_111
timestamp 1667941163
transform 1 0 11316 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_113
timestamp 1667941163
transform 1 0 11500 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_125
timestamp 1667941163
transform 1 0 12604 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_137
timestamp 1667941163
transform 1 0 13708 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_149
timestamp 1667941163
transform 1 0 14812 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_161
timestamp 1667941163
transform 1 0 15916 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_167
timestamp 1667941163
transform 1 0 16468 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_39_169
timestamp 1667941163
transform 1 0 16652 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_175
timestamp 1667941163
transform 1 0 17204 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_181
timestamp 1667941163
transform 1 0 17756 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_188
timestamp 1667941163
transform 1 0 18400 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_195
timestamp 1667941163
transform 1 0 19044 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_201
timestamp 1667941163
transform 1 0 19596 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_205
timestamp 1667941163
transform 1 0 19964 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_209
timestamp 1667941163
transform 1 0 20332 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_219
timestamp 1667941163
transform 1 0 21252 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_223
timestamp 1667941163
transform 1 0 21620 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_225
timestamp 1667941163
transform 1 0 21804 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_237
timestamp 1667941163
transform 1 0 22908 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_249
timestamp 1667941163
transform 1 0 24012 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_261
timestamp 1667941163
transform 1 0 25116 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_39_273
timestamp 1667941163
transform 1 0 26220 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_278
timestamp 1667941163
transform 1 0 26680 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_39_281
timestamp 1667941163
transform 1 0 26956 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_39_287
timestamp 1667941163
transform 1 0 27508 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_294
timestamp 1667941163
transform 1 0 28152 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_298
timestamp 1667941163
transform 1 0 28520 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_3
timestamp 1667941163
transform 1 0 1380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_15
timestamp 1667941163
transform 1 0 2484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_27
timestamp 1667941163
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_29
timestamp 1667941163
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_41
timestamp 1667941163
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_53
timestamp 1667941163
transform 1 0 5980 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_65
timestamp 1667941163
transform 1 0 7084 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_77
timestamp 1667941163
transform 1 0 8188 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_83
timestamp 1667941163
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_85
timestamp 1667941163
transform 1 0 8924 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_97
timestamp 1667941163
transform 1 0 10028 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_109
timestamp 1667941163
transform 1 0 11132 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_121
timestamp 1667941163
transform 1 0 12236 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_133
timestamp 1667941163
transform 1 0 13340 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_139
timestamp 1667941163
transform 1 0 13892 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_141
timestamp 1667941163
transform 1 0 14076 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_153
timestamp 1667941163
transform 1 0 15180 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_165
timestamp 1667941163
transform 1 0 16284 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_173
timestamp 1667941163
transform 1 0 17020 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_177
timestamp 1667941163
transform 1 0 17388 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_189
timestamp 1667941163
transform 1 0 18492 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_195
timestamp 1667941163
transform 1 0 19044 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_197
timestamp 1667941163
transform 1 0 19228 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_40_215
timestamp 1667941163
transform 1 0 20884 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_40_239
timestamp 1667941163
transform 1 0 23092 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_248
timestamp 1667941163
transform 1 0 23920 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_40_253
timestamp 1667941163
transform 1 0 24380 0 1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_40_259
timestamp 1667941163
transform 1 0 24932 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_271
timestamp 1667941163
transform 1 0 26036 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_275
timestamp 1667941163
transform 1 0 26404 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_297
timestamp 1667941163
transform 1 0 28428 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_3
timestamp 1667941163
transform 1 0 1380 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_41_8
timestamp 1667941163
transform 1 0 1840 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_20
timestamp 1667941163
transform 1 0 2944 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_32
timestamp 1667941163
transform 1 0 4048 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_44
timestamp 1667941163
transform 1 0 5152 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_57
timestamp 1667941163
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_69
timestamp 1667941163
transform 1 0 7452 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_81
timestamp 1667941163
transform 1 0 8556 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_93
timestamp 1667941163
transform 1 0 9660 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_105
timestamp 1667941163
transform 1 0 10764 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_111
timestamp 1667941163
transform 1 0 11316 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_113
timestamp 1667941163
transform 1 0 11500 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_125
timestamp 1667941163
transform 1 0 12604 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_137
timestamp 1667941163
transform 1 0 13708 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_149
timestamp 1667941163
transform 1 0 14812 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_161
timestamp 1667941163
transform 1 0 15916 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_167
timestamp 1667941163
transform 1 0 16468 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_169
timestamp 1667941163
transform 1 0 16652 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_41_194
timestamp 1667941163
transform 1 0 18952 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_41_207
timestamp 1667941163
transform 1 0 20148 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_220
timestamp 1667941163
transform 1 0 21344 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_225
timestamp 1667941163
transform 1 0 21804 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_237
timestamp 1667941163
transform 1 0 22908 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_41_250
timestamp 1667941163
transform 1 0 24104 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_41_258
timestamp 1667941163
transform 1 0 24840 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_41_271
timestamp 1667941163
transform 1 0 26036 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_279
timestamp 1667941163
transform 1 0 26772 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_41_281
timestamp 1667941163
transform 1 0 26956 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_286
timestamp 1667941163
transform 1 0 27416 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_41_293
timestamp 1667941163
transform 1 0 28060 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_42_3
timestamp 1667941163
transform 1 0 1380 0 1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_42_9
timestamp 1667941163
transform 1 0 1932 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_21
timestamp 1667941163
transform 1 0 3036 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_27
timestamp 1667941163
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_29
timestamp 1667941163
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_41
timestamp 1667941163
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_53
timestamp 1667941163
transform 1 0 5980 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_65
timestamp 1667941163
transform 1 0 7084 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_77
timestamp 1667941163
transform 1 0 8188 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_83
timestamp 1667941163
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_85
timestamp 1667941163
transform 1 0 8924 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_97
timestamp 1667941163
transform 1 0 10028 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_109
timestamp 1667941163
transform 1 0 11132 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_121
timestamp 1667941163
transform 1 0 12236 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_133
timestamp 1667941163
transform 1 0 13340 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_139
timestamp 1667941163
transform 1 0 13892 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_141
timestamp 1667941163
transform 1 0 14076 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_42_153
timestamp 1667941163
transform 1 0 15180 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_42_165
timestamp 1667941163
transform 1 0 16284 0 1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_42_174
timestamp 1667941163
transform 1 0 17112 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_42_186
timestamp 1667941163
transform 1 0 18216 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_42_192
timestamp 1667941163
transform 1 0 18768 0 1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_42_197
timestamp 1667941163
transform 1 0 19228 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_209
timestamp 1667941163
transform 1 0 20332 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_221
timestamp 1667941163
transform 1 0 21436 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_226
timestamp 1667941163
transform 1 0 21896 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_42_250
timestamp 1667941163
transform 1 0 24104 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_42_253
timestamp 1667941163
transform 1 0 24380 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_259
timestamp 1667941163
transform 1 0 24932 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_42_269
timestamp 1667941163
transform 1 0 25852 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_275
timestamp 1667941163
transform 1 0 26404 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_42_297
timestamp 1667941163
transform 1 0 28428 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_43_3
timestamp 1667941163
transform 1 0 1380 0 -1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_43_27
timestamp 1667941163
transform 1 0 3588 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_39
timestamp 1667941163
transform 1 0 4692 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_51
timestamp 1667941163
transform 1 0 5796 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_55
timestamp 1667941163
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_57
timestamp 1667941163
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_69
timestamp 1667941163
transform 1 0 7452 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_81
timestamp 1667941163
transform 1 0 8556 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_93
timestamp 1667941163
transform 1 0 9660 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_105
timestamp 1667941163
transform 1 0 10764 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_111
timestamp 1667941163
transform 1 0 11316 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_113
timestamp 1667941163
transform 1 0 11500 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_125
timestamp 1667941163
transform 1 0 12604 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_137
timestamp 1667941163
transform 1 0 13708 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_149
timestamp 1667941163
transform 1 0 14812 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_43_161
timestamp 1667941163
transform 1 0 15916 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_166
timestamp 1667941163
transform 1 0 16376 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_169
timestamp 1667941163
transform 1 0 16652 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_43_187
timestamp 1667941163
transform 1 0 18308 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_199
timestamp 1667941163
transform 1 0 19412 0 -1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_43_208
timestamp 1667941163
transform 1 0 20240 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_220
timestamp 1667941163
transform 1 0 21344 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_43_225
timestamp 1667941163
transform 1 0 21804 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_43_233
timestamp 1667941163
transform 1 0 22540 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_43_239
timestamp 1667941163
transform 1 0 23092 0 -1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_43_246
timestamp 1667941163
transform 1 0 23736 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_43_258
timestamp 1667941163
transform 1 0 24840 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_43_267
timestamp 1667941163
transform 1 0 25668 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_271
timestamp 1667941163
transform 1 0 26036 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_43_278
timestamp 1667941163
transform 1 0 26680 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_281
timestamp 1667941163
transform 1 0 26956 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_43_286
timestamp 1667941163
transform 1 0 27416 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_43_298
timestamp 1667941163
transform 1 0 28520 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_44_3
timestamp 1667941163
transform 1 0 1380 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_9
timestamp 1667941163
transform 1 0 1932 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_13
timestamp 1667941163
transform 1 0 2300 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_44_25
timestamp 1667941163
transform 1 0 3404 0 1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_44_29
timestamp 1667941163
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_41
timestamp 1667941163
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_53
timestamp 1667941163
transform 1 0 5980 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_65
timestamp 1667941163
transform 1 0 7084 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_77
timestamp 1667941163
transform 1 0 8188 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_83
timestamp 1667941163
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_85
timestamp 1667941163
transform 1 0 8924 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_97
timestamp 1667941163
transform 1 0 10028 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_109
timestamp 1667941163
transform 1 0 11132 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_121
timestamp 1667941163
transform 1 0 12236 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_133
timestamp 1667941163
transform 1 0 13340 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_139
timestamp 1667941163
transform 1 0 13892 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_141
timestamp 1667941163
transform 1 0 14076 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_44_153
timestamp 1667941163
transform 1 0 15180 0 1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_44_165
timestamp 1667941163
transform 1 0 16284 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_177
timestamp 1667941163
transform 1 0 17388 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_189
timestamp 1667941163
transform 1 0 18492 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_195
timestamp 1667941163
transform 1 0 19044 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_44_197
timestamp 1667941163
transform 1 0 19228 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_44_206
timestamp 1667941163
transform 1 0 20056 0 1 26112
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_44_228
timestamp 1667941163
transform 1 0 22080 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_240
timestamp 1667941163
transform 1 0 23184 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_246
timestamp 1667941163
transform 1 0 23736 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_250
timestamp 1667941163
transform 1 0 24104 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_253
timestamp 1667941163
transform 1 0 24380 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_44_261
timestamp 1667941163
transform 1 0 25116 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_269
timestamp 1667941163
transform 1 0 25852 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_286
timestamp 1667941163
transform 1 0 27416 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_298
timestamp 1667941163
transform 1 0 28520 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_3
timestamp 1667941163
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_15
timestamp 1667941163
transform 1 0 2484 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_27
timestamp 1667941163
transform 1 0 3588 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_39
timestamp 1667941163
transform 1 0 4692 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_51
timestamp 1667941163
transform 1 0 5796 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_55
timestamp 1667941163
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_57
timestamp 1667941163
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_69
timestamp 1667941163
transform 1 0 7452 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_81
timestamp 1667941163
transform 1 0 8556 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_93
timestamp 1667941163
transform 1 0 9660 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_105
timestamp 1667941163
transform 1 0 10764 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_111
timestamp 1667941163
transform 1 0 11316 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_113
timestamp 1667941163
transform 1 0 11500 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_125
timestamp 1667941163
transform 1 0 12604 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_137
timestamp 1667941163
transform 1 0 13708 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_149
timestamp 1667941163
transform 1 0 14812 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_45_166
timestamp 1667941163
transform 1 0 16376 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_169
timestamp 1667941163
transform 1 0 16652 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_189
timestamp 1667941163
transform 1 0 18492 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_209
timestamp 1667941163
transform 1 0 20332 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_45_217
timestamp 1667941163
transform 1 0 21068 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_45_222
timestamp 1667941163
transform 1 0 21528 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_225
timestamp 1667941163
transform 1 0 21804 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_235
timestamp 1667941163
transform 1 0 22724 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_242
timestamp 1667941163
transform 1 0 23368 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_45_250
timestamp 1667941163
transform 1 0 24104 0 -1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_45_257
timestamp 1667941163
transform 1 0 24748 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_269
timestamp 1667941163
transform 1 0 25852 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_45_277
timestamp 1667941163
transform 1 0 26588 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_45_281
timestamp 1667941163
transform 1 0 26956 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_45_292
timestamp 1667941163
transform 1 0 27968 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_298
timestamp 1667941163
transform 1 0 28520 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_3
timestamp 1667941163
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_15
timestamp 1667941163
transform 1 0 2484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_27
timestamp 1667941163
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_29
timestamp 1667941163
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_41
timestamp 1667941163
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_53
timestamp 1667941163
transform 1 0 5980 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_65
timestamp 1667941163
transform 1 0 7084 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_77
timestamp 1667941163
transform 1 0 8188 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_83
timestamp 1667941163
transform 1 0 8740 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_85
timestamp 1667941163
transform 1 0 8924 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_97
timestamp 1667941163
transform 1 0 10028 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_109
timestamp 1667941163
transform 1 0 11132 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_121
timestamp 1667941163
transform 1 0 12236 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_133
timestamp 1667941163
transform 1 0 13340 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_139
timestamp 1667941163
transform 1 0 13892 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_46_141
timestamp 1667941163
transform 1 0 14076 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_46_147
timestamp 1667941163
transform 1 0 14628 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_46_162
timestamp 1667941163
transform 1 0 16008 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_166
timestamp 1667941163
transform 1 0 16376 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_170
timestamp 1667941163
transform 1 0 16744 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_182
timestamp 1667941163
transform 1 0 17848 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_46_194
timestamp 1667941163
transform 1 0 18952 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_197
timestamp 1667941163
transform 1 0 19228 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_46_215
timestamp 1667941163
transform 1 0 20884 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_227
timestamp 1667941163
transform 1 0 21988 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_231
timestamp 1667941163
transform 1 0 22356 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_46_249
timestamp 1667941163
transform 1 0 24012 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_46_253
timestamp 1667941163
transform 1 0 24380 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_46_269
timestamp 1667941163
transform 1 0 25852 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_275
timestamp 1667941163
transform 1 0 26404 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_46_297
timestamp 1667941163
transform 1 0 28428 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_3
timestamp 1667941163
transform 1 0 1380 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_47_8
timestamp 1667941163
transform 1 0 1840 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_20
timestamp 1667941163
transform 1 0 2944 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_32
timestamp 1667941163
transform 1 0 4048 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_44
timestamp 1667941163
transform 1 0 5152 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_57
timestamp 1667941163
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_69
timestamp 1667941163
transform 1 0 7452 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_81
timestamp 1667941163
transform 1 0 8556 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_93
timestamp 1667941163
transform 1 0 9660 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_105
timestamp 1667941163
transform 1 0 10764 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_111
timestamp 1667941163
transform 1 0 11316 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_113
timestamp 1667941163
transform 1 0 11500 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_125
timestamp 1667941163
transform 1 0 12604 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_137
timestamp 1667941163
transform 1 0 13708 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_47_164
timestamp 1667941163
transform 1 0 16192 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_47_169
timestamp 1667941163
transform 1 0 16652 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_47_174
timestamp 1667941163
transform 1 0 17112 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_186
timestamp 1667941163
transform 1 0 18216 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_198
timestamp 1667941163
transform 1 0 19320 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_210
timestamp 1667941163
transform 1 0 20424 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_47_222
timestamp 1667941163
transform 1 0 21528 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_47_225
timestamp 1667941163
transform 1 0 21804 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_47_233
timestamp 1667941163
transform 1 0 22540 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_241
timestamp 1667941163
transform 1 0 23276 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_247
timestamp 1667941163
transform 1 0 23828 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_258
timestamp 1667941163
transform 1 0 24840 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_47_278
timestamp 1667941163
transform 1 0 26680 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_47_281
timestamp 1667941163
transform 1 0 26956 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_47_287
timestamp 1667941163
transform 1 0 27508 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_294
timestamp 1667941163
transform 1 0 28152 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_298
timestamp 1667941163
transform 1 0 28520 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_3
timestamp 1667941163
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_15
timestamp 1667941163
transform 1 0 2484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 1667941163
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_29
timestamp 1667941163
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_41
timestamp 1667941163
transform 1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_53
timestamp 1667941163
transform 1 0 5980 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_65
timestamp 1667941163
transform 1 0 7084 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_77
timestamp 1667941163
transform 1 0 8188 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_83
timestamp 1667941163
transform 1 0 8740 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_85
timestamp 1667941163
transform 1 0 8924 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_97
timestamp 1667941163
transform 1 0 10028 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_109
timestamp 1667941163
transform 1 0 11132 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_121
timestamp 1667941163
transform 1 0 12236 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_133
timestamp 1667941163
transform 1 0 13340 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_139
timestamp 1667941163
transform 1 0 13892 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_141
timestamp 1667941163
transform 1 0 14076 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_153
timestamp 1667941163
transform 1 0 15180 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_157
timestamp 1667941163
transform 1 0 15548 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_48_163
timestamp 1667941163
transform 1 0 16100 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_48_187
timestamp 1667941163
transform 1 0 18308 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_195
timestamp 1667941163
transform 1 0 19044 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_197
timestamp 1667941163
transform 1 0 19228 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_209
timestamp 1667941163
transform 1 0 20332 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_213
timestamp 1667941163
transform 1 0 20700 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_234
timestamp 1667941163
transform 1 0 22632 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_48_242
timestamp 1667941163
transform 1 0 23368 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_48_250
timestamp 1667941163
transform 1 0 24104 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_253
timestamp 1667941163
transform 1 0 24380 0 1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_48_260
timestamp 1667941163
transform 1 0 25024 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_272
timestamp 1667941163
transform 1 0 26128 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_48_297
timestamp 1667941163
transform 1 0 28428 0 1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_49_3
timestamp 1667941163
transform 1 0 1380 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_15
timestamp 1667941163
transform 1 0 2484 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_27
timestamp 1667941163
transform 1 0 3588 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_39
timestamp 1667941163
transform 1 0 4692 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_51
timestamp 1667941163
transform 1 0 5796 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_55
timestamp 1667941163
transform 1 0 6164 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_57
timestamp 1667941163
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_69
timestamp 1667941163
transform 1 0 7452 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_81
timestamp 1667941163
transform 1 0 8556 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_93
timestamp 1667941163
transform 1 0 9660 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_105
timestamp 1667941163
transform 1 0 10764 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_111
timestamp 1667941163
transform 1 0 11316 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_113
timestamp 1667941163
transform 1 0 11500 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_125
timestamp 1667941163
transform 1 0 12604 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_137
timestamp 1667941163
transform 1 0 13708 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_149
timestamp 1667941163
transform 1 0 14812 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_161
timestamp 1667941163
transform 1 0 15916 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_167
timestamp 1667941163
transform 1 0 16468 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_169
timestamp 1667941163
transform 1 0 16652 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_181
timestamp 1667941163
transform 1 0 17756 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_185
timestamp 1667941163
transform 1 0 18124 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_206
timestamp 1667941163
transform 1 0 20056 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_49_216
timestamp 1667941163
transform 1 0 20976 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_49_225
timestamp 1667941163
transform 1 0 21804 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_235
timestamp 1667941163
transform 1 0 22724 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_242
timestamp 1667941163
transform 1 0 23368 0 -1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_49_249
timestamp 1667941163
transform 1 0 24012 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_261
timestamp 1667941163
transform 1 0 25116 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_49_271
timestamp 1667941163
transform 1 0 26036 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_279
timestamp 1667941163
transform 1 0 26772 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_49_281
timestamp 1667941163
transform 1 0 26956 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_49_287
timestamp 1667941163
transform 1 0 27508 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_294
timestamp 1667941163
transform 1 0 28152 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_298
timestamp 1667941163
transform 1 0 28520 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_3
timestamp 1667941163
transform 1 0 1380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_15
timestamp 1667941163
transform 1 0 2484 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_27
timestamp 1667941163
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_29
timestamp 1667941163
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_41
timestamp 1667941163
transform 1 0 4876 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_53
timestamp 1667941163
transform 1 0 5980 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_65
timestamp 1667941163
transform 1 0 7084 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_77
timestamp 1667941163
transform 1 0 8188 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_83
timestamp 1667941163
transform 1 0 8740 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_85
timestamp 1667941163
transform 1 0 8924 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_97
timestamp 1667941163
transform 1 0 10028 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_109
timestamp 1667941163
transform 1 0 11132 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_121
timestamp 1667941163
transform 1 0 12236 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_133
timestamp 1667941163
transform 1 0 13340 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_139
timestamp 1667941163
transform 1 0 13892 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_141
timestamp 1667941163
transform 1 0 14076 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_153
timestamp 1667941163
transform 1 0 15180 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_165
timestamp 1667941163
transform 1 0 16284 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_172
timestamp 1667941163
transform 1 0 16928 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_192
timestamp 1667941163
transform 1 0 18768 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_50_197
timestamp 1667941163
transform 1 0 19228 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_215
timestamp 1667941163
transform 1 0 20884 0 1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_50_235
timestamp 1667941163
transform 1 0 22724 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_247
timestamp 1667941163
transform 1 0 23828 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_251
timestamp 1667941163
transform 1 0 24196 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_50_253
timestamp 1667941163
transform 1 0 24380 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_262
timestamp 1667941163
transform 1 0 25208 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_266
timestamp 1667941163
transform 1 0 25576 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_272
timestamp 1667941163
transform 1 0 26128 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_50_297
timestamp 1667941163
transform 1 0 28428 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_3
timestamp 1667941163
transform 1 0 1380 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_51_15
timestamp 1667941163
transform 1 0 2484 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_27
timestamp 1667941163
transform 1 0 3588 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_39
timestamp 1667941163
transform 1 0 4692 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_51
timestamp 1667941163
transform 1 0 5796 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_55
timestamp 1667941163
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_57
timestamp 1667941163
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_69
timestamp 1667941163
transform 1 0 7452 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_81
timestamp 1667941163
transform 1 0 8556 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_93
timestamp 1667941163
transform 1 0 9660 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_105
timestamp 1667941163
transform 1 0 10764 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_111
timestamp 1667941163
transform 1 0 11316 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_113
timestamp 1667941163
transform 1 0 11500 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_125
timestamp 1667941163
transform 1 0 12604 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_137
timestamp 1667941163
transform 1 0 13708 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_149
timestamp 1667941163
transform 1 0 14812 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_51_161
timestamp 1667941163
transform 1 0 15916 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_166
timestamp 1667941163
transform 1 0 16376 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_169
timestamp 1667941163
transform 1 0 16652 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_51_179
timestamp 1667941163
transform 1 0 17572 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_191
timestamp 1667941163
transform 1 0 18676 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_199
timestamp 1667941163
transform 1 0 19412 0 -1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_51_209
timestamp 1667941163
transform 1 0 20332 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_51_221
timestamp 1667941163
transform 1 0 21436 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_51_225
timestamp 1667941163
transform 1 0 21804 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_51_231
timestamp 1667941163
transform 1 0 22356 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_51_239
timestamp 1667941163
transform 1 0 23092 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_246
timestamp 1667941163
transform 1 0 23736 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_250
timestamp 1667941163
transform 1 0 24104 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_255
timestamp 1667941163
transform 1 0 24564 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_267
timestamp 1667941163
transform 1 0 25668 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_51_277
timestamp 1667941163
transform 1 0 26588 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_51_281
timestamp 1667941163
transform 1 0 26956 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_51_286
timestamp 1667941163
transform 1 0 27416 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_51_297
timestamp 1667941163
transform 1 0 28428 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_52_3
timestamp 1667941163
transform 1 0 1380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_15
timestamp 1667941163
transform 1 0 2484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_27
timestamp 1667941163
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_29
timestamp 1667941163
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_41
timestamp 1667941163
transform 1 0 4876 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_53
timestamp 1667941163
transform 1 0 5980 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_65
timestamp 1667941163
transform 1 0 7084 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_77
timestamp 1667941163
transform 1 0 8188 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_83
timestamp 1667941163
transform 1 0 8740 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_85
timestamp 1667941163
transform 1 0 8924 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_97
timestamp 1667941163
transform 1 0 10028 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_109
timestamp 1667941163
transform 1 0 11132 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_121
timestamp 1667941163
transform 1 0 12236 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_133
timestamp 1667941163
transform 1 0 13340 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_139
timestamp 1667941163
transform 1 0 13892 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_141
timestamp 1667941163
transform 1 0 14076 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_153
timestamp 1667941163
transform 1 0 15180 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_52_164
timestamp 1667941163
transform 1 0 16192 0 1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_52_173
timestamp 1667941163
transform 1 0 17020 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_185
timestamp 1667941163
transform 1 0 18124 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_192
timestamp 1667941163
transform 1 0 18768 0 1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_52_197
timestamp 1667941163
transform 1 0 19228 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_209
timestamp 1667941163
transform 1 0 20332 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_221
timestamp 1667941163
transform 1 0 21436 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_52_229
timestamp 1667941163
transform 1 0 22172 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_52_235
timestamp 1667941163
transform 1 0 22724 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_247
timestamp 1667941163
transform 1 0 23828 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_251
timestamp 1667941163
transform 1 0 24196 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_52_253
timestamp 1667941163
transform 1 0 24380 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_260
timestamp 1667941163
transform 1 0 25024 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_52_269
timestamp 1667941163
transform 1 0 25852 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_52_296
timestamp 1667941163
transform 1 0 28336 0 1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_53_3
timestamp 1667941163
transform 1 0 1380 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_15
timestamp 1667941163
transform 1 0 2484 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_27
timestamp 1667941163
transform 1 0 3588 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_39
timestamp 1667941163
transform 1 0 4692 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_51
timestamp 1667941163
transform 1 0 5796 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_55
timestamp 1667941163
transform 1 0 6164 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_57
timestamp 1667941163
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_69
timestamp 1667941163
transform 1 0 7452 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_81
timestamp 1667941163
transform 1 0 8556 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_93
timestamp 1667941163
transform 1 0 9660 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_105
timestamp 1667941163
transform 1 0 10764 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_111
timestamp 1667941163
transform 1 0 11316 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_113
timestamp 1667941163
transform 1 0 11500 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_125
timestamp 1667941163
transform 1 0 12604 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_137
timestamp 1667941163
transform 1 0 13708 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_149
timestamp 1667941163
transform 1 0 14812 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_53_166
timestamp 1667941163
transform 1 0 16376 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_169
timestamp 1667941163
transform 1 0 16652 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_174
timestamp 1667941163
transform 1 0 17112 0 -1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_53_194
timestamp 1667941163
transform 1 0 18952 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_53_206
timestamp 1667941163
transform 1 0 20056 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_210
timestamp 1667941163
transform 1 0 20424 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_53_222
timestamp 1667941163
transform 1 0 21528 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_225
timestamp 1667941163
transform 1 0 21804 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_230
timestamp 1667941163
transform 1 0 22264 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_53_241
timestamp 1667941163
transform 1 0 23276 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_53_252
timestamp 1667941163
transform 1 0 24288 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_256
timestamp 1667941163
transform 1 0 24656 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_53_278
timestamp 1667941163
transform 1 0 26680 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_53_281
timestamp 1667941163
transform 1 0 26956 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_53_292
timestamp 1667941163
transform 1 0 27968 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_298
timestamp 1667941163
transform 1 0 28520 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_3
timestamp 1667941163
transform 1 0 1380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_15
timestamp 1667941163
transform 1 0 2484 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_27
timestamp 1667941163
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_29
timestamp 1667941163
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_41
timestamp 1667941163
transform 1 0 4876 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_53
timestamp 1667941163
transform 1 0 5980 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_65
timestamp 1667941163
transform 1 0 7084 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_77
timestamp 1667941163
transform 1 0 8188 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_83
timestamp 1667941163
transform 1 0 8740 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_85
timestamp 1667941163
transform 1 0 8924 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_97
timestamp 1667941163
transform 1 0 10028 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_109
timestamp 1667941163
transform 1 0 11132 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_121
timestamp 1667941163
transform 1 0 12236 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_54_130
timestamp 1667941163
transform 1 0 13064 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_54_138
timestamp 1667941163
transform 1 0 13800 0 1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_54_141
timestamp 1667941163
transform 1 0 14076 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_153
timestamp 1667941163
transform 1 0 15180 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_54_173
timestamp 1667941163
transform 1 0 17020 0 1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_54_180
timestamp 1667941163
transform 1 0 17664 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_54_192
timestamp 1667941163
transform 1 0 18768 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_54_197
timestamp 1667941163
transform 1 0 19228 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_207
timestamp 1667941163
transform 1 0 20148 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_214
timestamp 1667941163
transform 1 0 20792 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_234
timestamp 1667941163
transform 1 0 22632 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_54_246
timestamp 1667941163
transform 1 0 23736 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_54_253
timestamp 1667941163
transform 1 0 24380 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_54_261
timestamp 1667941163
transform 1 0 25116 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_267
timestamp 1667941163
transform 1 0 25668 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_289
timestamp 1667941163
transform 1 0 27692 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_54_296
timestamp 1667941163
transform 1 0 28336 0 1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_55_3
timestamp 1667941163
transform 1 0 1380 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_15
timestamp 1667941163
transform 1 0 2484 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_27
timestamp 1667941163
transform 1 0 3588 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_39
timestamp 1667941163
transform 1 0 4692 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_51
timestamp 1667941163
transform 1 0 5796 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_55
timestamp 1667941163
transform 1 0 6164 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_57
timestamp 1667941163
transform 1 0 6348 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_69
timestamp 1667941163
transform 1 0 7452 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_81
timestamp 1667941163
transform 1 0 8556 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_93
timestamp 1667941163
transform 1 0 9660 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_105
timestamp 1667941163
transform 1 0 10764 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_111
timestamp 1667941163
transform 1 0 11316 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_113
timestamp 1667941163
transform 1 0 11500 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_55_125
timestamp 1667941163
transform 1 0 12604 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_147
timestamp 1667941163
transform 1 0 14628 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_159
timestamp 1667941163
transform 1 0 15732 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_55_167
timestamp 1667941163
transform 1 0 16468 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_169
timestamp 1667941163
transform 1 0 16652 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_181
timestamp 1667941163
transform 1 0 17756 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_55_189
timestamp 1667941163
transform 1 0 18492 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_194
timestamp 1667941163
transform 1 0 18952 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_214
timestamp 1667941163
transform 1 0 20792 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_55_221
timestamp 1667941163
transform 1 0 21436 0 -1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_55_225
timestamp 1667941163
transform 1 0 21804 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_55_237
timestamp 1667941163
transform 1 0 22908 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_55_243
timestamp 1667941163
transform 1 0 23460 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_255
timestamp 1667941163
transform 1 0 24564 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_55_267
timestamp 1667941163
transform 1 0 25668 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_55_272
timestamp 1667941163
transform 1 0 26128 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_55_281
timestamp 1667941163
transform 1 0 26956 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_55_287
timestamp 1667941163
transform 1 0 27508 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_294
timestamp 1667941163
transform 1 0 28152 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_298
timestamp 1667941163
transform 1 0 28520 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_3
timestamp 1667941163
transform 1 0 1380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_15
timestamp 1667941163
transform 1 0 2484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_27
timestamp 1667941163
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_29
timestamp 1667941163
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_41
timestamp 1667941163
transform 1 0 4876 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_53
timestamp 1667941163
transform 1 0 5980 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_65
timestamp 1667941163
transform 1 0 7084 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_77
timestamp 1667941163
transform 1 0 8188 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_83
timestamp 1667941163
transform 1 0 8740 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_85
timestamp 1667941163
transform 1 0 8924 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_97
timestamp 1667941163
transform 1 0 10028 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_109
timestamp 1667941163
transform 1 0 11132 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_121
timestamp 1667941163
transform 1 0 12236 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_133
timestamp 1667941163
transform 1 0 13340 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_139
timestamp 1667941163
transform 1 0 13892 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_141
timestamp 1667941163
transform 1 0 14076 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_153
timestamp 1667941163
transform 1 0 15180 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_56_161
timestamp 1667941163
transform 1 0 15916 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_168
timestamp 1667941163
transform 1 0 16560 0 1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_56_175
timestamp 1667941163
transform 1 0 17204 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_187
timestamp 1667941163
transform 1 0 18308 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_56_195
timestamp 1667941163
transform 1 0 19044 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_56_197
timestamp 1667941163
transform 1 0 19228 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_203
timestamp 1667941163
transform 1 0 19780 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_212
timestamp 1667941163
transform 1 0 20608 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_224
timestamp 1667941163
transform 1 0 21712 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_236
timestamp 1667941163
transform 1 0 22816 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_56_250
timestamp 1667941163
transform 1 0 24104 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_56_253
timestamp 1667941163
transform 1 0 24380 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_56_261
timestamp 1667941163
transform 1 0 25116 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_265
timestamp 1667941163
transform 1 0 25484 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_56_270
timestamp 1667941163
transform 1 0 25944 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_56_297
timestamp 1667941163
transform 1 0 28428 0 1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_57_3
timestamp 1667941163
transform 1 0 1380 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_15
timestamp 1667941163
transform 1 0 2484 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_27
timestamp 1667941163
transform 1 0 3588 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_39
timestamp 1667941163
transform 1 0 4692 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_51
timestamp 1667941163
transform 1 0 5796 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_55
timestamp 1667941163
transform 1 0 6164 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_57
timestamp 1667941163
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_69
timestamp 1667941163
transform 1 0 7452 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_81
timestamp 1667941163
transform 1 0 8556 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_93
timestamp 1667941163
transform 1 0 9660 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_105
timestamp 1667941163
transform 1 0 10764 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_111
timestamp 1667941163
transform 1 0 11316 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_113
timestamp 1667941163
transform 1 0 11500 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_125
timestamp 1667941163
transform 1 0 12604 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_137
timestamp 1667941163
transform 1 0 13708 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_149
timestamp 1667941163
transform 1 0 14812 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_57_157
timestamp 1667941163
transform 1 0 15548 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_166
timestamp 1667941163
transform 1 0 16376 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_169
timestamp 1667941163
transform 1 0 16652 0 -1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_57_189
timestamp 1667941163
transform 1 0 18492 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_201
timestamp 1667941163
transform 1 0 19596 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_213
timestamp 1667941163
transform 1 0 20700 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_217
timestamp 1667941163
transform 1 0 21068 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_57_221
timestamp 1667941163
transform 1 0 21436 0 -1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_57_225
timestamp 1667941163
transform 1 0 21804 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_237
timestamp 1667941163
transform 1 0 22908 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_243
timestamp 1667941163
transform 1 0 23460 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_57_260
timestamp 1667941163
transform 1 0 25024 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_57_268
timestamp 1667941163
transform 1 0 25760 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_57_278
timestamp 1667941163
transform 1 0 26680 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_281
timestamp 1667941163
transform 1 0 26956 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_288
timestamp 1667941163
transform 1 0 27600 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_295
timestamp 1667941163
transform 1 0 28244 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_58_3
timestamp 1667941163
transform 1 0 1380 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_9
timestamp 1667941163
transform 1 0 1932 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_13
timestamp 1667941163
transform 1 0 2300 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_58_25
timestamp 1667941163
transform 1 0 3404 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_58_29
timestamp 1667941163
transform 1 0 3772 0 1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_58_43
timestamp 1667941163
transform 1 0 5060 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_55
timestamp 1667941163
transform 1 0 6164 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_67
timestamp 1667941163
transform 1 0 7268 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_58_79
timestamp 1667941163
transform 1 0 8372 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_83
timestamp 1667941163
transform 1 0 8740 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_85
timestamp 1667941163
transform 1 0 8924 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_97
timestamp 1667941163
transform 1 0 10028 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_109
timestamp 1667941163
transform 1 0 11132 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_121
timestamp 1667941163
transform 1 0 12236 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_133
timestamp 1667941163
transform 1 0 13340 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_139
timestamp 1667941163
transform 1 0 13892 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_141
timestamp 1667941163
transform 1 0 14076 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_153
timestamp 1667941163
transform 1 0 15180 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_58_161
timestamp 1667941163
transform 1 0 15916 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_165
timestamp 1667941163
transform 1 0 16284 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_177
timestamp 1667941163
transform 1 0 17388 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_189
timestamp 1667941163
transform 1 0 18492 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_195
timestamp 1667941163
transform 1 0 19044 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_197
timestamp 1667941163
transform 1 0 19228 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_209
timestamp 1667941163
transform 1 0 20332 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_58_213
timestamp 1667941163
transform 1 0 20700 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_58_236
timestamp 1667941163
transform 1 0 22816 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_242
timestamp 1667941163
transform 1 0 23368 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_58_250
timestamp 1667941163
transform 1 0 24104 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_58_253
timestamp 1667941163
transform 1 0 24380 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_58_272
timestamp 1667941163
transform 1 0 26128 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_58_297
timestamp 1667941163
transform 1 0 28428 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_59_3
timestamp 1667941163
transform 1 0 1380 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_59_27
timestamp 1667941163
transform 1 0 3588 0 -1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_59_43
timestamp 1667941163
transform 1 0 5060 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_59_55
timestamp 1667941163
transform 1 0 6164 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_57
timestamp 1667941163
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_69
timestamp 1667941163
transform 1 0 7452 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_81
timestamp 1667941163
transform 1 0 8556 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_93
timestamp 1667941163
transform 1 0 9660 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_105
timestamp 1667941163
transform 1 0 10764 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_111
timestamp 1667941163
transform 1 0 11316 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_113
timestamp 1667941163
transform 1 0 11500 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_125
timestamp 1667941163
transform 1 0 12604 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_137
timestamp 1667941163
transform 1 0 13708 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_149
timestamp 1667941163
transform 1 0 14812 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_155
timestamp 1667941163
transform 1 0 15364 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_59_161
timestamp 1667941163
transform 1 0 15916 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_167
timestamp 1667941163
transform 1 0 16468 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_169
timestamp 1667941163
transform 1 0 16652 0 -1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_59_189
timestamp 1667941163
transform 1 0 18492 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_201
timestamp 1667941163
transform 1 0 19596 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_59_214
timestamp 1667941163
transform 1 0 20792 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_59_222
timestamp 1667941163
transform 1 0 21528 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_59_225
timestamp 1667941163
transform 1 0 21804 0 -1 34816
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_59_249
timestamp 1667941163
transform 1 0 24012 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_59_261
timestamp 1667941163
transform 1 0 25116 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_59_278
timestamp 1667941163
transform 1 0 26680 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_281
timestamp 1667941163
transform 1 0 26956 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_59_291
timestamp 1667941163
transform 1 0 27876 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_60_3
timestamp 1667941163
transform 1 0 1380 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_60_9
timestamp 1667941163
transform 1 0 1932 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_13
timestamp 1667941163
transform 1 0 2300 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_60_26
timestamp 1667941163
transform 1 0 3496 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_60_29
timestamp 1667941163
transform 1 0 3772 0 1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_60_43
timestamp 1667941163
transform 1 0 5060 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_55
timestamp 1667941163
transform 1 0 6164 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_67
timestamp 1667941163
transform 1 0 7268 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_60_79
timestamp 1667941163
transform 1 0 8372 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_83
timestamp 1667941163
transform 1 0 8740 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_85
timestamp 1667941163
transform 1 0 8924 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_97
timestamp 1667941163
transform 1 0 10028 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_109
timestamp 1667941163
transform 1 0 11132 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_121
timestamp 1667941163
transform 1 0 12236 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_133
timestamp 1667941163
transform 1 0 13340 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_139
timestamp 1667941163
transform 1 0 13892 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_141
timestamp 1667941163
transform 1 0 14076 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_153
timestamp 1667941163
transform 1 0 15180 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_165
timestamp 1667941163
transform 1 0 16284 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_60_187
timestamp 1667941163
transform 1 0 18308 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_60_195
timestamp 1667941163
transform 1 0 19044 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_60_197
timestamp 1667941163
transform 1 0 19228 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_60_215
timestamp 1667941163
transform 1 0 20884 0 1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_60_235
timestamp 1667941163
transform 1 0 22724 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_60_247
timestamp 1667941163
transform 1 0 23828 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_251
timestamp 1667941163
transform 1 0 24196 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_60_253
timestamp 1667941163
transform 1 0 24380 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_259
timestamp 1667941163
transform 1 0 24932 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_276
timestamp 1667941163
transform 1 0 26496 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_60_296
timestamp 1667941163
transform 1 0 28336 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_61_3
timestamp 1667941163
transform 1 0 1380 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_61_23
timestamp 1667941163
transform 1 0 3220 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_39
timestamp 1667941163
transform 1 0 4692 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_52
timestamp 1667941163
transform 1 0 5888 0 -1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_61_57
timestamp 1667941163
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_69
timestamp 1667941163
transform 1 0 7452 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_81
timestamp 1667941163
transform 1 0 8556 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_93
timestamp 1667941163
transform 1 0 9660 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_105
timestamp 1667941163
transform 1 0 10764 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_111
timestamp 1667941163
transform 1 0 11316 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_113
timestamp 1667941163
transform 1 0 11500 0 -1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_61_129
timestamp 1667941163
transform 1 0 12972 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_141
timestamp 1667941163
transform 1 0 14076 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_153
timestamp 1667941163
transform 1 0 15180 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_61_162
timestamp 1667941163
transform 1 0 16008 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_61_169
timestamp 1667941163
transform 1 0 16652 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_61_174
timestamp 1667941163
transform 1 0 17112 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_61_182
timestamp 1667941163
transform 1 0 17848 0 -1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_61_201
timestamp 1667941163
transform 1 0 19596 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_213
timestamp 1667941163
transform 1 0 20700 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_61_221
timestamp 1667941163
transform 1 0 21436 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_61_225
timestamp 1667941163
transform 1 0 21804 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_61_233
timestamp 1667941163
transform 1 0 22540 0 -1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_61_239
timestamp 1667941163
transform 1 0 23092 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_251
timestamp 1667941163
transform 1 0 24196 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_61_259
timestamp 1667941163
transform 1 0 24932 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_61_269
timestamp 1667941163
transform 1 0 25852 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_276
timestamp 1667941163
transform 1 0 26496 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_61_281
timestamp 1667941163
transform 1 0 26956 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_61_286
timestamp 1667941163
transform 1 0 27416 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_61_293
timestamp 1667941163
transform 1 0 28060 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_62_3
timestamp 1667941163
transform 1 0 1380 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_62_26
timestamp 1667941163
transform 1 0 3496 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_62_29
timestamp 1667941163
transform 1 0 3772 0 1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_62_44
timestamp 1667941163
transform 1 0 5152 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_56
timestamp 1667941163
transform 1 0 6256 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_68
timestamp 1667941163
transform 1 0 7360 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_62_80
timestamp 1667941163
transform 1 0 8464 0 1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_62_85
timestamp 1667941163
transform 1 0 8924 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_97
timestamp 1667941163
transform 1 0 10028 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_109
timestamp 1667941163
transform 1 0 11132 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_121
timestamp 1667941163
transform 1 0 12236 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_133
timestamp 1667941163
transform 1 0 13340 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_139
timestamp 1667941163
transform 1 0 13892 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_141
timestamp 1667941163
transform 1 0 14076 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_153
timestamp 1667941163
transform 1 0 15180 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_165
timestamp 1667941163
transform 1 0 16284 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_171
timestamp 1667941163
transform 1 0 16836 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_175
timestamp 1667941163
transform 1 0 17204 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_187
timestamp 1667941163
transform 1 0 18308 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_62_195
timestamp 1667941163
transform 1 0 19044 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_62_197
timestamp 1667941163
transform 1 0 19228 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_62_210
timestamp 1667941163
transform 1 0 20424 0 1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_62_217
timestamp 1667941163
transform 1 0 21068 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_229
timestamp 1667941163
transform 1 0 22172 0 1 35904
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_62_240
timestamp 1667941163
transform 1 0 23184 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_253
timestamp 1667941163
transform 1 0 24380 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_265
timestamp 1667941163
transform 1 0 25484 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_62_273
timestamp 1667941163
transform 1 0 26220 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_62_297
timestamp 1667941163
transform 1 0 28428 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_63_3
timestamp 1667941163
transform 1 0 1380 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_63_9
timestamp 1667941163
transform 1 0 1932 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_24
timestamp 1667941163
transform 1 0 3312 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_40
timestamp 1667941163
transform 1 0 4784 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_63_47
timestamp 1667941163
transform 1 0 5428 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_55
timestamp 1667941163
transform 1 0 6164 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_57
timestamp 1667941163
transform 1 0 6348 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_69
timestamp 1667941163
transform 1 0 7452 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_81
timestamp 1667941163
transform 1 0 8556 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_93
timestamp 1667941163
transform 1 0 9660 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_105
timestamp 1667941163
transform 1 0 10764 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_111
timestamp 1667941163
transform 1 0 11316 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_113
timestamp 1667941163
transform 1 0 11500 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_125
timestamp 1667941163
transform 1 0 12604 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_137
timestamp 1667941163
transform 1 0 13708 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_149
timestamp 1667941163
transform 1 0 14812 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_63_166
timestamp 1667941163
transform 1 0 16376 0 -1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_63_169
timestamp 1667941163
transform 1 0 16652 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_181
timestamp 1667941163
transform 1 0 17756 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_63_193
timestamp 1667941163
transform 1 0 18860 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_63_198
timestamp 1667941163
transform 1 0 19320 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_206
timestamp 1667941163
transform 1 0 20056 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_215
timestamp 1667941163
transform 1 0 20884 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_63_222
timestamp 1667941163
transform 1 0 21528 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_63_225
timestamp 1667941163
transform 1 0 21804 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_229
timestamp 1667941163
transform 1 0 22172 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_236
timestamp 1667941163
transform 1 0 22816 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_248
timestamp 1667941163
transform 1 0 23920 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_260
timestamp 1667941163
transform 1 0 25024 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_268
timestamp 1667941163
transform 1 0 25760 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_272
timestamp 1667941163
transform 1 0 26128 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_63_281
timestamp 1667941163
transform 1 0 26956 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_63_286
timestamp 1667941163
transform 1 0 27416 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_290
timestamp 1667941163
transform 1 0 27784 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_294
timestamp 1667941163
transform 1 0 28152 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_298
timestamp 1667941163
transform 1 0 28520 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_3
timestamp 1667941163
transform 1 0 1380 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_26
timestamp 1667941163
transform 1 0 3496 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_29
timestamp 1667941163
transform 1 0 3772 0 1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_64_52
timestamp 1667941163
transform 1 0 5888 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_64
timestamp 1667941163
transform 1 0 6992 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_76
timestamp 1667941163
transform 1 0 8096 0 1 36992
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_64_85
timestamp 1667941163
transform 1 0 8924 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_97
timestamp 1667941163
transform 1 0 10028 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_109
timestamp 1667941163
transform 1 0 11132 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_121
timestamp 1667941163
transform 1 0 12236 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_133
timestamp 1667941163
transform 1 0 13340 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_139
timestamp 1667941163
transform 1 0 13892 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_141
timestamp 1667941163
transform 1 0 14076 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_64_153
timestamp 1667941163
transform 1 0 15180 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_163
timestamp 1667941163
transform 1 0 16100 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_171
timestamp 1667941163
transform 1 0 16836 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_177
timestamp 1667941163
transform 1 0 17388 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_64_188
timestamp 1667941163
transform 1 0 18400 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_197
timestamp 1667941163
transform 1 0 19228 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_202
timestamp 1667941163
transform 1 0 19688 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_213
timestamp 1667941163
transform 1 0 20700 0 1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_64_220
timestamp 1667941163
transform 1 0 21344 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_232
timestamp 1667941163
transform 1 0 22448 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_236
timestamp 1667941163
transform 1 0 22816 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_64_246
timestamp 1667941163
transform 1 0 23736 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_64_253
timestamp 1667941163
transform 1 0 24380 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_258
timestamp 1667941163
transform 1 0 24840 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_64_266
timestamp 1667941163
transform 1 0 25576 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_64_290
timestamp 1667941163
transform 1 0 27784 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_64_297
timestamp 1667941163
transform 1 0 28428 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_65_3
timestamp 1667941163
transform 1 0 1380 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_65_32
timestamp 1667941163
transform 1 0 4048 0 -1 38080
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_65_39
timestamp 1667941163
transform 1 0 4692 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_51
timestamp 1667941163
transform 1 0 5796 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_55
timestamp 1667941163
transform 1 0 6164 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_57
timestamp 1667941163
transform 1 0 6348 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_69
timestamp 1667941163
transform 1 0 7452 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_81
timestamp 1667941163
transform 1 0 8556 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_93
timestamp 1667941163
transform 1 0 9660 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_105
timestamp 1667941163
transform 1 0 10764 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_111
timestamp 1667941163
transform 1 0 11316 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_113
timestamp 1667941163
transform 1 0 11500 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_125
timestamp 1667941163
transform 1 0 12604 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_137
timestamp 1667941163
transform 1 0 13708 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_149
timestamp 1667941163
transform 1 0 14812 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_65_161
timestamp 1667941163
transform 1 0 15916 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_65_166
timestamp 1667941163
transform 1 0 16376 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_65_169
timestamp 1667941163
transform 1 0 16652 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_65_179
timestamp 1667941163
transform 1 0 17572 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_183
timestamp 1667941163
transform 1 0 17940 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_65_193
timestamp 1667941163
transform 1 0 18860 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_199
timestamp 1667941163
transform 1 0 19412 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_204
timestamp 1667941163
transform 1 0 19872 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_65_216
timestamp 1667941163
transform 1 0 20976 0 -1 38080
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_65_225
timestamp 1667941163
transform 1 0 21804 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_237
timestamp 1667941163
transform 1 0 22908 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_249
timestamp 1667941163
transform 1 0 24012 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_261
timestamp 1667941163
transform 1 0 25116 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_273
timestamp 1667941163
transform 1 0 26220 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_279
timestamp 1667941163
transform 1 0 26772 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_65_281
timestamp 1667941163
transform 1 0 26956 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_65_286
timestamp 1667941163
transform 1 0 27416 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_65_293
timestamp 1667941163
transform 1 0 28060 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_66_3
timestamp 1667941163
transform 1 0 1380 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_66_9
timestamp 1667941163
transform 1 0 1932 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_66_17
timestamp 1667941163
transform 1 0 2668 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_66_21
timestamp 1667941163
transform 1 0 3036 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_27
timestamp 1667941163
transform 1 0 3588 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_29
timestamp 1667941163
transform 1 0 3772 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_41
timestamp 1667941163
transform 1 0 4876 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_53
timestamp 1667941163
transform 1 0 5980 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_65
timestamp 1667941163
transform 1 0 7084 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_77
timestamp 1667941163
transform 1 0 8188 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_83
timestamp 1667941163
transform 1 0 8740 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_85
timestamp 1667941163
transform 1 0 8924 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_97
timestamp 1667941163
transform 1 0 10028 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_109
timestamp 1667941163
transform 1 0 11132 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_121
timestamp 1667941163
transform 1 0 12236 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_133
timestamp 1667941163
transform 1 0 13340 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_139
timestamp 1667941163
transform 1 0 13892 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_66_141
timestamp 1667941163
transform 1 0 14076 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_66_149
timestamp 1667941163
transform 1 0 14812 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_66_157
timestamp 1667941163
transform 1 0 15548 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_66_168
timestamp 1667941163
transform 1 0 16560 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_174
timestamp 1667941163
transform 1 0 17112 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_66_182
timestamp 1667941163
transform 1 0 17848 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_66_189
timestamp 1667941163
transform 1 0 18492 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_195
timestamp 1667941163
transform 1 0 19044 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_197
timestamp 1667941163
transform 1 0 19228 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_66_209
timestamp 1667941163
transform 1 0 20332 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_66_217
timestamp 1667941163
transform 1 0 21068 0 1 38080
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_66_222
timestamp 1667941163
transform 1 0 21528 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_234
timestamp 1667941163
transform 1 0 22632 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_246
timestamp 1667941163
transform 1 0 23736 0 1 38080
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_66_253
timestamp 1667941163
transform 1 0 24380 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_66_265
timestamp 1667941163
transform 1 0 25484 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_66_273
timestamp 1667941163
transform 1 0 26220 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_66_297
timestamp 1667941163
transform 1 0 28428 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_67_3
timestamp 1667941163
transform 1 0 1380 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_67_12
timestamp 1667941163
transform 1 0 2208 0 -1 39168
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_67_19
timestamp 1667941163
transform 1 0 2852 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_31
timestamp 1667941163
transform 1 0 3956 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_43
timestamp 1667941163
transform 1 0 5060 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_67_55
timestamp 1667941163
transform 1 0 6164 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_57
timestamp 1667941163
transform 1 0 6348 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_69
timestamp 1667941163
transform 1 0 7452 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_81
timestamp 1667941163
transform 1 0 8556 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_93
timestamp 1667941163
transform 1 0 9660 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_105
timestamp 1667941163
transform 1 0 10764 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_111
timestamp 1667941163
transform 1 0 11316 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_113
timestamp 1667941163
transform 1 0 11500 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_125
timestamp 1667941163
transform 1 0 12604 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_137
timestamp 1667941163
transform 1 0 13708 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_149
timestamp 1667941163
transform 1 0 14812 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_161
timestamp 1667941163
transform 1 0 15916 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_167
timestamp 1667941163
transform 1 0 16468 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_169
timestamp 1667941163
transform 1 0 16652 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_181
timestamp 1667941163
transform 1 0 17756 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_185
timestamp 1667941163
transform 1 0 18124 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_67_189
timestamp 1667941163
transform 1 0 18492 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_67_200
timestamp 1667941163
transform 1 0 19504 0 -1 39168
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_67_207
timestamp 1667941163
transform 1 0 20148 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_219
timestamp 1667941163
transform 1 0 21252 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_223
timestamp 1667941163
transform 1 0 21620 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_67_225
timestamp 1667941163
transform 1 0 21804 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_67_248
timestamp 1667941163
transform 1 0 23920 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_67_256
timestamp 1667941163
transform 1 0 24656 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_67_278
timestamp 1667941163
transform 1 0 26680 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_67_281
timestamp 1667941163
transform 1 0 26956 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_67_292
timestamp 1667941163
transform 1 0 27968 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_298
timestamp 1667941163
transform 1 0 28520 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_68_3
timestamp 1667941163
transform 1 0 1380 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_68_8
timestamp 1667941163
transform 1 0 1840 0 1 39168
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_68_15
timestamp 1667941163
transform 1 0 2484 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_68_27
timestamp 1667941163
transform 1 0 3588 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_29
timestamp 1667941163
transform 1 0 3772 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_41
timestamp 1667941163
transform 1 0 4876 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_53
timestamp 1667941163
transform 1 0 5980 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_65
timestamp 1667941163
transform 1 0 7084 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_77
timestamp 1667941163
transform 1 0 8188 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_83
timestamp 1667941163
transform 1 0 8740 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_85
timestamp 1667941163
transform 1 0 8924 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_97
timestamp 1667941163
transform 1 0 10028 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_109
timestamp 1667941163
transform 1 0 11132 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_121
timestamp 1667941163
transform 1 0 12236 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_133
timestamp 1667941163
transform 1 0 13340 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_139
timestamp 1667941163
transform 1 0 13892 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_141
timestamp 1667941163
transform 1 0 14076 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_153
timestamp 1667941163
transform 1 0 15180 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_165
timestamp 1667941163
transform 1 0 16284 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_68_177
timestamp 1667941163
transform 1 0 17388 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_68_182
timestamp 1667941163
transform 1 0 17848 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_68_194
timestamp 1667941163
transform 1 0 18952 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_68_197
timestamp 1667941163
transform 1 0 19228 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_68_208
timestamp 1667941163
transform 1 0 20240 0 1 39168
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_68_215
timestamp 1667941163
transform 1 0 20884 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_227
timestamp 1667941163
transform 1 0 21988 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_239
timestamp 1667941163
transform 1 0 23092 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_68_251
timestamp 1667941163
transform 1 0 24196 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_253
timestamp 1667941163
transform 1 0 24380 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_68_265
timestamp 1667941163
transform 1 0 25484 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_68_273
timestamp 1667941163
transform 1 0 26220 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_68_297
timestamp 1667941163
transform 1 0 28428 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_69_3
timestamp 1667941163
transform 1 0 1380 0 -1 40256
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_69_27
timestamp 1667941163
transform 1 0 3588 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_39
timestamp 1667941163
transform 1 0 4692 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_69_51
timestamp 1667941163
transform 1 0 5796 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_55
timestamp 1667941163
transform 1 0 6164 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_57
timestamp 1667941163
transform 1 0 6348 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_69
timestamp 1667941163
transform 1 0 7452 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_81
timestamp 1667941163
transform 1 0 8556 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_93
timestamp 1667941163
transform 1 0 9660 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_105
timestamp 1667941163
transform 1 0 10764 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_111
timestamp 1667941163
transform 1 0 11316 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_113
timestamp 1667941163
transform 1 0 11500 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_125
timestamp 1667941163
transform 1 0 12604 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_137
timestamp 1667941163
transform 1 0 13708 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_149
timestamp 1667941163
transform 1 0 14812 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_161
timestamp 1667941163
transform 1 0 15916 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_167
timestamp 1667941163
transform 1 0 16468 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_69_169
timestamp 1667941163
transform 1 0 16652 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_181
timestamp 1667941163
transform 1 0 17756 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_69_190
timestamp 1667941163
transform 1 0 18584 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_69_198
timestamp 1667941163
transform 1 0 19320 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_204
timestamp 1667941163
transform 1 0 19872 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_69_216
timestamp 1667941163
transform 1 0 20976 0 -1 40256
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_69_225
timestamp 1667941163
transform 1 0 21804 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_237
timestamp 1667941163
transform 1 0 22908 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_249
timestamp 1667941163
transform 1 0 24012 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_261
timestamp 1667941163
transform 1 0 25116 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_273
timestamp 1667941163
transform 1 0 26220 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_279
timestamp 1667941163
transform 1 0 26772 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_69_281
timestamp 1667941163
transform 1 0 26956 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_288
timestamp 1667941163
transform 1 0 27600 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_295
timestamp 1667941163
transform 1 0 28244 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_3
timestamp 1667941163
transform 1 0 1380 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_10
timestamp 1667941163
transform 1 0 2024 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_70_17
timestamp 1667941163
transform 1 0 2668 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_70_25
timestamp 1667941163
transform 1 0 3404 0 1 40256
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_70_29
timestamp 1667941163
transform 1 0 3772 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_41
timestamp 1667941163
transform 1 0 4876 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_53
timestamp 1667941163
transform 1 0 5980 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_65
timestamp 1667941163
transform 1 0 7084 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_77
timestamp 1667941163
transform 1 0 8188 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_83
timestamp 1667941163
transform 1 0 8740 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_85
timestamp 1667941163
transform 1 0 8924 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_97
timestamp 1667941163
transform 1 0 10028 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_109
timestamp 1667941163
transform 1 0 11132 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_121
timestamp 1667941163
transform 1 0 12236 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_133
timestamp 1667941163
transform 1 0 13340 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_139
timestamp 1667941163
transform 1 0 13892 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_141
timestamp 1667941163
transform 1 0 14076 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_153
timestamp 1667941163
transform 1 0 15180 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_165
timestamp 1667941163
transform 1 0 16284 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_70_177
timestamp 1667941163
transform 1 0 17388 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_70_182
timestamp 1667941163
transform 1 0 17848 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_70_193
timestamp 1667941163
transform 1 0 18860 0 1 40256
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_70_197
timestamp 1667941163
transform 1 0 19228 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_209
timestamp 1667941163
transform 1 0 20332 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_221
timestamp 1667941163
transform 1 0 21436 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_233
timestamp 1667941163
transform 1 0 22540 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_245
timestamp 1667941163
transform 1 0 23644 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_251
timestamp 1667941163
transform 1 0 24196 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_253
timestamp 1667941163
transform 1 0 24380 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_70_265
timestamp 1667941163
transform 1 0 25484 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_70_273
timestamp 1667941163
transform 1 0 26220 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_70_297
timestamp 1667941163
transform 1 0 28428 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_71_3
timestamp 1667941163
transform 1 0 1380 0 -1 41344
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_71_27
timestamp 1667941163
transform 1 0 3588 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_39
timestamp 1667941163
transform 1 0 4692 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_71_51
timestamp 1667941163
transform 1 0 5796 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_55
timestamp 1667941163
transform 1 0 6164 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_57
timestamp 1667941163
transform 1 0 6348 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_69
timestamp 1667941163
transform 1 0 7452 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_81
timestamp 1667941163
transform 1 0 8556 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_93
timestamp 1667941163
transform 1 0 9660 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_105
timestamp 1667941163
transform 1 0 10764 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_111
timestamp 1667941163
transform 1 0 11316 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_113
timestamp 1667941163
transform 1 0 11500 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_125
timestamp 1667941163
transform 1 0 12604 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_137
timestamp 1667941163
transform 1 0 13708 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_149
timestamp 1667941163
transform 1 0 14812 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_161
timestamp 1667941163
transform 1 0 15916 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_167
timestamp 1667941163
transform 1 0 16468 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_169
timestamp 1667941163
transform 1 0 16652 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_181
timestamp 1667941163
transform 1 0 17756 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_193
timestamp 1667941163
transform 1 0 18860 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_205
timestamp 1667941163
transform 1 0 19964 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_217
timestamp 1667941163
transform 1 0 21068 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_223
timestamp 1667941163
transform 1 0 21620 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_225
timestamp 1667941163
transform 1 0 21804 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_237
timestamp 1667941163
transform 1 0 22908 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_249
timestamp 1667941163
transform 1 0 24012 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_261
timestamp 1667941163
transform 1 0 25116 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_273
timestamp 1667941163
transform 1 0 26220 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_279
timestamp 1667941163
transform 1 0 26772 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_71_281
timestamp 1667941163
transform 1 0 26956 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_285
timestamp 1667941163
transform 1 0 27324 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_71_289
timestamp 1667941163
transform 1 0 27692 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_71_296
timestamp 1667941163
transform 1 0 28336 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_72_3
timestamp 1667941163
transform 1 0 1380 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_72_26
timestamp 1667941163
transform 1 0 3496 0 1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_72_29
timestamp 1667941163
transform 1 0 3772 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_41
timestamp 1667941163
transform 1 0 4876 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_53
timestamp 1667941163
transform 1 0 5980 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_65
timestamp 1667941163
transform 1 0 7084 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_77
timestamp 1667941163
transform 1 0 8188 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_83
timestamp 1667941163
transform 1 0 8740 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_85
timestamp 1667941163
transform 1 0 8924 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_97
timestamp 1667941163
transform 1 0 10028 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_109
timestamp 1667941163
transform 1 0 11132 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_121
timestamp 1667941163
transform 1 0 12236 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_133
timestamp 1667941163
transform 1 0 13340 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_139
timestamp 1667941163
transform 1 0 13892 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_141
timestamp 1667941163
transform 1 0 14076 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_153
timestamp 1667941163
transform 1 0 15180 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_165
timestamp 1667941163
transform 1 0 16284 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_177
timestamp 1667941163
transform 1 0 17388 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_189
timestamp 1667941163
transform 1 0 18492 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_195
timestamp 1667941163
transform 1 0 19044 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_197
timestamp 1667941163
transform 1 0 19228 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_209
timestamp 1667941163
transform 1 0 20332 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_221
timestamp 1667941163
transform 1 0 21436 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_233
timestamp 1667941163
transform 1 0 22540 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_245
timestamp 1667941163
transform 1 0 23644 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_251
timestamp 1667941163
transform 1 0 24196 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_253
timestamp 1667941163
transform 1 0 24380 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_72_265
timestamp 1667941163
transform 1 0 25484 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_72_273
timestamp 1667941163
transform 1 0 26220 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_72_297
timestamp 1667941163
transform 1 0 28428 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_73_3
timestamp 1667941163
transform 1 0 1380 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_73_9
timestamp 1667941163
transform 1 0 1932 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_73_18
timestamp 1667941163
transform 1 0 2760 0 -1 42432
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_73_25
timestamp 1667941163
transform 1 0 3404 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_37
timestamp 1667941163
transform 1 0 4508 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_49
timestamp 1667941163
transform 1 0 5612 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_55
timestamp 1667941163
transform 1 0 6164 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_57
timestamp 1667941163
transform 1 0 6348 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_69
timestamp 1667941163
transform 1 0 7452 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_81
timestamp 1667941163
transform 1 0 8556 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_93
timestamp 1667941163
transform 1 0 9660 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_105
timestamp 1667941163
transform 1 0 10764 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_111
timestamp 1667941163
transform 1 0 11316 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_113
timestamp 1667941163
transform 1 0 11500 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_125
timestamp 1667941163
transform 1 0 12604 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_137
timestamp 1667941163
transform 1 0 13708 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_149
timestamp 1667941163
transform 1 0 14812 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_161
timestamp 1667941163
transform 1 0 15916 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_167
timestamp 1667941163
transform 1 0 16468 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_169
timestamp 1667941163
transform 1 0 16652 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_181
timestamp 1667941163
transform 1 0 17756 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_193
timestamp 1667941163
transform 1 0 18860 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_205
timestamp 1667941163
transform 1 0 19964 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_217
timestamp 1667941163
transform 1 0 21068 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_223
timestamp 1667941163
transform 1 0 21620 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_225
timestamp 1667941163
transform 1 0 21804 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_237
timestamp 1667941163
transform 1 0 22908 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_249
timestamp 1667941163
transform 1 0 24012 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_261
timestamp 1667941163
transform 1 0 25116 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_273
timestamp 1667941163
transform 1 0 26220 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_279
timestamp 1667941163
transform 1 0 26772 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_73_281
timestamp 1667941163
transform 1 0 26956 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_73_292
timestamp 1667941163
transform 1 0 27968 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_298
timestamp 1667941163
transform 1 0 28520 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_74_3
timestamp 1667941163
transform 1 0 1380 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_74_26
timestamp 1667941163
transform 1 0 3496 0 1 42432
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_74_29
timestamp 1667941163
transform 1 0 3772 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_41
timestamp 1667941163
transform 1 0 4876 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_53
timestamp 1667941163
transform 1 0 5980 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_65
timestamp 1667941163
transform 1 0 7084 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_77
timestamp 1667941163
transform 1 0 8188 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_83
timestamp 1667941163
transform 1 0 8740 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_85
timestamp 1667941163
transform 1 0 8924 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_97
timestamp 1667941163
transform 1 0 10028 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_109
timestamp 1667941163
transform 1 0 11132 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_121
timestamp 1667941163
transform 1 0 12236 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_133
timestamp 1667941163
transform 1 0 13340 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_139
timestamp 1667941163
transform 1 0 13892 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_141
timestamp 1667941163
transform 1 0 14076 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_153
timestamp 1667941163
transform 1 0 15180 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_165
timestamp 1667941163
transform 1 0 16284 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_177
timestamp 1667941163
transform 1 0 17388 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_189
timestamp 1667941163
transform 1 0 18492 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_195
timestamp 1667941163
transform 1 0 19044 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_197
timestamp 1667941163
transform 1 0 19228 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_209
timestamp 1667941163
transform 1 0 20332 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_221
timestamp 1667941163
transform 1 0 21436 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_233
timestamp 1667941163
transform 1 0 22540 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_245
timestamp 1667941163
transform 1 0 23644 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_251
timestamp 1667941163
transform 1 0 24196 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_253
timestamp 1667941163
transform 1 0 24380 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_74_265
timestamp 1667941163
transform 1 0 25484 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_74_273
timestamp 1667941163
transform 1 0 26220 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_74_297
timestamp 1667941163
transform 1 0 28428 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_75_3
timestamp 1667941163
transform 1 0 1380 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_9
timestamp 1667941163
transform 1 0 1932 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_75_13
timestamp 1667941163
transform 1 0 2300 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_19
timestamp 1667941163
transform 1 0 2852 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_41
timestamp 1667941163
transform 1 0 4876 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_75_53
timestamp 1667941163
transform 1 0 5980 0 -1 43520
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_75_57
timestamp 1667941163
transform 1 0 6348 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_69
timestamp 1667941163
transform 1 0 7452 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_81
timestamp 1667941163
transform 1 0 8556 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_93
timestamp 1667941163
transform 1 0 9660 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_105
timestamp 1667941163
transform 1 0 10764 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_111
timestamp 1667941163
transform 1 0 11316 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_113
timestamp 1667941163
transform 1 0 11500 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_125
timestamp 1667941163
transform 1 0 12604 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_137
timestamp 1667941163
transform 1 0 13708 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_149
timestamp 1667941163
transform 1 0 14812 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_161
timestamp 1667941163
transform 1 0 15916 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_167
timestamp 1667941163
transform 1 0 16468 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_169
timestamp 1667941163
transform 1 0 16652 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_181
timestamp 1667941163
transform 1 0 17756 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_193
timestamp 1667941163
transform 1 0 18860 0 -1 43520
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_75_202
timestamp 1667941163
transform 1 0 19688 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_75_214
timestamp 1667941163
transform 1 0 20792 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_75_222
timestamp 1667941163
transform 1 0 21528 0 -1 43520
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_75_225
timestamp 1667941163
transform 1 0 21804 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_237
timestamp 1667941163
transform 1 0 22908 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_249
timestamp 1667941163
transform 1 0 24012 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_75_261
timestamp 1667941163
transform 1 0 25116 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_75_269
timestamp 1667941163
transform 1 0 25852 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_75_275
timestamp 1667941163
transform 1 0 26404 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_279
timestamp 1667941163
transform 1 0 26772 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_75_281
timestamp 1667941163
transform 1 0 26956 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_75_286
timestamp 1667941163
transform 1 0 27416 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_290
timestamp 1667941163
transform 1 0 27784 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_75_294
timestamp 1667941163
transform 1 0 28152 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_298
timestamp 1667941163
transform 1 0 28520 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_76_3
timestamp 1667941163
transform 1 0 1380 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_76_9
timestamp 1667941163
transform 1 0 1932 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_76_16
timestamp 1667941163
transform 1 0 2576 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_76_25
timestamp 1667941163
transform 1 0 3404 0 1 43520
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_76_29
timestamp 1667941163
transform 1 0 3772 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_41
timestamp 1667941163
transform 1 0 4876 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_53
timestamp 1667941163
transform 1 0 5980 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_65
timestamp 1667941163
transform 1 0 7084 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_77
timestamp 1667941163
transform 1 0 8188 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_83
timestamp 1667941163
transform 1 0 8740 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_85
timestamp 1667941163
transform 1 0 8924 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_97
timestamp 1667941163
transform 1 0 10028 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_109
timestamp 1667941163
transform 1 0 11132 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_121
timestamp 1667941163
transform 1 0 12236 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_133
timestamp 1667941163
transform 1 0 13340 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_139
timestamp 1667941163
transform 1 0 13892 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_141
timestamp 1667941163
transform 1 0 14076 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_153
timestamp 1667941163
transform 1 0 15180 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_165
timestamp 1667941163
transform 1 0 16284 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_177
timestamp 1667941163
transform 1 0 17388 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_189
timestamp 1667941163
transform 1 0 18492 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_195
timestamp 1667941163
transform 1 0 19044 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_76_197
timestamp 1667941163
transform 1 0 19228 0 1 43520
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_76_220
timestamp 1667941163
transform 1 0 21344 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_232
timestamp 1667941163
transform 1 0 22448 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_76_244
timestamp 1667941163
transform 1 0 23552 0 1 43520
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_76_253
timestamp 1667941163
transform 1 0 24380 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_76_265
timestamp 1667941163
transform 1 0 25484 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_76_294
timestamp 1667941163
transform 1 0 28152 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_76_298
timestamp 1667941163
transform 1 0 28520 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_77_3
timestamp 1667941163
transform 1 0 1380 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_9
timestamp 1667941163
transform 1 0 1932 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_77_13
timestamp 1667941163
transform 1 0 2300 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_19
timestamp 1667941163
transform 1 0 2852 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_23
timestamp 1667941163
transform 1 0 3220 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_35
timestamp 1667941163
transform 1 0 4324 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_77_47
timestamp 1667941163
transform 1 0 5428 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_77_55
timestamp 1667941163
transform 1 0 6164 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_57
timestamp 1667941163
transform 1 0 6348 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_69
timestamp 1667941163
transform 1 0 7452 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_81
timestamp 1667941163
transform 1 0 8556 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_93
timestamp 1667941163
transform 1 0 9660 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_105
timestamp 1667941163
transform 1 0 10764 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_111
timestamp 1667941163
transform 1 0 11316 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_113
timestamp 1667941163
transform 1 0 11500 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_125
timestamp 1667941163
transform 1 0 12604 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_77_137
timestamp 1667941163
transform 1 0 13708 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_141
timestamp 1667941163
transform 1 0 14076 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_145
timestamp 1667941163
transform 1 0 14444 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_77_157
timestamp 1667941163
transform 1 0 15548 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_77_165
timestamp 1667941163
transform 1 0 16284 0 -1 44608
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_77_169
timestamp 1667941163
transform 1 0 16652 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_181
timestamp 1667941163
transform 1 0 17756 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_193
timestamp 1667941163
transform 1 0 18860 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_205
timestamp 1667941163
transform 1 0 19964 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_217
timestamp 1667941163
transform 1 0 21068 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_223
timestamp 1667941163
transform 1 0 21620 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_225
timestamp 1667941163
transform 1 0 21804 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_237
timestamp 1667941163
transform 1 0 22908 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_77_249
timestamp 1667941163
transform 1 0 24012 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_77_278
timestamp 1667941163
transform 1 0 26680 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_77_281
timestamp 1667941163
transform 1 0 26956 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_77_286
timestamp 1667941163
transform 1 0 27416 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_77_293
timestamp 1667941163
transform 1 0 28060 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_78_3
timestamp 1667941163
transform 1 0 1380 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_78_12
timestamp 1667941163
transform 1 0 2208 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_78_20
timestamp 1667941163
transform 1 0 2944 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_78_25
timestamp 1667941163
transform 1 0 3404 0 1 44608
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_78_29
timestamp 1667941163
transform 1 0 3772 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_41
timestamp 1667941163
transform 1 0 4876 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_53
timestamp 1667941163
transform 1 0 5980 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_65
timestamp 1667941163
transform 1 0 7084 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_77
timestamp 1667941163
transform 1 0 8188 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_83
timestamp 1667941163
transform 1 0 8740 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_85
timestamp 1667941163
transform 1 0 8924 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_97
timestamp 1667941163
transform 1 0 10028 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_109
timestamp 1667941163
transform 1 0 11132 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_121
timestamp 1667941163
transform 1 0 12236 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_133
timestamp 1667941163
transform 1 0 13340 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_139
timestamp 1667941163
transform 1 0 13892 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_141
timestamp 1667941163
transform 1 0 14076 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_153
timestamp 1667941163
transform 1 0 15180 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_165
timestamp 1667941163
transform 1 0 16284 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_177
timestamp 1667941163
transform 1 0 17388 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_189
timestamp 1667941163
transform 1 0 18492 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_195
timestamp 1667941163
transform 1 0 19044 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_197
timestamp 1667941163
transform 1 0 19228 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_209
timestamp 1667941163
transform 1 0 20332 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_221
timestamp 1667941163
transform 1 0 21436 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_233
timestamp 1667941163
transform 1 0 22540 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_245
timestamp 1667941163
transform 1 0 23644 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_251
timestamp 1667941163
transform 1 0 24196 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_253
timestamp 1667941163
transform 1 0 24380 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_78_265
timestamp 1667941163
transform 1 0 25484 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_272
timestamp 1667941163
transform 1 0 26128 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_78_297
timestamp 1667941163
transform 1 0 28428 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_79_3
timestamp 1667941163
transform 1 0 1380 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_79_27
timestamp 1667941163
transform 1 0 3588 0 -1 45696
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_79_34
timestamp 1667941163
transform 1 0 4232 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_79_46
timestamp 1667941163
transform 1 0 5336 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_79_54
timestamp 1667941163
transform 1 0 6072 0 -1 45696
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_79_57
timestamp 1667941163
transform 1 0 6348 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_69
timestamp 1667941163
transform 1 0 7452 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_81
timestamp 1667941163
transform 1 0 8556 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_79_96
timestamp 1667941163
transform 1 0 9936 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_100
timestamp 1667941163
transform 1 0 10304 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_79_104
timestamp 1667941163
transform 1 0 10672 0 -1 45696
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_79_113
timestamp 1667941163
transform 1 0 11500 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_79_125
timestamp 1667941163
transform 1 0 12604 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_129
timestamp 1667941163
transform 1 0 12972 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_79_133
timestamp 1667941163
transform 1 0 13340 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_79_141
timestamp 1667941163
transform 1 0 14076 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_79_163
timestamp 1667941163
transform 1 0 16100 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_167
timestamp 1667941163
transform 1 0 16468 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_169
timestamp 1667941163
transform 1 0 16652 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_181
timestamp 1667941163
transform 1 0 17756 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_193
timestamp 1667941163
transform 1 0 18860 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_79_205
timestamp 1667941163
transform 1 0 19964 0 -1 45696
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_79_212
timestamp 1667941163
transform 1 0 20608 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_225
timestamp 1667941163
transform 1 0 21804 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_237
timestamp 1667941163
transform 1 0 22908 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_79_249
timestamp 1667941163
transform 1 0 24012 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_79_278
timestamp 1667941163
transform 1 0 26680 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_79_281
timestamp 1667941163
transform 1 0 26956 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_79_292
timestamp 1667941163
transform 1 0 27968 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_298
timestamp 1667941163
transform 1 0 28520 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_80_3
timestamp 1667941163
transform 1 0 1380 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_80_26
timestamp 1667941163
transform 1 0 3496 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_80_29
timestamp 1667941163
transform 1 0 3772 0 1 45696
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_80_52
timestamp 1667941163
transform 1 0 5888 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_80_64
timestamp 1667941163
transform 1 0 6992 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_80_72
timestamp 1667941163
transform 1 0 7728 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_80_76
timestamp 1667941163
transform 1 0 8096 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_80_85
timestamp 1667941163
transform 1 0 8924 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_80_89
timestamp 1667941163
transform 1 0 9292 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_80_93
timestamp 1667941163
transform 1 0 9660 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_100
timestamp 1667941163
transform 1 0 10304 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_107
timestamp 1667941163
transform 1 0 10948 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_80_132
timestamp 1667941163
transform 1 0 13248 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_80_141
timestamp 1667941163
transform 1 0 14076 0 1 45696
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_80_146
timestamp 1667941163
transform 1 0 14536 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_80_158
timestamp 1667941163
transform 1 0 15640 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_80_182
timestamp 1667941163
transform 1 0 17848 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_80_186
timestamp 1667941163
transform 1 0 18216 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_80_190
timestamp 1667941163
transform 1 0 18584 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_80_197
timestamp 1667941163
transform 1 0 19228 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_80_205
timestamp 1667941163
transform 1 0 19964 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_80_229
timestamp 1667941163
transform 1 0 22172 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_80_237
timestamp 1667941163
transform 1 0 22908 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_80_241
timestamp 1667941163
transform 1 0 23276 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_80_249
timestamp 1667941163
transform 1 0 24012 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_80_253
timestamp 1667941163
transform 1 0 24380 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_80_261
timestamp 1667941163
transform 1 0 25116 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_80_265
timestamp 1667941163
transform 1 0 25484 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_272
timestamp 1667941163
transform 1 0 26128 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_80_297
timestamp 1667941163
transform 1 0 28428 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_81_3
timestamp 1667941163
transform 1 0 1380 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_81_9
timestamp 1667941163
transform 1 0 1932 0 -1 46784
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_81_34
timestamp 1667941163
transform 1 0 4232 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_81_46
timestamp 1667941163
transform 1 0 5336 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_81_54
timestamp 1667941163
transform 1 0 6072 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_81_57
timestamp 1667941163
transform 1 0 6348 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_63
timestamp 1667941163
transform 1 0 6900 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_81_85
timestamp 1667941163
transform 1 0 8924 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_81_110
timestamp 1667941163
transform 1 0 11224 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_81_113
timestamp 1667941163
transform 1 0 11500 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_81_118
timestamp 1667941163
transform 1 0 11960 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_81_126
timestamp 1667941163
transform 1 0 12696 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_81_149
timestamp 1667941163
transform 1 0 14812 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_81_157
timestamp 1667941163
transform 1 0 15548 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_81_163
timestamp 1667941163
transform 1 0 16100 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_167
timestamp 1667941163
transform 1 0 16468 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_81_169
timestamp 1667941163
transform 1 0 16652 0 -1 46784
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_81_174
timestamp 1667941163
transform 1 0 17112 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_81_207
timestamp 1667941163
transform 1 0 20148 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_81_214
timestamp 1667941163
transform 1 0 20792 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_81_222
timestamp 1667941163
transform 1 0 21528 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_81_225
timestamp 1667941163
transform 1 0 21804 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_81_233
timestamp 1667941163
transform 1 0 22540 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_81_257
timestamp 1667941163
transform 1 0 24748 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_81_265
timestamp 1667941163
transform 1 0 25484 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_81_270
timestamp 1667941163
transform 1 0 25944 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_81_277
timestamp 1667941163
transform 1 0 26588 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_81_281
timestamp 1667941163
transform 1 0 26956 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_81_286
timestamp 1667941163
transform 1 0 27416 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_81_293
timestamp 1667941163
transform 1 0 28060 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_82_3
timestamp 1667941163
transform 1 0 1380 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_9
timestamp 1667941163
transform 1 0 1932 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_13
timestamp 1667941163
transform 1 0 2300 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_82_20
timestamp 1667941163
transform 1 0 2944 0 1 46784
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_82_29
timestamp 1667941163
transform 1 0 3772 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_82_41
timestamp 1667941163
transform 1 0 4876 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_82_49
timestamp 1667941163
transform 1 0 5612 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_82_54
timestamp 1667941163
transform 1 0 6072 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_82_57
timestamp 1667941163
transform 1 0 6348 0 1 46784
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_82_62
timestamp 1667941163
transform 1 0 6808 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_77
timestamp 1667941163
transform 1 0 8188 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_83
timestamp 1667941163
transform 1 0 8740 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_85
timestamp 1667941163
transform 1 0 8924 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_82_110
timestamp 1667941163
transform 1 0 11224 0 1 46784
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_82_113
timestamp 1667941163
transform 1 0 11500 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_82_125
timestamp 1667941163
transform 1 0 12604 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_82_132
timestamp 1667941163
transform 1 0 13248 0 1 46784
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_82_141
timestamp 1667941163
transform 1 0 14076 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_153
timestamp 1667941163
transform 1 0 15180 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_82_165
timestamp 1667941163
transform 1 0 16284 0 1 46784
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_82_169
timestamp 1667941163
transform 1 0 16652 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_181
timestamp 1667941163
transform 1 0 17756 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_82_190
timestamp 1667941163
transform 1 0 18584 0 1 46784
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_82_197
timestamp 1667941163
transform 1 0 19228 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_209
timestamp 1667941163
transform 1 0 20332 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_82_221
timestamp 1667941163
transform 1 0 21436 0 1 46784
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_82_225
timestamp 1667941163
transform 1 0 21804 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_240
timestamp 1667941163
transform 1 0 23184 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_246
timestamp 1667941163
transform 1 0 23736 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_82_250
timestamp 1667941163
transform 1 0 24104 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_82_253
timestamp 1667941163
transform 1 0 24380 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_82_278
timestamp 1667941163
transform 1 0 26680 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_82_281
timestamp 1667941163
transform 1 0 26956 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_82_287
timestamp 1667941163
transform 1 0 27508 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_294
timestamp 1667941163
transform 1 0 28152 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_82_298
timestamp 1667941163
transform 1 0 28520 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1667941163
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1667941163
transform -1 0 28888 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1667941163
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1667941163
transform -1 0 28888 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1667941163
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1667941163
transform -1 0 28888 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1667941163
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1667941163
transform -1 0 28888 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1667941163
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1667941163
transform -1 0 28888 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1667941163
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1667941163
transform -1 0 28888 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1667941163
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1667941163
transform -1 0 28888 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1667941163
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1667941163
transform -1 0 28888 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1667941163
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1667941163
transform -1 0 28888 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1667941163
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1667941163
transform -1 0 28888 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1667941163
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1667941163
transform -1 0 28888 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1667941163
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1667941163
transform -1 0 28888 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1667941163
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1667941163
transform -1 0 28888 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1667941163
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1667941163
transform -1 0 28888 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1667941163
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1667941163
transform -1 0 28888 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1667941163
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1667941163
transform -1 0 28888 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1667941163
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1667941163
transform -1 0 28888 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1667941163
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1667941163
transform -1 0 28888 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1667941163
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1667941163
transform -1 0 28888 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1667941163
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1667941163
transform -1 0 28888 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1667941163
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1667941163
transform -1 0 28888 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1667941163
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1667941163
transform -1 0 28888 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1667941163
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1667941163
transform -1 0 28888 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1667941163
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1667941163
transform -1 0 28888 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1667941163
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1667941163
transform -1 0 28888 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1667941163
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1667941163
transform -1 0 28888 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1667941163
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1667941163
transform -1 0 28888 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1667941163
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1667941163
transform -1 0 28888 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1667941163
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1667941163
transform -1 0 28888 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1667941163
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1667941163
transform -1 0 28888 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1667941163
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1667941163
transform -1 0 28888 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1667941163
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1667941163
transform -1 0 28888 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1667941163
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1667941163
transform -1 0 28888 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1667941163
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1667941163
transform -1 0 28888 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1667941163
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1667941163
transform -1 0 28888 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1667941163
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1667941163
transform -1 0 28888 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1667941163
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1667941163
transform -1 0 28888 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1667941163
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1667941163
transform -1 0 28888 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1667941163
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1667941163
transform -1 0 28888 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1667941163
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1667941163
transform -1 0 28888 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1667941163
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1667941163
transform -1 0 28888 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1667941163
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1667941163
transform -1 0 28888 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1667941163
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1667941163
transform -1 0 28888 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1667941163
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1667941163
transform -1 0 28888 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1667941163
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1667941163
transform -1 0 28888 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1667941163
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1667941163
transform -1 0 28888 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1667941163
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1667941163
transform -1 0 28888 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1667941163
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1667941163
transform -1 0 28888 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1667941163
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1667941163
transform -1 0 28888 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1667941163
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1667941163
transform -1 0 28888 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1667941163
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1667941163
transform -1 0 28888 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1667941163
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1667941163
transform -1 0 28888 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1667941163
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1667941163
transform -1 0 28888 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1667941163
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1667941163
transform -1 0 28888 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1667941163
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1667941163
transform -1 0 28888 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1667941163
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1667941163
transform -1 0 28888 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1667941163
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1667941163
transform -1 0 28888 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1667941163
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1667941163
transform -1 0 28888 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1667941163
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1667941163
transform -1 0 28888 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1667941163
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1667941163
transform -1 0 28888 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1667941163
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1667941163
transform -1 0 28888 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1667941163
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1667941163
transform -1 0 28888 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1667941163
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1667941163
transform -1 0 28888 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1667941163
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1667941163
transform -1 0 28888 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1667941163
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1667941163
transform -1 0 28888 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 1667941163
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 1667941163
transform -1 0 28888 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 1667941163
transform 1 0 1104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 1667941163
transform -1 0 28888 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_134
timestamp 1667941163
transform 1 0 1104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_135
timestamp 1667941163
transform -1 0 28888 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_136
timestamp 1667941163
transform 1 0 1104 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_137
timestamp 1667941163
transform -1 0 28888 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_138
timestamp 1667941163
transform 1 0 1104 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_139
timestamp 1667941163
transform -1 0 28888 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_140
timestamp 1667941163
transform 1 0 1104 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_141
timestamp 1667941163
transform -1 0 28888 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_142
timestamp 1667941163
transform 1 0 1104 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_143
timestamp 1667941163
transform -1 0 28888 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_144
timestamp 1667941163
transform 1 0 1104 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_145
timestamp 1667941163
transform -1 0 28888 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_146
timestamp 1667941163
transform 1 0 1104 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_147
timestamp 1667941163
transform -1 0 28888 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_148
timestamp 1667941163
transform 1 0 1104 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_149
timestamp 1667941163
transform -1 0 28888 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_150
timestamp 1667941163
transform 1 0 1104 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_151
timestamp 1667941163
transform -1 0 28888 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_152
timestamp 1667941163
transform 1 0 1104 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_153
timestamp 1667941163
transform -1 0 28888 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_154
timestamp 1667941163
transform 1 0 1104 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_155
timestamp 1667941163
transform -1 0 28888 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_156
timestamp 1667941163
transform 1 0 1104 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_157
timestamp 1667941163
transform -1 0 28888 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_158
timestamp 1667941163
transform 1 0 1104 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_159
timestamp 1667941163
transform -1 0 28888 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_160
timestamp 1667941163
transform 1 0 1104 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_161
timestamp 1667941163
transform -1 0 28888 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_162
timestamp 1667941163
transform 1 0 1104 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_163
timestamp 1667941163
transform -1 0 28888 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_164
timestamp 1667941163
transform 1 0 1104 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_165
timestamp 1667941163
transform -1 0 28888 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1667941163
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1667941163
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1667941163
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1667941163
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1667941163
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1667941163
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1667941163
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1667941163
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1667941163
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1667941163
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1667941163
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1667941163
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1667941163
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1667941163
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1667941163
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1667941163
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1667941163
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1667941163
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1667941163
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1667941163
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1667941163
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1667941163
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1667941163
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1667941163
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1667941163
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1667941163
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1667941163
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1667941163
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1667941163
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1667941163
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1667941163
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1667941163
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1667941163
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1667941163
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1667941163
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1667941163
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1667941163
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1667941163
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1667941163
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1667941163
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1667941163
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1667941163
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1667941163
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1667941163
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1667941163
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1667941163
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1667941163
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1667941163
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1667941163
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1667941163
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1667941163
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1667941163
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1667941163
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1667941163
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1667941163
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1667941163
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1667941163
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1667941163
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1667941163
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1667941163
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1667941163
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1667941163
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1667941163
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1667941163
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1667941163
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1667941163
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1667941163
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1667941163
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1667941163
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1667941163
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1667941163
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1667941163
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1667941163
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1667941163
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1667941163
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1667941163
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1667941163
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1667941163
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1667941163
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1667941163
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1667941163
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1667941163
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1667941163
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1667941163
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1667941163
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1667941163
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1667941163
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1667941163
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1667941163
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1667941163
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1667941163
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1667941163
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1667941163
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1667941163
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1667941163
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1667941163
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1667941163
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1667941163
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1667941163
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1667941163
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1667941163
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1667941163
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1667941163
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1667941163
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1667941163
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1667941163
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1667941163
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1667941163
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1667941163
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1667941163
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1667941163
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1667941163
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1667941163
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1667941163
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1667941163
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1667941163
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1667941163
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1667941163
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1667941163
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1667941163
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1667941163
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1667941163
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1667941163
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1667941163
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1667941163
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1667941163
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1667941163
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1667941163
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1667941163
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1667941163
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1667941163
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1667941163
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1667941163
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1667941163
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1667941163
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1667941163
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1667941163
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1667941163
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1667941163
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1667941163
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1667941163
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1667941163
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1667941163
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1667941163
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1667941163
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1667941163
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1667941163
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1667941163
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1667941163
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1667941163
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1667941163
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1667941163
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1667941163
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1667941163
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1667941163
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1667941163
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1667941163
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1667941163
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1667941163
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1667941163
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1667941163
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1667941163
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1667941163
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1667941163
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1667941163
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1667941163
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1667941163
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1667941163
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1667941163
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1667941163
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1667941163
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1667941163
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1667941163
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1667941163
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1667941163
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1667941163
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1667941163
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1667941163
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1667941163
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1667941163
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1667941163
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1667941163
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1667941163
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1667941163
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1667941163
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1667941163
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1667941163
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1667941163
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1667941163
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1667941163
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1667941163
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1667941163
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1667941163
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1667941163
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1667941163
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1667941163
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1667941163
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1667941163
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1667941163
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1667941163
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1667941163
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1667941163
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1667941163
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1667941163
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1667941163
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1667941163
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1667941163
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1667941163
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1667941163
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1667941163
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1667941163
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1667941163
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1667941163
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1667941163
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1667941163
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1667941163
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1667941163
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1667941163
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1667941163
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1667941163
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1667941163
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1667941163
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1667941163
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1667941163
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1667941163
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1667941163
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1667941163
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1667941163
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1667941163
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1667941163
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1667941163
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1667941163
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1667941163
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1667941163
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1667941163
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1667941163
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1667941163
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1667941163
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1667941163
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1667941163
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1667941163
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1667941163
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1667941163
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1667941163
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1667941163
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1667941163
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1667941163
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1667941163
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1667941163
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1667941163
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1667941163
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1667941163
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1667941163
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1667941163
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1667941163
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1667941163
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1667941163
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1667941163
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1667941163
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1667941163
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1667941163
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1667941163
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1667941163
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1667941163
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1667941163
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1667941163
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1667941163
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1667941163
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1667941163
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1667941163
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1667941163
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1667941163
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1667941163
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1667941163
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1667941163
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1667941163
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1667941163
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1667941163
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1667941163
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1667941163
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1667941163
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1667941163
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1667941163
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1667941163
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1667941163
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1667941163
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1667941163
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1667941163
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1667941163
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1667941163
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1667941163
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1667941163
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1667941163
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1667941163
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1667941163
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1667941163
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1667941163
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1667941163
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1667941163
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1667941163
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1667941163
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1667941163
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1667941163
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1667941163
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1667941163
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1667941163
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1667941163
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1667941163
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1667941163
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1667941163
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1667941163
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1667941163
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1667941163
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1667941163
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1667941163
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1667941163
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1667941163
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1667941163
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1667941163
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1667941163
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1667941163
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1667941163
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1667941163
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1667941163
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1667941163
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1667941163
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1667941163
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1667941163
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1667941163
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1667941163
transform 1 0 6256 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1667941163
transform 1 0 11408 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1667941163
transform 1 0 16560 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1667941163
transform 1 0 21712 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1667941163
transform 1 0 26864 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1667941163
transform 1 0 3680 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1667941163
transform 1 0 8832 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1667941163
transform 1 0 13984 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1667941163
transform 1 0 19136 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1667941163
transform 1 0 24288 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1667941163
transform 1 0 6256 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1667941163
transform 1 0 11408 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1667941163
transform 1 0 16560 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1667941163
transform 1 0 21712 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1667941163
transform 1 0 26864 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1667941163
transform 1 0 3680 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1667941163
transform 1 0 8832 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1667941163
transform 1 0 13984 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1667941163
transform 1 0 19136 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1667941163
transform 1 0 24288 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1667941163
transform 1 0 6256 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1667941163
transform 1 0 11408 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1667941163
transform 1 0 16560 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1667941163
transform 1 0 21712 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1667941163
transform 1 0 26864 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1667941163
transform 1 0 3680 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1667941163
transform 1 0 8832 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1667941163
transform 1 0 13984 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1667941163
transform 1 0 19136 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1667941163
transform 1 0 24288 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1667941163
transform 1 0 6256 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1667941163
transform 1 0 11408 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1667941163
transform 1 0 16560 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1667941163
transform 1 0 21712 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1667941163
transform 1 0 26864 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1667941163
transform 1 0 3680 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1667941163
transform 1 0 8832 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1667941163
transform 1 0 13984 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1667941163
transform 1 0 19136 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1667941163
transform 1 0 24288 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1667941163
transform 1 0 6256 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1667941163
transform 1 0 11408 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1667941163
transform 1 0 16560 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1667941163
transform 1 0 21712 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1667941163
transform 1 0 26864 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1667941163
transform 1 0 3680 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1667941163
transform 1 0 8832 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1667941163
transform 1 0 13984 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1667941163
transform 1 0 19136 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1667941163
transform 1 0 24288 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1667941163
transform 1 0 6256 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1667941163
transform 1 0 11408 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1667941163
transform 1 0 16560 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1667941163
transform 1 0 21712 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1667941163
transform 1 0 26864 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1667941163
transform 1 0 3680 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1667941163
transform 1 0 8832 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1667941163
transform 1 0 13984 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1667941163
transform 1 0 19136 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1667941163
transform 1 0 24288 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1667941163
transform 1 0 6256 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1667941163
transform 1 0 11408 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1667941163
transform 1 0 16560 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1667941163
transform 1 0 21712 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1667941163
transform 1 0 26864 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1667941163
transform 1 0 3680 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1667941163
transform 1 0 8832 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1667941163
transform 1 0 13984 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1667941163
transform 1 0 19136 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1667941163
transform 1 0 24288 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1667941163
transform 1 0 6256 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1667941163
transform 1 0 11408 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1667941163
transform 1 0 16560 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1667941163
transform 1 0 21712 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1667941163
transform 1 0 26864 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1667941163
transform 1 0 3680 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1667941163
transform 1 0 8832 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1667941163
transform 1 0 13984 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1667941163
transform 1 0 19136 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1667941163
transform 1 0 24288 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1667941163
transform 1 0 6256 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1667941163
transform 1 0 11408 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1667941163
transform 1 0 16560 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1667941163
transform 1 0 21712 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1667941163
transform 1 0 26864 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1667941163
transform 1 0 3680 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1667941163
transform 1 0 6256 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1667941163
transform 1 0 8832 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1667941163
transform 1 0 11408 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1667941163
transform 1 0 13984 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1667941163
transform 1 0 16560 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1667941163
transform 1 0 19136 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1667941163
transform 1 0 21712 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1667941163
transform 1 0 24288 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1667941163
transform 1 0 26864 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_8  _0470_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 3312 0 -1 36992
box -38 -48 1050 592
use sky130_fd_sc_hd__buf_8  _0471_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 4048 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_6  _0472_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 25208 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0473_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 2116 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0474_
timestamp 1667941163
transform -1 0 2576 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0475_
timestamp 1667941163
transform -1 0 2116 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0476_
timestamp 1667941163
transform -1 0 2024 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0477_
timestamp 1667941163
transform 1 0 27692 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0478_
timestamp 1667941163
transform -1 0 2024 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0479_
timestamp 1667941163
transform 1 0 27692 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0480_
timestamp 1667941163
transform -1 0 2484 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0481_
timestamp 1667941163
transform -1 0 27416 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0482_
timestamp 1667941163
transform 1 0 27692 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _0483_
timestamp 1667941163
transform 1 0 11868 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0484_
timestamp 1667941163
transform -1 0 13340 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0485_
timestamp 1667941163
transform 1 0 27692 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0486_
timestamp 1667941163
transform 1 0 27600 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0487_
timestamp 1667941163
transform -1 0 10304 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0488_
timestamp 1667941163
transform 1 0 9384 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0489_
timestamp 1667941163
transform -1 0 4876 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0490_
timestamp 1667941163
transform -1 0 2760 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0491_
timestamp 1667941163
transform 1 0 27692 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0492_
timestamp 1667941163
transform -1 0 2944 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0493_
timestamp 1667941163
transform 1 0 18308 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _0494_
timestamp 1667941163
transform -1 0 3220 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0495_
timestamp 1667941163
transform 1 0 10488 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0496_
timestamp 1667941163
transform -1 0 27508 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0497_
timestamp 1667941163
transform -1 0 2208 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0498_
timestamp 1667941163
transform -1 0 2576 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0499_
timestamp 1667941163
transform -1 0 27508 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0500_
timestamp 1667941163
transform 1 0 27784 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0501_
timestamp 1667941163
transform 1 0 28060 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0502_
timestamp 1667941163
transform -1 0 2208 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0503_
timestamp 1667941163
transform 1 0 3956 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0504_
timestamp 1667941163
transform 1 0 27784 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _0505_
timestamp 1667941163
transform -1 0 4784 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0506_
timestamp 1667941163
transform -1 0 27416 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0507_
timestamp 1667941163
transform -1 0 23276 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0508_
timestamp 1667941163
transform 1 0 18676 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0509_
timestamp 1667941163
transform 1 0 27600 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0510_
timestamp 1667941163
transform -1 0 2300 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0511_
timestamp 1667941163
transform -1 0 27508 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0512_
timestamp 1667941163
transform -1 0 2300 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0513_
timestamp 1667941163
transform 1 0 2576 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0514_
timestamp 1667941163
transform 1 0 27692 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0515_
timestamp 1667941163
transform -1 0 27508 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _0516_
timestamp 1667941163
transform 1 0 3588 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0517_
timestamp 1667941163
transform -1 0 27416 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0518_
timestamp 1667941163
transform 1 0 23828 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0519_
timestamp 1667941163
transform -1 0 27508 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0520_
timestamp 1667941163
transform 1 0 22172 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0521_
timestamp 1667941163
transform -1 0 6808 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0522_
timestamp 1667941163
transform -1 0 1932 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0523_
timestamp 1667941163
transform 1 0 16652 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0524_
timestamp 1667941163
transform -1 0 2300 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0525_
timestamp 1667941163
transform 1 0 27416 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0526_
timestamp 1667941163
transform 1 0 2392 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _0527_
timestamp 1667941163
transform -1 0 5060 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0528_
timestamp 1667941163
transform -1 0 27508 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0529_
timestamp 1667941163
transform -1 0 2024 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0530_
timestamp 1667941163
transform 1 0 27416 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0531_
timestamp 1667941163
transform 1 0 25852 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0532_
timestamp 1667941163
transform 1 0 27784 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0533_
timestamp 1667941163
transform 1 0 18124 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0534_
timestamp 1667941163
transform 1 0 27784 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0535_
timestamp 1667941163
transform -1 0 3404 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0536_
timestamp 1667941163
transform 1 0 10672 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0537_
timestamp 1667941163
transform -1 0 2484 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _0538_
timestamp 1667941163
transform 1 0 2392 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0539_
timestamp 1667941163
transform -1 0 27416 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0540_
timestamp 1667941163
transform 1 0 27692 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0541_
timestamp 1667941163
transform -1 0 2300 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0542_
timestamp 1667941163
transform 1 0 21252 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0543_
timestamp 1667941163
transform -1 0 27508 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0544_
timestamp 1667941163
transform 1 0 15824 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0545_
timestamp 1667941163
transform 1 0 2300 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0546_
timestamp 1667941163
transform 1 0 5336 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0547_
timestamp 1667941163
transform -1 0 2300 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0548_
timestamp 1667941163
transform 1 0 20332 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _0549_
timestamp 1667941163
transform 1 0 3956 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0550_
timestamp 1667941163
transform 1 0 27968 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0551_
timestamp 1667941163
transform -1 0 8096 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0552_
timestamp 1667941163
transform 1 0 12788 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0553_
timestamp 1667941163
transform -1 0 26588 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0554_
timestamp 1667941163
transform -1 0 2208 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0555_
timestamp 1667941163
transform 1 0 26404 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0556_
timestamp 1667941163
transform 1 0 13524 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0557_
timestamp 1667941163
transform 1 0 9660 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0558_
timestamp 1667941163
transform -1 0 2300 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0559_
timestamp 1667941163
transform -1 0 2576 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _0560_
timestamp 1667941163
transform 1 0 5060 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0561_
timestamp 1667941163
transform 1 0 27784 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0562_
timestamp 1667941163
transform -1 0 27416 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0563_
timestamp 1667941163
transform 1 0 8372 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0564_
timestamp 1667941163
transform 1 0 10948 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0565_
timestamp 1667941163
transform -1 0 27416 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0566_
timestamp 1667941163
transform -1 0 3036 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0567_
timestamp 1667941163
transform 1 0 25852 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0568_
timestamp 1667941163
transform 1 0 27416 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0569_
timestamp 1667941163
transform 1 0 12788 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0570_
timestamp 1667941163
transform 1 0 25852 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _0571_
timestamp 1667941163
transform 1 0 3956 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0572_
timestamp 1667941163
transform -1 0 5428 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0573_
timestamp 1667941163
transform -1 0 26036 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0574_
timestamp 1667941163
transform 1 0 21252 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0575_
timestamp 1667941163
transform 1 0 19412 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0576_
timestamp 1667941163
transform 1 0 14352 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0577_
timestamp 1667941163
transform 1 0 26128 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0578_
timestamp 1667941163
transform -1 0 4232 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0579_
timestamp 1667941163
transform 1 0 27140 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0580_
timestamp 1667941163
transform 1 0 14168 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0581_
timestamp 1667941163
transform 1 0 9292 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0582_
timestamp 1667941163
transform 1 0 27140 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0583_
timestamp 1667941163
transform -1 0 4416 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0584_
timestamp 1667941163
transform 1 0 26312 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0585_
timestamp 1667941163
transform -1 0 3312 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0586_
timestamp 1667941163
transform -1 0 4692 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0587_
timestamp 1667941163
transform -1 0 8280 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0588_
timestamp 1667941163
transform -1 0 21344 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0589_
timestamp 1667941163
transform 1 0 27140 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _0590_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 21252 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0591_
timestamp 1667941163
transform -1 0 17112 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0592_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 19964 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_2  _0593_
timestamp 1667941163
transform 1 0 20700 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _0594_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 12512 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _0595_
timestamp 1667941163
transform 1 0 20056 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _0596_
timestamp 1667941163
transform 1 0 14444 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0597_
timestamp 1667941163
transform -1 0 13800 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0598_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 13248 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _0599_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 14996 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_1  _0600_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 16376 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0601_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 15732 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__or2b_1  _0602_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 16100 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0603_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 16008 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__o21bai_1  _0604_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 12880 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0605_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 14260 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0606_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 14168 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0607_
timestamp 1667941163
transform 1 0 14904 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _0608_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 14260 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0609_
timestamp 1667941163
transform -1 0 15272 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0610_
timestamp 1667941163
transform 1 0 15732 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0611_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 24840 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _0612_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 14444 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _0613_
timestamp 1667941163
transform 1 0 13248 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _0614_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 26036 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _0615_
timestamp 1667941163
transform -1 0 22816 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0616_
timestamp 1667941163
transform -1 0 21436 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0617_
timestamp 1667941163
transform 1 0 26404 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0618_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 24932 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _0619_
timestamp 1667941163
transform 1 0 21988 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0620_
timestamp 1667941163
transform 1 0 21988 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0621_
timestamp 1667941163
transform -1 0 23092 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0622_
timestamp 1667941163
transform -1 0 19780 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _0623_
timestamp 1667941163
transform 1 0 20424 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0624_
timestamp 1667941163
transform -1 0 19964 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0625_
timestamp 1667941163
transform 1 0 19412 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0626_
timestamp 1667941163
transform 1 0 20332 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0627_
timestamp 1667941163
transform -1 0 19872 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0628_
timestamp 1667941163
transform -1 0 19688 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0629_
timestamp 1667941163
transform 1 0 21068 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0630_
timestamp 1667941163
transform 1 0 20700 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0631_
timestamp 1667941163
transform 1 0 21528 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0632_
timestamp 1667941163
transform 1 0 20700 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0633_
timestamp 1667941163
transform 1 0 20516 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0634_
timestamp 1667941163
transform 1 0 20700 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0635_
timestamp 1667941163
transform 1 0 20424 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0636_
timestamp 1667941163
transform -1 0 20148 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0637_
timestamp 1667941163
transform 1 0 19688 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0638_
timestamp 1667941163
transform 1 0 20240 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0639_
timestamp 1667941163
transform -1 0 19872 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0640_
timestamp 1667941163
transform -1 0 18952 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0641_
timestamp 1667941163
transform 1 0 20516 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0642_
timestamp 1667941163
transform -1 0 20240 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0643_
timestamp 1667941163
transform 1 0 19780 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _0644_
timestamp 1667941163
transform 1 0 18216 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  _0645_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 15732 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _0646_
timestamp 1667941163
transform -1 0 16284 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _0647_
timestamp 1667941163
transform 1 0 16652 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0648_
timestamp 1667941163
transform -1 0 16376 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0649_
timestamp 1667941163
transform -1 0 16284 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _0650_
timestamp 1667941163
transform 1 0 15916 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0651_
timestamp 1667941163
transform -1 0 16744 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0652_
timestamp 1667941163
transform 1 0 22908 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _0653_
timestamp 1667941163
transform 1 0 22724 0 1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0654_
timestamp 1667941163
transform 1 0 22816 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0655_
timestamp 1667941163
transform -1 0 26680 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _0656_
timestamp 1667941163
transform 1 0 27140 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0657_
timestamp 1667941163
transform 1 0 26220 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0658_
timestamp 1667941163
transform 1 0 15548 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0659_
timestamp 1667941163
transform 1 0 15548 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0660_
timestamp 1667941163
transform -1 0 17112 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0661_
timestamp 1667941163
transform 1 0 15180 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _0662_
timestamp 1667941163
transform 1 0 15456 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0663_
timestamp 1667941163
transform -1 0 16284 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0664_
timestamp 1667941163
transform -1 0 16100 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0665_
timestamp 1667941163
transform 1 0 15456 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0666_
timestamp 1667941163
transform -1 0 16284 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0667_
timestamp 1667941163
transform -1 0 16008 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _0668_
timestamp 1667941163
transform 1 0 15640 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0669_
timestamp 1667941163
transform -1 0 17112 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0670_
timestamp 1667941163
transform 1 0 16836 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0671_
timestamp 1667941163
transform -1 0 17020 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0672_
timestamp 1667941163
transform -1 0 16376 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0673_
timestamp 1667941163
transform 1 0 27140 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0674_
timestamp 1667941163
transform 1 0 27140 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0675_
timestamp 1667941163
transform 1 0 27968 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0676_
timestamp 1667941163
transform 1 0 15364 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _0677_
timestamp 1667941163
transform 1 0 15640 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0678_
timestamp 1667941163
transform -1 0 17112 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0679_
timestamp 1667941163
transform 1 0 25300 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0680_
timestamp 1667941163
transform -1 0 25852 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0681_
timestamp 1667941163
transform -1 0 24840 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0682_
timestamp 1667941163
transform -1 0 19872 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0683_
timestamp 1667941163
transform -1 0 18952 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_1  _0684_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 18400 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0685_
timestamp 1667941163
transform 1 0 19504 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0686_
timestamp 1667941163
transform 1 0 20792 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0687_
timestamp 1667941163
transform -1 0 19780 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0688_
timestamp 1667941163
transform -1 0 16192 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0689_
timestamp 1667941163
transform -1 0 17848 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__a22oi_1  _0690_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 15548 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0691_
timestamp 1667941163
transform -1 0 20700 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0692_
timestamp 1667941163
transform 1 0 20148 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _0693_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 19412 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0694_
timestamp 1667941163
transform 1 0 21252 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _0695_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 20424 0 1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0696_
timestamp 1667941163
transform -1 0 20884 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _0697_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 20056 0 1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _0698_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 19504 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0699_
timestamp 1667941163
transform -1 0 17204 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _0700_
timestamp 1667941163
transform -1 0 16376 0 -1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0701_
timestamp 1667941163
transform 1 0 18216 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _0702_
timestamp 1667941163
transform 1 0 17204 0 1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0703_
timestamp 1667941163
transform 1 0 18216 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0704_
timestamp 1667941163
transform -1 0 19688 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _0705_
timestamp 1667941163
transform 1 0 16008 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _0706_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 18860 0 -1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _0707_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 16928 0 1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0708_
timestamp 1667941163
transform -1 0 16560 0 1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _0709_
timestamp 1667941163
transform 1 0 16008 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__a32o_1  _0710_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 17572 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0711_
timestamp 1667941163
transform -1 0 18124 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0712_
timestamp 1667941163
transform 1 0 17756 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _0713_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 18860 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0714_
timestamp 1667941163
transform -1 0 18400 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0715_
timestamp 1667941163
transform 1 0 16100 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _0716_
timestamp 1667941163
transform 1 0 16836 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0717_
timestamp 1667941163
transform -1 0 18768 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__o2111a_1  _0718_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 16836 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__and3b_1  _0719_
timestamp 1667941163
transform 1 0 16836 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0720_
timestamp 1667941163
transform -1 0 17204 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0721_
timestamp 1667941163
transform 1 0 19412 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _0722_
timestamp 1667941163
transform 1 0 19412 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _0723_
timestamp 1667941163
transform 1 0 27140 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _0724_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 26680 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _0725_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 26128 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__clkinv_2  _0726_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 24932 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0727_
timestamp 1667941163
transform -1 0 23552 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _0728_
timestamp 1667941163
transform -1 0 22724 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _0729_
timestamp 1667941163
transform -1 0 23736 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _0730_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 23828 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0731_
timestamp 1667941163
transform 1 0 23736 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0732_
timestamp 1667941163
transform -1 0 23000 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0733_
timestamp 1667941163
transform -1 0 23368 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _0734_
timestamp 1667941163
transform -1 0 22172 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0735_
timestamp 1667941163
transform 1 0 22080 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0736_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 23000 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0737_
timestamp 1667941163
transform 1 0 23092 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_1  _0738_
timestamp 1667941163
transform 1 0 21988 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _0739_
timestamp 1667941163
transform 1 0 21988 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0740_
timestamp 1667941163
transform 1 0 22816 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_1  _0741_
timestamp 1667941163
transform 1 0 21988 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _0742_
timestamp 1667941163
transform 1 0 21160 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0743_
timestamp 1667941163
transform 1 0 22724 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_1  _0744_
timestamp 1667941163
transform 1 0 22264 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _0745_
timestamp 1667941163
transform 1 0 22264 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0746_
timestamp 1667941163
transform 1 0 23460 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_1  _0747_
timestamp 1667941163
transform 1 0 22172 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _0748_
timestamp 1667941163
transform 1 0 21528 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0749_
timestamp 1667941163
transform -1 0 25484 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _0750_
timestamp 1667941163
transform -1 0 25208 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _0751_
timestamp 1667941163
transform 1 0 24564 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _0752_
timestamp 1667941163
transform 1 0 25668 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _0753_
timestamp 1667941163
transform 1 0 24196 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _0754_
timestamp 1667941163
transform -1 0 24840 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _0755_
timestamp 1667941163
transform 1 0 22356 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0756_
timestamp 1667941163
transform -1 0 22816 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__a41o_1  _0757_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 23644 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _0758_
timestamp 1667941163
transform 1 0 23092 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__a41o_1  _0759_
timestamp 1667941163
transform 1 0 22172 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0760_
timestamp 1667941163
transform 1 0 22264 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _0761_
timestamp 1667941163
transform 1 0 23276 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _0762_
timestamp 1667941163
transform 1 0 21988 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _0763_
timestamp 1667941163
transform 1 0 20608 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0764_
timestamp 1667941163
transform 1 0 19780 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _0765_
timestamp 1667941163
transform -1 0 19412 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _0766_
timestamp 1667941163
transform 1 0 19412 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0767_
timestamp 1667941163
transform 1 0 21160 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0768_
timestamp 1667941163
transform -1 0 20792 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _0769_
timestamp 1667941163
transform 1 0 20424 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__o32a_1  _0770_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 19872 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _0771_
timestamp 1667941163
transform -1 0 18952 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0772_
timestamp 1667941163
transform 1 0 20792 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0773_
timestamp 1667941163
transform -1 0 20792 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__o32a_1  _0774_
timestamp 1667941163
transform -1 0 20884 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _0775_
timestamp 1667941163
transform 1 0 21068 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0776_
timestamp 1667941163
transform 1 0 19872 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0777_
timestamp 1667941163
transform -1 0 19872 0 -1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__o32a_1  _0778_
timestamp 1667941163
transform 1 0 19504 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _0779_
timestamp 1667941163
transform -1 0 19320 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0780_
timestamp 1667941163
transform 1 0 18584 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0781_
timestamp 1667941163
transform -1 0 19504 0 -1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__o32a_1  _0782_
timestamp 1667941163
transform 1 0 18216 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _0783_
timestamp 1667941163
transform -1 0 18400 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0784_
timestamp 1667941163
transform 1 0 17480 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0785_
timestamp 1667941163
transform -1 0 18584 0 -1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__o32a_1  _0786_
timestamp 1667941163
transform 1 0 17020 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _0787_
timestamp 1667941163
transform -1 0 17204 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0788_
timestamp 1667941163
transform -1 0 16376 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0789_
timestamp 1667941163
transform 1 0 16560 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__o32a_1  _0790_
timestamp 1667941163
transform 1 0 16836 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _0791_
timestamp 1667941163
transform -1 0 16928 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0792_
timestamp 1667941163
transform -1 0 17112 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0793_
timestamp 1667941163
transform -1 0 16376 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__o32a_1  _0794_
timestamp 1667941163
transform -1 0 17020 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _0795_
timestamp 1667941163
transform 1 0 17388 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0796_
timestamp 1667941163
transform -1 0 15916 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0797_
timestamp 1667941163
transform 1 0 16284 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__o32a_1  _0798_
timestamp 1667941163
transform 1 0 16836 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _0799_
timestamp 1667941163
transform -1 0 16284 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0800_
timestamp 1667941163
transform 1 0 18308 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0801_
timestamp 1667941163
transform -1 0 17756 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__o32a_1  _0802_
timestamp 1667941163
transform 1 0 17204 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _0803_
timestamp 1667941163
transform -1 0 17388 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0804_
timestamp 1667941163
transform -1 0 19872 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0805_
timestamp 1667941163
transform -1 0 19044 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__o32a_1  _0806_
timestamp 1667941163
transform 1 0 18492 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _0807_
timestamp 1667941163
transform 1 0 18492 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__o211ai_1  _0808_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 19688 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0809_
timestamp 1667941163
transform 1 0 18676 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0810_
timestamp 1667941163
transform 1 0 17848 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0811_
timestamp 1667941163
transform 1 0 18676 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0812_
timestamp 1667941163
transform -1 0 24012 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0813_
timestamp 1667941163
transform 1 0 25392 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0814_
timestamp 1667941163
transform -1 0 25116 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _0815_
timestamp 1667941163
transform -1 0 25944 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0816_
timestamp 1667941163
transform -1 0 25116 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0817_
timestamp 1667941163
transform -1 0 24288 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0818_
timestamp 1667941163
transform -1 0 25024 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _0819_
timestamp 1667941163
transform -1 0 24564 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _0820_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 24932 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__o221ai_1  _0821_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 24932 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _0822_
timestamp 1667941163
transform -1 0 25668 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _0823_
timestamp 1667941163
transform -1 0 23828 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0824_
timestamp 1667941163
transform 1 0 23460 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _0825_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 23644 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__o32a_1  _0826_
timestamp 1667941163
transform 1 0 23644 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0827_
timestamp 1667941163
transform 1 0 23828 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _0828_
timestamp 1667941163
transform -1 0 25300 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _0829_
timestamp 1667941163
transform 1 0 27140 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _0830_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 25392 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0831_
timestamp 1667941163
transform 1 0 23644 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0832_
timestamp 1667941163
transform -1 0 24104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _0833_
timestamp 1667941163
transform 1 0 24472 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0834_
timestamp 1667941163
transform 1 0 24656 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _0835_
timestamp 1667941163
transform 1 0 25024 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _0836_
timestamp 1667941163
transform 1 0 24564 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _0837_
timestamp 1667941163
transform 1 0 25116 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__a21bo_1  _0838_
timestamp 1667941163
transform -1 0 25668 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__or3b_1  _0839_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 24564 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _0840_
timestamp 1667941163
transform -1 0 25852 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _0841_
timestamp 1667941163
transform -1 0 24748 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0842_
timestamp 1667941163
transform -1 0 23828 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _0843_
timestamp 1667941163
transform 1 0 24564 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _0844_
timestamp 1667941163
transform 1 0 25668 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _0845_
timestamp 1667941163
transform -1 0 26588 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0846_
timestamp 1667941163
transform -1 0 24840 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__o21ba_1  _0847_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 24564 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_1  _0848_
timestamp 1667941163
transform 1 0 23092 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _0849_
timestamp 1667941163
transform -1 0 22724 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _0850_
timestamp 1667941163
transform 1 0 22632 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_2  _0851_
timestamp 1667941163
transform 1 0 23092 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__o2bb2a_1  _0852_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 23000 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _0853_
timestamp 1667941163
transform -1 0 22264 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _0854_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 23460 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__o21ba_1  _0855_
timestamp 1667941163
transform 1 0 23368 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_2  _0856_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 21252 0 1 33728
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _0857_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 23368 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0858_
timestamp 1667941163
transform 1 0 19044 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0859_
timestamp 1667941163
transform 1 0 19412 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0860_
timestamp 1667941163
transform 1 0 21252 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0861_
timestamp 1667941163
transform 1 0 20424 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0862_
timestamp 1667941163
transform 1 0 19412 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0863_
timestamp 1667941163
transform 1 0 19228 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0864_
timestamp 1667941163
transform 1 0 19412 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0865_
timestamp 1667941163
transform -1 0 28336 0 1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0866_
timestamp 1667941163
transform -1 0 26680 0 -1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0867_
timestamp 1667941163
transform 1 0 24656 0 1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0868_
timestamp 1667941163
transform 1 0 16836 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0869_
timestamp 1667941163
transform 1 0 17020 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0870_
timestamp 1667941163
transform 1 0 22540 0 -1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0871_
timestamp 1667941163
transform -1 0 26496 0 1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0872_
timestamp 1667941163
transform 1 0 16836 0 1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0873_
timestamp 1667941163
transform 1 0 16836 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0874_
timestamp 1667941163
transform -1 0 18492 0 -1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0875_
timestamp 1667941163
transform -1 0 18308 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0876_
timestamp 1667941163
transform 1 0 16836 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0877_
timestamp 1667941163
transform 1 0 26312 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0878_
timestamp 1667941163
transform 1 0 16836 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0879_
timestamp 1667941163
transform 1 0 25208 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _0880_
timestamp 1667941163
transform 1 0 23552 0 -1 17408
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _0881_
timestamp 1667941163
transform -1 0 24012 0 1 27200
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _0882_
timestamp 1667941163
transform -1 0 23552 0 -1 19584
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _0883_
timestamp 1667941163
transform -1 0 22724 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0884_
timestamp 1667941163
transform 1 0 20608 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0885_
timestamp 1667941163
transform -1 0 23460 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0886_
timestamp 1667941163
transform -1 0 23092 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _0887_
timestamp 1667941163
transform 1 0 24564 0 1 14144
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _0888_
timestamp 1667941163
transform 1 0 24196 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0889_
timestamp 1667941163
transform -1 0 23920 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0890_
timestamp 1667941163
transform 1 0 21988 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0891_
timestamp 1667941163
transform 1 0 19412 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0892_
timestamp 1667941163
transform 1 0 19320 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0893_
timestamp 1667941163
transform -1 0 22724 0 1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0894_
timestamp 1667941163
transform 1 0 19412 0 1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0895_
timestamp 1667941163
transform 1 0 18124 0 -1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0896_
timestamp 1667941163
transform 1 0 17020 0 -1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0897_
timestamp 1667941163
transform -1 0 18768 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0898_
timestamp 1667941163
transform -1 0 18952 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0899_
timestamp 1667941163
transform 1 0 16836 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _0900_
timestamp 1667941163
transform 1 0 17388 0 -1 25024
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _0901_
timestamp 1667941163
transform 1 0 18860 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0902_
timestamp 1667941163
transform 1 0 18216 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0903_
timestamp 1667941163
transform 1 0 25208 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _0904_
timestamp 1667941163
transform 1 0 25116 0 -1 22848
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _0905_
timestamp 1667941163
transform -1 0 27416 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0906_
timestamp 1667941163
transform 1 0 25208 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _0907_
timestamp 1667941163
transform 1 0 24564 0 1 17408
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _0908_
timestamp 1667941163
transform 1 0 21160 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0909_
timestamp 1667941163
transform 1 0 23552 0 -1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__ebufn_8  _1001_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 5704 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1001__17 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 5060 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1002__18
timestamp 1667941163
transform -1 0 1932 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1002_
timestamp 1667941163
transform 1 0 1564 0 1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1003__19
timestamp 1667941163
transform 1 0 16008 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1003_
timestamp 1667941163
transform 1 0 16836 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1004__20
timestamp 1667941163
transform -1 0 2024 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1004_
timestamp 1667941163
transform 1 0 1656 0 -1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1005__21
timestamp 1667941163
transform -1 0 27876 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1005_
timestamp 1667941163
transform -1 0 26680 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1006_
timestamp 1667941163
transform 1 0 2944 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1006__22
timestamp 1667941163
transform -1 0 3220 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1007__23
timestamp 1667941163
transform -1 0 28152 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1007_
timestamp 1667941163
transform 1 0 26496 0 1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1008__24
timestamp 1667941163
transform -1 0 1840 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1008_
timestamp 1667941163
transform 1 0 1564 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1009__25
timestamp 1667941163
transform 1 0 28060 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1009_
timestamp 1667941163
transform -1 0 28428 0 1 40256
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1010__26
timestamp 1667941163
transform -1 0 27416 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1010_
timestamp 1667941163
transform 1 0 26496 0 1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1011__27
timestamp 1667941163
transform 1 0 28152 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1011_
timestamp 1667941163
transform -1 0 28428 0 1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1012__28
timestamp 1667941163
transform 1 0 17480 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1012_
timestamp 1667941163
transform 1 0 19136 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1013__29
timestamp 1667941163
transform -1 0 28152 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1013_
timestamp 1667941163
transform -1 0 26680 0 -1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1014__30
timestamp 1667941163
transform -1 0 3220 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1014_
timestamp 1667941163
transform 1 0 2944 0 -1 43520
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1015__31
timestamp 1667941163
transform -1 0 11960 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1015_
timestamp 1667941163
transform 1 0 11316 0 1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1016_
timestamp 1667941163
transform 1 0 1748 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1016__32
timestamp 1667941163
transform -1 0 2116 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1017__33
timestamp 1667941163
transform 1 0 26404 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1017_
timestamp 1667941163
transform 1 0 26496 0 1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1018__34
timestamp 1667941163
transform -1 0 28244 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1018_
timestamp 1667941163
transform -1 0 26680 0 -1 39168
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1019__35
timestamp 1667941163
transform -1 0 1932 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1019_
timestamp 1667941163
transform 1 0 1564 0 1 42432
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1020__36
timestamp 1667941163
transform -1 0 28152 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1020_
timestamp 1667941163
transform -1 0 26680 0 -1 31552
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1021_
timestamp 1667941163
transform 1 0 3036 0 -1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1021__37
timestamp 1667941163
transform -1 0 3312 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1022__38
timestamp 1667941163
transform 1 0 25852 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1022_
timestamp 1667941163
transform 1 0 26220 0 1 43520
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1023__39
timestamp 1667941163
transform -1 0 14536 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1023_
timestamp 1667941163
transform 1 0 14168 0 -1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1024__40
timestamp 1667941163
transform 1 0 9108 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1024_
timestamp 1667941163
transform 1 0 9200 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1025_
timestamp 1667941163
transform 1 0 26496 0 1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1025__41
timestamp 1667941163
transform -1 0 28060 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1026__42
timestamp 1667941163
transform -1 0 4232 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1026_
timestamp 1667941163
transform 1 0 3680 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1027__43
timestamp 1667941163
transform -1 0 28152 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1027_
timestamp 1667941163
transform 1 0 26496 0 1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1028__44
timestamp 1667941163
transform 1 0 2576 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1028_
timestamp 1667941163
transform -1 0 4048 0 -1 38080
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1029_
timestamp 1667941163
transform 1 0 26404 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1029__45
timestamp 1667941163
transform -1 0 27416 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1030__46
timestamp 1667941163
transform -1 0 4968 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1030_
timestamp 1667941163
transform 1 0 4140 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1031__47
timestamp 1667941163
transform -1 0 28152 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1031_
timestamp 1667941163
transform 1 0 26496 0 1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1032__48
timestamp 1667941163
transform -1 0 25484 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1032_
timestamp 1667941163
transform 1 0 24748 0 -1 44608
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1033_
timestamp 1667941163
transform 1 0 26496 0 1 38080
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1033__49
timestamp 1667941163
transform -1 0 27416 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1034__50
timestamp 1667941163
transform -1 0 17112 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1034_
timestamp 1667941163
transform 1 0 15916 0 1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1035_
timestamp 1667941163
transform 1 0 5244 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1035__51
timestamp 1667941163
transform 1 0 4600 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1036__52
timestamp 1667941163
transform -1 0 1932 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1036_
timestamp 1667941163
transform 1 0 1656 0 -1 34816
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1037__53
timestamp 1667941163
transform 1 0 27784 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1037_
timestamp 1667941163
transform -1 0 28428 0 1 33728
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1038__54
timestamp 1667941163
transform -1 0 8188 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1038_
timestamp 1667941163
transform 1 0 6992 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1039_
timestamp 1667941163
transform -1 0 26680 0 1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1039__55
timestamp 1667941163
transform 1 0 25668 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1040_
timestamp 1667941163
transform 1 0 1656 0 -1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1040__56
timestamp 1667941163
transform -1 0 1932 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1041__57
timestamp 1667941163
transform -1 0 14536 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1041_
timestamp 1667941163
transform 1 0 13984 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1042_
timestamp 1667941163
transform -1 0 11500 0 1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1043_
timestamp 1667941163
transform 1 0 26404 0 1 30464
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1044_
timestamp 1667941163
transform -1 0 10212 0 -1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1045_
timestamp 1667941163
transform -1 0 13616 0 -1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1046_
timestamp 1667941163
transform 1 0 26496 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1047_
timestamp 1667941163
transform 1 0 25852 0 1 36992
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1048_
timestamp 1667941163
transform 1 0 12696 0 -1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1049_
timestamp 1667941163
transform 1 0 25760 0 1 31552
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1050_
timestamp 1667941163
transform 1 0 3956 0 1 36992
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1051_
timestamp 1667941163
transform 1 0 25576 0 1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1052_
timestamp 1667941163
transform -1 0 22356 0 1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1053_
timestamp 1667941163
transform 1 0 19412 0 1 43520
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1054_
timestamp 1667941163
transform -1 0 16192 0 -1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1055_
timestamp 1667941163
transform 1 0 24564 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1056_
timestamp 1667941163
transform 1 0 26496 0 1 29376
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1057_
timestamp 1667941163
transform -1 0 24012 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1058_
timestamp 1667941163
transform 1 0 21988 0 -1 39168
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1059__58
timestamp 1667941163
transform -1 0 3312 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1059_
timestamp 1667941163
transform 1 0 2944 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1060__59
timestamp 1667941163
transform -1 0 20792 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1060_
timestamp 1667941163
transform 1 0 20240 0 1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1061_
timestamp 1667941163
transform 1 0 12788 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1061__60
timestamp 1667941163
transform -1 0 13156 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1062__61
timestamp 1667941163
transform -1 0 27416 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1062_
timestamp 1667941163
transform 1 0 26496 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1063_
timestamp 1667941163
transform 1 0 1564 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1063__62
timestamp 1667941163
transform -1 0 1932 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1064_
timestamp 1667941163
transform 1 0 1656 0 -1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1064__63
timestamp 1667941163
transform -1 0 1932 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1065__64
timestamp 1667941163
transform 1 0 1932 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1065_
timestamp 1667941163
transform -1 0 3496 0 1 36992
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1066__65
timestamp 1667941163
transform 1 0 28060 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1066_
timestamp 1667941163
transform -1 0 28428 0 1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1067__66
timestamp 1667941163
transform -1 0 27416 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1067_
timestamp 1667941163
transform 1 0 26496 0 1 42432
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1068__67
timestamp 1667941163
transform -1 0 27600 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1068_
timestamp 1667941163
transform 1 0 26496 0 1 39168
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1069_
timestamp 1667941163
transform 1 0 3956 0 1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1069__68
timestamp 1667941163
transform 1 0 3128 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1070__69
timestamp 1667941163
transform 1 0 27692 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1070_
timestamp 1667941163
transform -1 0 28428 0 1 44608
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1071__70
timestamp 1667941163
transform -1 0 20700 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1071_
timestamp 1667941163
transform 1 0 20332 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1072__71
timestamp 1667941163
transform 1 0 25852 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1072_
timestamp 1667941163
transform 1 0 26496 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1073__72
timestamp 1667941163
transform -1 0 23184 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1073_
timestamp 1667941163
transform 1 0 22816 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1074__73
timestamp 1667941163
transform -1 0 19688 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1074_
timestamp 1667941163
transform 1 0 19412 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1075_
timestamp 1667941163
transform -1 0 28428 0 1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1075__74
timestamp 1667941163
transform 1 0 27876 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1076_
timestamp 1667941163
transform 1 0 1656 0 -1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1076__75
timestamp 1667941163
transform -1 0 1932 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1077__76
timestamp 1667941163
transform -1 0 28152 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1077_
timestamp 1667941163
transform 1 0 26496 0 1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1078_
timestamp 1667941163
transform -1 0 3496 0 1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1078__77
timestamp 1667941163
transform 1 0 2300 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1079__78
timestamp 1667941163
transform 1 0 3220 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1079_
timestamp 1667941163
transform 1 0 3956 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1080__79
timestamp 1667941163
transform -1 0 8004 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1080_
timestamp 1667941163
transform 1 0 6900 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1081__80
timestamp 1667941163
transform 1 0 2300 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1081_
timestamp 1667941163
transform -1 0 3496 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1082_
timestamp 1667941163
transform -1 0 28428 0 1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1082__81
timestamp 1667941163
transform 1 0 27232 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1083__82
timestamp 1667941163
transform 1 0 27876 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1083_
timestamp 1667941163
transform -1 0 28428 0 1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1084_
timestamp 1667941163
transform 1 0 26496 0 1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1084__83
timestamp 1667941163
transform -1 0 28152 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1085_
timestamp 1667941163
transform 1 0 1564 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1085__84
timestamp 1667941163
transform -1 0 1932 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1086__85
timestamp 1667941163
transform -1 0 1932 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1086_
timestamp 1667941163
transform 1 0 1656 0 -1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1087__86
timestamp 1667941163
transform -1 0 28152 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1087_
timestamp 1667941163
transform 1 0 26496 0 1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1088__87
timestamp 1667941163
transform 1 0 9752 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1088_
timestamp 1667941163
transform 1 0 10396 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1089__88
timestamp 1667941163
transform -1 0 18584 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1089_
timestamp 1667941163
transform 1 0 18216 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1090__89
timestamp 1667941163
transform 1 0 2024 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1090_
timestamp 1667941163
transform 1 0 2300 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1091__90
timestamp 1667941163
transform 1 0 27876 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1091_
timestamp 1667941163
transform -1 0 28428 0 1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1092__91
timestamp 1667941163
transform 1 0 3128 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1092_
timestamp 1667941163
transform -1 0 3496 0 1 41344
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1093__92
timestamp 1667941163
transform -1 0 4232 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1093_
timestamp 1667941163
transform 1 0 3956 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1094_
timestamp 1667941163
transform 1 0 9292 0 1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1094__93
timestamp 1667941163
transform -1 0 9936 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1095_
timestamp 1667941163
transform 1 0 9292 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1095__94
timestamp 1667941163
transform -1 0 10672 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1096__95
timestamp 1667941163
transform 1 0 26404 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1096_
timestamp 1667941163
transform -1 0 26680 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1097__96
timestamp 1667941163
transform 1 0 27876 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1097_
timestamp 1667941163
transform -1 0 28428 0 1 41344
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1098__97
timestamp 1667941163
transform -1 0 13248 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1098_
timestamp 1667941163
transform 1 0 12880 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1099_
timestamp 1667941163
transform -1 0 28428 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1099__98
timestamp 1667941163
transform 1 0 27876 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1100__99
timestamp 1667941163
transform -1 0 28152 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1100_
timestamp 1667941163
transform 1 0 26496 0 1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1101__100
timestamp 1667941163
transform -1 0 1932 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1101_
timestamp 1667941163
transform 1 0 1656 0 -1 41344
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1102__101
timestamp 1667941163
transform -1 0 28152 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1102_
timestamp 1667941163
transform -1 0 26680 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1103_
timestamp 1667941163
transform 1 0 1564 0 1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1103__102
timestamp 1667941163
transform -1 0 1932 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1104__103
timestamp 1667941163
transform 1 0 27876 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1104_
timestamp 1667941163
transform -1 0 28428 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1105__104
timestamp 1667941163
transform -1 0 2668 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1105_
timestamp 1667941163
transform 1 0 1656 0 -1 40256
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1106__105
timestamp 1667941163
transform -1 0 1932 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1106_
timestamp 1667941163
transform 1 0 1564 0 1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1107__106
timestamp 1667941163
transform -1 0 1932 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1107_
timestamp 1667941163
transform 1 0 1564 0 1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1108_
timestamp 1667941163
transform 1 0 1564 0 1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1108__107
timestamp 1667941163
transform -1 0 1932 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_wb_clk_i $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 24104 0 1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_0__f_wb_clk_i
timestamp 1667941163
transform -1 0 20056 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_1__f_wb_clk_i
timestamp 1667941163
transform 1 0 23368 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_2__f_wb_clk_i
timestamp 1667941163
transform -1 0 20056 0 -1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_3__f_wb_clk_i
timestamp 1667941163
transform 1 0 20792 0 1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 27876 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 1667941163
transform -1 0 25852 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1667941163
transform -1 0 1840 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1667941163
transform 1 0 28152 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1667941163
transform 1 0 27140 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1667941163
transform 1 0 17572 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1667941163
transform 1 0 28152 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input6 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 1564 0 -1 30464
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1667941163
transform 1 0 26404 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input8
timestamp 1667941163
transform -1 0 17204 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input9
timestamp 1667941163
transform 1 0 9108 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1667941163
transform -1 0 1840 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1667941163
transform 1 0 23828 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1667941163
transform 1 0 28152 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1667941163
transform -1 0 6072 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1667941163
transform -1 0 1840 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input15
timestamp 1667941163
transform -1 0 6808 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input16
timestamp 1667941163
transform -1 0 1840 0 -1 28288
box -38 -48 314 592
<< labels >>
flabel metal3 s 200 36668 800 36908 0 FreeSans 960 0 0 0 active
port 0 nsew signal input
flabel metal2 s 12226 200 12338 800 0 FreeSans 448 90 0 0 io_in[0]
port 1 nsew signal input
flabel metal2 s 12226 49200 12338 49800 0 FreeSans 448 90 0 0 io_in[10]
port 2 nsew signal input
flabel metal3 s 200 40068 800 40308 0 FreeSans 960 0 0 0 io_in[11]
port 3 nsew signal input
flabel metal3 s 29200 43468 29800 43708 0 FreeSans 960 0 0 0 io_in[12]
port 4 nsew signal input
flabel metal2 s 18666 200 18778 800 0 FreeSans 448 90 0 0 io_in[13]
port 5 nsew signal input
flabel metal2 s 5142 49200 5254 49800 0 FreeSans 448 90 0 0 io_in[14]
port 6 nsew signal input
flabel metal3 s 29200 45508 29800 45748 0 FreeSans 960 0 0 0 io_in[15]
port 7 nsew signal input
flabel metal3 s 29200 13548 29800 13788 0 FreeSans 960 0 0 0 io_in[16]
port 8 nsew signal input
flabel metal3 s 200 48228 800 48468 0 FreeSans 960 0 0 0 io_in[17]
port 9 nsew signal input
flabel metal2 s -10 49200 102 49800 0 FreeSans 448 90 0 0 io_in[18]
port 10 nsew signal input
flabel metal3 s 29200 4028 29800 4268 0 FreeSans 960 0 0 0 io_in[19]
port 11 nsew signal input
flabel metal3 s 200 12868 800 13108 0 FreeSans 960 0 0 0 io_in[1]
port 12 nsew signal input
flabel metal3 s 200 23068 800 23308 0 FreeSans 960 0 0 0 io_in[20]
port 13 nsew signal input
flabel metal3 s 200 14908 800 15148 0 FreeSans 960 0 0 0 io_in[21]
port 14 nsew signal input
flabel metal3 s 29200 23068 29800 23308 0 FreeSans 960 0 0 0 io_in[22]
port 15 nsew signal input
flabel metal3 s 200 47548 800 47788 0 FreeSans 960 0 0 0 io_in[23]
port 16 nsew signal input
flabel metal3 s 200 45508 800 45748 0 FreeSans 960 0 0 0 io_in[24]
port 17 nsew signal input
flabel metal2 s 29614 200 29726 800 0 FreeSans 448 90 0 0 io_in[25]
port 18 nsew signal input
flabel metal2 s 28970 200 29082 800 0 FreeSans 448 90 0 0 io_in[26]
port 19 nsew signal input
flabel metal3 s 29200 18988 29800 19228 0 FreeSans 960 0 0 0 io_in[27]
port 20 nsew signal input
flabel metal2 s 26394 200 26506 800 0 FreeSans 448 90 0 0 io_in[28]
port 21 nsew signal input
flabel metal2 s 29614 49200 29726 49800 0 FreeSans 448 90 0 0 io_in[29]
port 22 nsew signal input
flabel metal2 s 12870 200 12982 800 0 FreeSans 448 90 0 0 io_in[2]
port 23 nsew signal input
flabel metal3 s 29200 25788 29800 26028 0 FreeSans 960 0 0 0 io_in[30]
port 24 nsew signal input
flabel metal3 s 200 35308 800 35548 0 FreeSans 960 0 0 0 io_in[31]
port 25 nsew signal input
flabel metal2 s 24462 200 24574 800 0 FreeSans 448 90 0 0 io_in[32]
port 26 nsew signal input
flabel metal3 s 200 20348 800 20588 0 FreeSans 960 0 0 0 io_in[33]
port 27 nsew signal input
flabel metal2 s 20598 49200 20710 49800 0 FreeSans 448 90 0 0 io_in[34]
port 28 nsew signal input
flabel metal2 s 25106 49200 25218 49800 0 FreeSans 448 90 0 0 io_in[35]
port 29 nsew signal input
flabel metal3 s 29200 35308 29800 35548 0 FreeSans 960 0 0 0 io_in[36]
port 30 nsew signal input
flabel metal2 s 25750 49200 25862 49800 0 FreeSans 448 90 0 0 io_in[37]
port 31 nsew signal input
flabel metal2 s 12870 49200 12982 49800 0 FreeSans 448 90 0 0 io_in[3]
port 32 nsew signal input
flabel metal3 s 29200 34628 29800 34868 0 FreeSans 960 0 0 0 io_in[4]
port 33 nsew signal input
flabel metal3 s 29200 48228 29800 48468 0 FreeSans 960 0 0 0 io_in[5]
port 34 nsew signal input
flabel metal3 s 200 24428 800 24668 0 FreeSans 960 0 0 0 io_in[6]
port 35 nsew signal input
flabel metal3 s 200 16948 800 17188 0 FreeSans 960 0 0 0 io_in[7]
port 36 nsew signal input
flabel metal3 s 29200 36668 29800 36908 0 FreeSans 960 0 0 0 io_in[8]
port 37 nsew signal input
flabel metal3 s 200 46868 800 47108 0 FreeSans 960 0 0 0 io_in[9]
port 38 nsew signal input
flabel metal2 s 21242 200 21354 800 0 FreeSans 448 90 0 0 io_oeb[0]
port 39 nsew signal tristate
flabel metal3 s 200 13548 800 13788 0 FreeSans 960 0 0 0 io_oeb[10]
port 40 nsew signal tristate
flabel metal3 s 29200 32588 29800 32828 0 FreeSans 960 0 0 0 io_oeb[11]
port 41 nsew signal tristate
flabel metal3 s 29200 21708 29800 21948 0 FreeSans 960 0 0 0 io_oeb[12]
port 42 nsew signal tristate
flabel metal3 s 29200 21028 29800 21268 0 FreeSans 960 0 0 0 io_oeb[13]
port 43 nsew signal tristate
flabel metal3 s 200 3348 800 3588 0 FreeSans 960 0 0 0 io_oeb[14]
port 44 nsew signal tristate
flabel metal2 s 1278 49200 1390 49800 0 FreeSans 448 90 0 0 io_oeb[15]
port 45 nsew signal tristate
flabel metal3 s 29200 12188 29800 12428 0 FreeSans 960 0 0 0 io_oeb[16]
port 46 nsew signal tristate
flabel metal2 s 10938 200 11050 800 0 FreeSans 448 90 0 0 io_oeb[17]
port 47 nsew signal tristate
flabel metal2 s 18666 49200 18778 49800 0 FreeSans 448 90 0 0 io_oeb[18]
port 48 nsew signal tristate
flabel metal2 s 1922 49200 2034 49800 0 FreeSans 448 90 0 0 io_oeb[19]
port 49 nsew signal tristate
flabel metal3 s 29200 1308 29800 1548 0 FreeSans 960 0 0 0 io_oeb[1]
port 50 nsew signal tristate
flabel metal3 s 29200 27148 29800 27388 0 FreeSans 960 0 0 0 io_oeb[20]
port 51 nsew signal tristate
flabel metal3 s 200 41428 800 41668 0 FreeSans 960 0 0 0 io_oeb[21]
port 52 nsew signal tristate
flabel metal2 s 3854 200 3966 800 0 FreeSans 448 90 0 0 io_oeb[22]
port 53 nsew signal tristate
flabel metal2 s 10294 49200 10406 49800 0 FreeSans 448 90 0 0 io_oeb[23]
port 54 nsew signal tristate
flabel metal2 s 10938 49200 11050 49800 0 FreeSans 448 90 0 0 io_oeb[24]
port 55 nsew signal tristate
flabel metal3 s 29200 8108 29800 8348 0 FreeSans 960 0 0 0 io_oeb[25]
port 56 nsew signal tristate
flabel metal3 s 29200 41428 29800 41668 0 FreeSans 960 0 0 0 io_oeb[26]
port 57 nsew signal tristate
flabel metal2 s 13514 49200 13626 49800 0 FreeSans 448 90 0 0 io_oeb[27]
port 58 nsew signal tristate
flabel metal3 s 29200 3348 29800 3588 0 FreeSans 960 0 0 0 io_oeb[28]
port 59 nsew signal tristate
flabel metal3 s 29200 35988 29800 36228 0 FreeSans 960 0 0 0 io_oeb[29]
port 60 nsew signal tristate
flabel metal2 s 23174 49200 23286 49800 0 FreeSans 448 90 0 0 io_oeb[2]
port 61 nsew signal tristate
flabel metal3 s 200 42108 800 42348 0 FreeSans 960 0 0 0 io_oeb[30]
port 62 nsew signal tristate
flabel metal3 s 29200 2668 29800 2908 0 FreeSans 960 0 0 0 io_oeb[31]
port 63 nsew signal tristate
flabel metal3 s 200 19668 800 19908 0 FreeSans 960 0 0 0 io_oeb[32]
port 64 nsew signal tristate
flabel metal3 s 29200 8788 29800 9028 0 FreeSans 960 0 0 0 io_oeb[33]
port 65 nsew signal tristate
flabel metal3 s 200 49588 800 49828 0 FreeSans 960 0 0 0 io_oeb[34]
port 66 nsew signal tristate
flabel metal3 s 200 17628 800 17868 0 FreeSans 960 0 0 0 io_oeb[35]
port 67 nsew signal tristate
flabel metal3 s 200 8788 800 9028 0 FreeSans 960 0 0 0 io_oeb[36]
port 68 nsew signal tristate
flabel metal3 s 200 14228 800 14468 0 FreeSans 960 0 0 0 io_oeb[37]
port 69 nsew signal tristate
flabel metal2 s 19954 200 20066 800 0 FreeSans 448 90 0 0 io_oeb[3]
port 70 nsew signal tristate
flabel metal3 s 29200 10148 29800 10388 0 FreeSans 960 0 0 0 io_oeb[4]
port 71 nsew signal tristate
flabel metal3 s 200 25788 800 26028 0 FreeSans 960 0 0 0 io_oeb[5]
port 72 nsew signal tristate
flabel metal3 s 29200 24428 29800 24668 0 FreeSans 960 0 0 0 io_oeb[6]
port 73 nsew signal tristate
flabel metal2 s 634 49200 746 49800 0 FreeSans 448 90 0 0 io_oeb[7]
port 74 nsew signal tristate
flabel metal2 s 3210 200 3322 800 0 FreeSans 448 90 0 0 io_oeb[8]
port 75 nsew signal tristate
flabel metal2 s 8362 200 8474 800 0 FreeSans 448 90 0 0 io_oeb[9]
port 76 nsew signal tristate
flabel metal3 s 29200 47548 29800 47788 0 FreeSans 960 0 0 0 io_out[0]
port 77 nsew signal tristate
flabel metal3 s 29200 31908 29800 32148 0 FreeSans 960 0 0 0 io_out[10]
port 78 nsew signal tristate
flabel metal3 s 200 1988 800 2228 0 FreeSans 960 0 0 0 io_out[11]
port 79 nsew signal tristate
flabel metal3 s 200 6068 800 6308 0 FreeSans 960 0 0 0 io_out[12]
port 80 nsew signal tristate
flabel metal3 s 29200 1988 29800 2228 0 FreeSans 960 0 0 0 io_out[13]
port 81 nsew signal tristate
flabel metal3 s 29200 42108 29800 42348 0 FreeSans 960 0 0 0 io_out[14]
port 82 nsew signal tristate
flabel metal3 s 200 33268 800 33508 0 FreeSans 960 0 0 0 io_out[15]
port 83 nsew signal tristate
flabel metal3 s 29200 31228 29800 31468 0 FreeSans 960 0 0 0 io_out[16]
port 84 nsew signal tristate
flabel metal2 s 27038 49200 27150 49800 0 FreeSans 448 90 0 0 io_out[17]
port 85 nsew signal tristate
flabel metal3 s 29200 7428 29800 7668 0 FreeSans 960 0 0 0 io_out[18]
port 86 nsew signal tristate
flabel metal3 s 200 18988 800 19228 0 FreeSans 960 0 0 0 io_out[19]
port 87 nsew signal tristate
flabel metal2 s 16734 49200 16846 49800 0 FreeSans 448 90 0 0 io_out[1]
port 88 nsew signal tristate
flabel metal2 s 22530 49200 22642 49800 0 FreeSans 448 90 0 0 io_out[20]
port 89 nsew signal tristate
flabel metal3 s 200 31908 800 32148 0 FreeSans 960 0 0 0 io_out[21]
port 90 nsew signal tristate
flabel metal2 s 25106 200 25218 800 0 FreeSans 448 90 0 0 io_out[22]
port 91 nsew signal tristate
flabel metal3 s 29200 28508 29800 28748 0 FreeSans 960 0 0 0 io_out[23]
port 92 nsew signal tristate
flabel metal2 s 21886 200 21998 800 0 FreeSans 448 90 0 0 io_out[24]
port 93 nsew signal tristate
flabel metal2 s 19954 49200 20066 49800 0 FreeSans 448 90 0 0 io_out[25]
port 94 nsew signal tristate
flabel metal3 s 200 4028 800 4268 0 FreeSans 960 0 0 0 io_out[26]
port 95 nsew signal tristate
flabel metal2 s 21242 49200 21354 49800 0 FreeSans 448 90 0 0 io_out[27]
port 96 nsew signal tristate
flabel metal2 s 13514 200 13626 800 0 FreeSans 448 90 0 0 io_out[28]
port 97 nsew signal tristate
flabel metal3 s 29200 10828 29800 11068 0 FreeSans 960 0 0 0 io_out[29]
port 98 nsew signal tristate
flabel metal2 s 5786 200 5898 800 0 FreeSans 448 90 0 0 io_out[2]
port 99 nsew signal tristate
flabel metal3 s 200 4708 800 4948 0 FreeSans 960 0 0 0 io_out[30]
port 100 nsew signal tristate
flabel metal3 s 200 11508 800 11748 0 FreeSans 960 0 0 0 io_out[31]
port 101 nsew signal tristate
flabel metal3 s 200 37348 800 37588 0 FreeSans 960 0 0 0 io_out[32]
port 102 nsew signal tristate
flabel metal3 s 29200 15588 29800 15828 0 FreeSans 960 0 0 0 io_out[33]
port 103 nsew signal tristate
flabel metal3 s 29200 42788 29800 43028 0 FreeSans 960 0 0 0 io_out[34]
port 104 nsew signal tristate
flabel metal3 s 29200 40748 29800 40988 0 FreeSans 960 0 0 0 io_out[35]
port 105 nsew signal tristate
flabel metal2 s 2566 49200 2678 49800 0 FreeSans 448 90 0 0 io_out[36]
port 106 nsew signal tristate
flabel metal3 s 29200 46188 29800 46428 0 FreeSans 960 0 0 0 io_out[37]
port 107 nsew signal tristate
flabel metal3 s 200 34628 800 34868 0 FreeSans 960 0 0 0 io_out[3]
port 108 nsew signal tristate
flabel metal3 s 29200 33948 29800 34188 0 FreeSans 960 0 0 0 io_out[4]
port 109 nsew signal tristate
flabel metal2 s 8362 49200 8474 49800 0 FreeSans 448 90 0 0 io_out[5]
port 110 nsew signal tristate
flabel metal2 s 28326 49200 28438 49800 0 FreeSans 448 90 0 0 io_out[6]
port 111 nsew signal tristate
flabel metal3 s 200 15588 800 15828 0 FreeSans 960 0 0 0 io_out[7]
port 112 nsew signal tristate
flabel metal2 s 14802 200 14914 800 0 FreeSans 448 90 0 0 io_out[8]
port 113 nsew signal tristate
flabel metal3 s 200 12188 800 12428 0 FreeSans 960 0 0 0 io_out[9]
port 114 nsew signal tristate
flabel metal3 s 29200 16268 29800 16508 0 FreeSans 960 0 0 0 la1_data_in[0]
port 115 nsew signal input
flabel metal2 s 17378 200 17490 800 0 FreeSans 448 90 0 0 la1_data_in[10]
port 116 nsew signal input
flabel metal3 s 29200 14908 29800 15148 0 FreeSans 960 0 0 0 la1_data_in[11]
port 117 nsew signal input
flabel metal3 s 200 29868 800 30108 0 FreeSans 960 0 0 0 la1_data_in[12]
port 118 nsew signal input
flabel metal2 s 27038 200 27150 800 0 FreeSans 448 90 0 0 la1_data_in[13]
port 119 nsew signal input
flabel metal3 s 200 10148 800 10388 0 FreeSans 960 0 0 0 la1_data_in[14]
port 120 nsew signal input
flabel metal2 s 3210 49200 3322 49800 0 FreeSans 448 90 0 0 la1_data_in[15]
port 121 nsew signal input
flabel metal2 s 15446 49200 15558 49800 0 FreeSans 448 90 0 0 la1_data_in[16]
port 122 nsew signal input
flabel metal2 s 9650 49200 9762 49800 0 FreeSans 448 90 0 0 la1_data_in[17]
port 123 nsew signal input
flabel metal3 s 29200 4708 29800 4948 0 FreeSans 960 0 0 0 la1_data_in[18]
port 124 nsew signal input
flabel metal2 s 4498 49200 4610 49800 0 FreeSans 448 90 0 0 la1_data_in[19]
port 125 nsew signal input
flabel metal2 s 16090 200 16202 800 0 FreeSans 448 90 0 0 la1_data_in[1]
port 126 nsew signal input
flabel metal3 s 200 29188 800 29428 0 FreeSans 960 0 0 0 la1_data_in[20]
port 127 nsew signal input
flabel metal2 s 28970 49200 29082 49800 0 FreeSans 448 90 0 0 la1_data_in[21]
port 128 nsew signal input
flabel metal3 s 29200 17628 29800 17868 0 FreeSans 960 0 0 0 la1_data_in[22]
port 129 nsew signal input
flabel metal3 s 200 628 800 868 0 FreeSans 960 0 0 0 la1_data_in[23]
port 130 nsew signal input
flabel metal2 s 11582 200 11694 800 0 FreeSans 448 90 0 0 la1_data_in[24]
port 131 nsew signal input
flabel metal3 s 200 30548 800 30788 0 FreeSans 960 0 0 0 la1_data_in[25]
port 132 nsew signal input
flabel metal3 s 29200 12868 29800 13108 0 FreeSans 960 0 0 0 la1_data_in[26]
port 133 nsew signal input
flabel metal2 s 23174 200 23286 800 0 FreeSans 448 90 0 0 la1_data_in[27]
port 134 nsew signal input
flabel metal3 s 200 26468 800 26708 0 FreeSans 960 0 0 0 la1_data_in[28]
port 135 nsew signal input
flabel metal3 s 200 40748 800 40988 0 FreeSans 960 0 0 0 la1_data_in[29]
port 136 nsew signal input
flabel metal2 s 9006 200 9118 800 0 FreeSans 448 90 0 0 la1_data_in[2]
port 137 nsew signal input
flabel metal2 s 1278 200 1390 800 0 FreeSans 448 90 0 0 la1_data_in[30]
port 138 nsew signal input
flabel metal3 s 29200 -52 29800 188 0 FreeSans 960 0 0 0 la1_data_in[31]
port 139 nsew signal input
flabel metal3 s 200 25108 800 25348 0 FreeSans 960 0 0 0 la1_data_in[3]
port 140 nsew signal input
flabel metal2 s 23818 49200 23930 49800 0 FreeSans 448 90 0 0 la1_data_in[4]
port 141 nsew signal input
flabel metal3 s 29200 29868 29800 30108 0 FreeSans 960 0 0 0 la1_data_in[5]
port 142 nsew signal input
flabel metal2 s 5786 49200 5898 49800 0 FreeSans 448 90 0 0 la1_data_in[6]
port 143 nsew signal input
flabel metal3 s 200 18308 800 18548 0 FreeSans 960 0 0 0 la1_data_in[7]
port 144 nsew signal input
flabel metal2 s 6430 49200 6542 49800 0 FreeSans 448 90 0 0 la1_data_in[8]
port 145 nsew signal input
flabel metal3 s 200 27828 800 28068 0 FreeSans 960 0 0 0 la1_data_in[9]
port 146 nsew signal input
flabel metal2 s 6430 200 6542 800 0 FreeSans 448 90 0 0 la1_data_out[0]
port 147 nsew signal tristate
flabel metal3 s 29200 19668 29800 19908 0 FreeSans 960 0 0 0 la1_data_out[10]
port 148 nsew signal tristate
flabel metal2 s 18022 200 18134 800 0 FreeSans 448 90 0 0 la1_data_out[11]
port 149 nsew signal tristate
flabel metal3 s 29200 46868 29800 47108 0 FreeSans 960 0 0 0 la1_data_out[12]
port 150 nsew signal tristate
flabel metal3 s 200 44148 800 44388 0 FreeSans 960 0 0 0 la1_data_out[13]
port 151 nsew signal tristate
flabel metal2 s 11582 49200 11694 49800 0 FreeSans 448 90 0 0 la1_data_out[14]
port 152 nsew signal tristate
flabel metal3 s 200 1308 800 1548 0 FreeSans 960 0 0 0 la1_data_out[15]
port 153 nsew signal tristate
flabel metal3 s 29200 23748 29800 23988 0 FreeSans 960 0 0 0 la1_data_out[16]
port 154 nsew signal tristate
flabel metal3 s 29200 39388 29800 39628 0 FreeSans 960 0 0 0 la1_data_out[17]
port 155 nsew signal tristate
flabel metal3 s 200 44828 800 45068 0 FreeSans 960 0 0 0 la1_data_out[18]
port 156 nsew signal tristate
flabel metal3 s 29200 30548 29800 30788 0 FreeSans 960 0 0 0 la1_data_out[19]
port 157 nsew signal tristate
flabel metal3 s 200 35988 800 36228 0 FreeSans 960 0 0 0 la1_data_out[1]
port 158 nsew signal tristate
flabel metal3 s 200 8108 800 8348 0 FreeSans 960 0 0 0 la1_data_out[20]
port 159 nsew signal tristate
flabel metal3 s 29200 44828 29800 45068 0 FreeSans 960 0 0 0 la1_data_out[21]
port 160 nsew signal tristate
flabel metal2 s 14802 49200 14914 49800 0 FreeSans 448 90 0 0 la1_data_out[22]
port 161 nsew signal tristate
flabel metal2 s 9650 200 9762 800 0 FreeSans 448 90 0 0 la1_data_out[23]
port 162 nsew signal tristate
flabel metal3 s 29200 25108 29800 25348 0 FreeSans 960 0 0 0 la1_data_out[24]
port 163 nsew signal tristate
flabel metal3 s 200 2668 800 2908 0 FreeSans 960 0 0 0 la1_data_out[25]
port 164 nsew signal tristate
flabel metal3 s 29200 14228 29800 14468 0 FreeSans 960 0 0 0 la1_data_out[26]
port 165 nsew signal tristate
flabel metal3 s 200 38708 800 38948 0 FreeSans 960 0 0 0 la1_data_out[27]
port 166 nsew signal tristate
flabel metal3 s 29200 5388 29800 5628 0 FreeSans 960 0 0 0 la1_data_out[28]
port 167 nsew signal tristate
flabel metal2 s 4498 200 4610 800 0 FreeSans 448 90 0 0 la1_data_out[29]
port 168 nsew signal tristate
flabel metal2 s 16734 200 16846 800 0 FreeSans 448 90 0 0 la1_data_out[2]
port 169 nsew signal tristate
flabel metal3 s 29200 20348 29800 20588 0 FreeSans 960 0 0 0 la1_data_out[30]
port 170 nsew signal tristate
flabel metal3 s 29200 48908 29800 49148 0 FreeSans 960 0 0 0 la1_data_out[31]
port 171 nsew signal tristate
flabel metal3 s 200 7428 800 7668 0 FreeSans 960 0 0 0 la1_data_out[3]
port 172 nsew signal tristate
flabel metal3 s 29200 6748 29800 6988 0 FreeSans 960 0 0 0 la1_data_out[4]
port 173 nsew signal tristate
flabel metal2 s 2566 200 2678 800 0 FreeSans 448 90 0 0 la1_data_out[5]
port 174 nsew signal tristate
flabel metal3 s 29200 26468 29800 26708 0 FreeSans 960 0 0 0 la1_data_out[6]
port 175 nsew signal tristate
flabel metal2 s 634 200 746 800 0 FreeSans 448 90 0 0 la1_data_out[7]
port 176 nsew signal tristate
flabel metal3 s 29200 40068 29800 40308 0 FreeSans 960 0 0 0 la1_data_out[8]
port 177 nsew signal tristate
flabel metal2 s 27682 49200 27794 49800 0 FreeSans 448 90 0 0 la1_data_out[9]
port 178 nsew signal tristate
flabel metal3 s 29200 9468 29800 9708 0 FreeSans 960 0 0 0 la1_oenb[0]
port 179 nsew signal input
flabel metal2 s 26394 49200 26506 49800 0 FreeSans 448 90 0 0 la1_oenb[10]
port 180 nsew signal input
flabel metal3 s 200 22388 800 22628 0 FreeSans 960 0 0 0 la1_oenb[11]
port 181 nsew signal input
flabel metal3 s 200 23748 800 23988 0 FreeSans 960 0 0 0 la1_oenb[12]
port 182 nsew signal input
flabel metal2 s 23818 200 23930 800 0 FreeSans 448 90 0 0 la1_oenb[13]
port 183 nsew signal input
flabel metal2 s -10 200 102 800 0 FreeSans 448 90 0 0 la1_oenb[14]
port 184 nsew signal input
flabel metal2 s 28326 200 28438 800 0 FreeSans 448 90 0 0 la1_oenb[15]
port 185 nsew signal input
flabel metal3 s 200 28508 800 28748 0 FreeSans 960 0 0 0 la1_oenb[16]
port 186 nsew signal input
flabel metal3 s 200 42788 800 43028 0 FreeSans 960 0 0 0 la1_oenb[17]
port 187 nsew signal input
flabel metal2 s 7718 49200 7830 49800 0 FreeSans 448 90 0 0 la1_oenb[18]
port 188 nsew signal input
flabel metal3 s 200 21028 800 21268 0 FreeSans 960 0 0 0 la1_oenb[19]
port 189 nsew signal input
flabel metal2 s 7074 200 7186 800 0 FreeSans 448 90 0 0 la1_oenb[1]
port 190 nsew signal input
flabel metal2 s 1922 200 2034 800 0 FreeSans 448 90 0 0 la1_oenb[20]
port 191 nsew signal input
flabel metal2 s 16090 49200 16202 49800 0 FreeSans 448 90 0 0 la1_oenb[21]
port 192 nsew signal input
flabel metal2 s 7074 49200 7186 49800 0 FreeSans 448 90 0 0 la1_oenb[22]
port 193 nsew signal input
flabel metal2 s 19310 200 19422 800 0 FreeSans 448 90 0 0 la1_oenb[23]
port 194 nsew signal input
flabel metal2 s 21886 49200 21998 49800 0 FreeSans 448 90 0 0 la1_oenb[24]
port 195 nsew signal input
flabel metal3 s 29200 18308 29800 18548 0 FreeSans 960 0 0 0 la1_oenb[25]
port 196 nsew signal input
flabel metal3 s 200 31228 800 31468 0 FreeSans 960 0 0 0 la1_oenb[26]
port 197 nsew signal input
flabel metal3 s 29200 38028 29800 38268 0 FreeSans 960 0 0 0 la1_oenb[27]
port 198 nsew signal input
flabel metal2 s 7718 200 7830 800 0 FreeSans 448 90 0 0 la1_oenb[28]
port 199 nsew signal input
flabel metal2 s 14158 200 14270 800 0 FreeSans 448 90 0 0 la1_oenb[29]
port 200 nsew signal input
flabel metal3 s 200 6748 800 6988 0 FreeSans 960 0 0 0 la1_oenb[2]
port 201 nsew signal input
flabel metal3 s 29200 37348 29800 37588 0 FreeSans 960 0 0 0 la1_oenb[30]
port 202 nsew signal input
flabel metal2 s 22530 200 22642 800 0 FreeSans 448 90 0 0 la1_oenb[31]
port 203 nsew signal input
flabel metal2 s 18022 49200 18134 49800 0 FreeSans 448 90 0 0 la1_oenb[3]
port 204 nsew signal input
flabel metal2 s 17378 49200 17490 49800 0 FreeSans 448 90 0 0 la1_oenb[4]
port 205 nsew signal input
flabel metal3 s 200 39388 800 39628 0 FreeSans 960 0 0 0 la1_oenb[5]
port 206 nsew signal input
flabel metal3 s 200 46188 800 46428 0 FreeSans 960 0 0 0 la1_oenb[6]
port 207 nsew signal input
flabel metal2 s 27682 200 27794 800 0 FreeSans 448 90 0 0 la1_oenb[7]
port 208 nsew signal input
flabel metal3 s 200 9468 800 9708 0 FreeSans 960 0 0 0 la1_oenb[8]
port 209 nsew signal input
flabel metal3 s 200 33948 800 34188 0 FreeSans 960 0 0 0 la1_oenb[9]
port 210 nsew signal input
flabel metal4 s 4417 2128 4737 47376 0 FreeSans 1920 90 0 0 vccd1
port 211 nsew power bidirectional
flabel metal4 s 11363 2128 11683 47376 0 FreeSans 1920 90 0 0 vccd1
port 211 nsew power bidirectional
flabel metal4 s 18309 2128 18629 47376 0 FreeSans 1920 90 0 0 vccd1
port 211 nsew power bidirectional
flabel metal4 s 25255 2128 25575 47376 0 FreeSans 1920 90 0 0 vccd1
port 211 nsew power bidirectional
flabel metal4 s 7890 2128 8210 47376 0 FreeSans 1920 90 0 0 vssd1
port 212 nsew ground bidirectional
flabel metal4 s 14836 2128 15156 47376 0 FreeSans 1920 90 0 0 vssd1
port 212 nsew ground bidirectional
flabel metal4 s 21782 2128 22102 47376 0 FreeSans 1920 90 0 0 vssd1
port 212 nsew ground bidirectional
flabel metal4 s 28728 2128 29048 47376 0 FreeSans 1920 90 0 0 vssd1
port 212 nsew ground bidirectional
flabel metal3 s 29200 29188 29800 29428 0 FreeSans 960 0 0 0 wb_clk_i
port 213 nsew signal input
rlabel metal1 14996 47328 14996 47328 0 vccd1
rlabel via1 15076 46784 15076 46784 0 vssd1
rlabel metal1 21344 33626 21344 33626 0 _0000_
rlabel via1 23050 16558 23050 16558 0 _0001_
rlabel metal1 19412 12954 19412 12954 0 _0002_
rlabel metal1 19688 12410 19688 12410 0 _0003_
rlabel via1 21569 14314 21569 14314 0 _0004_
rlabel metal2 20746 21794 20746 21794 0 _0005_
rlabel metal2 19734 23970 19734 23970 0 _0006_
rlabel via1 19545 20502 19545 20502 0 _0007_
rlabel metal2 19826 26962 19826 26962 0 _0008_
rlabel metal1 16728 25942 16728 25942 0 _0009_
rlabel metal1 17240 26962 17240 26962 0 _0010_
rlabel via1 22857 34646 22857 34646 0 _0011_
rlabel metal2 26266 35224 26266 35224 0 _0012_
rlabel via1 17153 35054 17153 35054 0 _0013_
rlabel metal1 17056 20434 17056 20434 0 _0014_
rlabel metal1 17208 33558 17208 33558 0 _0015_
rlabel metal2 17066 28322 17066 28322 0 _0016_
rlabel metal2 16330 14178 16330 14178 0 _0017_
rlabel metal2 28014 18530 28014 18530 0 _0018_
rlabel via1 17153 16558 17153 16558 0 _0019_
rlabel metal1 25146 16150 25146 16150 0 _0020_
rlabel metal1 23772 17170 23772 17170 0 _0021_
rlabel metal2 23230 27234 23230 27234 0 _0022_
rlabel via1 23234 19414 23234 19414 0 _0023_
rlabel metal2 22034 29784 22034 29784 0 _0024_
rlabel metal1 21063 26350 21063 26350 0 _0025_
rlabel via1 23142 20910 23142 20910 0 _0026_
rlabel metal2 22402 24786 22402 24786 0 _0027_
rlabel metal1 24732 14314 24732 14314 0 _0028_
rlabel metal2 24794 13430 24794 13430 0 _0029_
rlabel metal1 23372 14994 23372 14994 0 _0030_
rlabel metal1 21850 11866 21850 11866 0 _0031_
rlabel metal1 19632 29614 19632 29614 0 _0032_
rlabel metal1 19212 32470 19212 32470 0 _0033_
rlabel via1 22406 35054 22406 35054 0 _0034_
rlabel metal1 19632 35054 19632 35054 0 _0035_
rlabel metal1 18344 35666 18344 35666 0 _0036_
rlabel via1 17337 34578 17337 34578 0 _0037_
rlabel metal1 17622 29546 17622 29546 0 _0038_
rlabel metal1 18078 31858 18078 31858 0 _0039_
rlabel metal1 16636 21590 16636 21590 0 _0040_
rlabel metal1 17434 24378 17434 24378 0 _0041_
rlabel metal1 18768 25466 18768 25466 0 _0042_
rlabel via1 18533 13906 18533 13906 0 _0043_
rlabel metal2 25622 19992 25622 19992 0 _0044_
rlabel metal1 25208 22202 25208 22202 0 _0045_
rlabel metal1 26036 25466 26036 25466 0 _0046_
rlabel metal2 25806 27846 25806 27846 0 _0047_
rlabel via1 24881 17646 24881 17646 0 _0048_
rlabel metal1 21845 31790 21845 31790 0 _0049_
rlabel metal1 23460 33082 23460 33082 0 _0050_
rlabel metal2 4278 36448 4278 36448 0 _0051_
rlabel metal1 4370 3468 4370 3468 0 _0052_
rlabel metal1 2438 39440 2438 39440 0 _0053_
rlabel metal1 2806 42194 2806 42194 0 _0054_
rlabel metal1 2530 5236 2530 5236 0 _0055_
rlabel metal2 5198 44608 5198 44608 0 _0056_
rlabel metal1 5934 4114 5934 4114 0 _0057_
rlabel metal1 1978 4182 1978 4182 0 _0058_
rlabel metal1 2346 6222 2346 6222 0 _0059_
rlabel metal1 2392 11118 2392 11118 0 _0060_
rlabel metal1 4278 38318 4278 38318 0 _0061_
rlabel metal1 4876 36686 4876 36686 0 _0062_
rlabel metal1 17066 15028 17066 15028 0 _0063_
rlabel metal2 15594 14586 15594 14586 0 _0064_
rlabel metal1 12282 14416 12282 14416 0 _0065_
rlabel metal1 15870 14892 15870 14892 0 _0066_
rlabel metal1 13202 14348 13202 14348 0 _0067_
rlabel metal1 16054 14926 16054 14926 0 _0068_
rlabel metal1 13110 14926 13110 14926 0 _0069_
rlabel metal1 13800 15674 13800 15674 0 _0070_
rlabel metal1 13570 15130 13570 15130 0 _0071_
rlabel metal1 15732 15130 15732 15130 0 _0072_
rlabel metal2 15318 14756 15318 14756 0 _0073_
rlabel metal2 15502 14858 15502 14858 0 _0074_
rlabel metal1 14444 13498 14444 13498 0 _0075_
rlabel metal1 14858 13294 14858 13294 0 _0076_
rlabel metal2 15226 15470 15226 15470 0 _0077_
rlabel metal1 24564 37230 24564 37230 0 _0078_
rlabel metal2 13754 16388 13754 16388 0 _0079_
rlabel metal1 23552 36074 23552 36074 0 _0080_
rlabel metal1 21436 33490 21436 33490 0 _0081_
rlabel metal1 18400 19414 18400 19414 0 _0082_
rlabel metal1 21666 19890 21666 19890 0 _0083_
rlabel metal2 22218 16694 22218 16694 0 _0084_
rlabel metal1 22632 17170 22632 17170 0 _0085_
rlabel metal1 20332 11118 20332 11118 0 _0086_
rlabel metal2 19734 11322 19734 11322 0 _0087_
rlabel metal1 19596 11322 19596 11322 0 _0088_
rlabel metal1 20010 11730 20010 11730 0 _0089_
rlabel metal2 19458 12036 19458 12036 0 _0090_
rlabel metal2 20930 10812 20930 10812 0 _0091_
rlabel metal2 21114 11492 21114 11492 0 _0092_
rlabel metal2 20746 22916 20746 22916 0 _0093_
rlabel metal2 20930 22236 20930 22236 0 _0094_
rlabel metal2 20470 24310 20470 24310 0 _0095_
rlabel metal2 19918 24140 19918 24140 0 _0096_
rlabel metal1 19642 20944 19642 20944 0 _0097_
rlabel metal1 19090 20910 19090 20910 0 _0098_
rlabel metal1 20286 24922 20286 24922 0 _0099_
rlabel metal1 19918 26010 19918 26010 0 _0100_
rlabel metal1 16606 22066 16606 22066 0 _0101_
rlabel metal1 23506 37332 23506 37332 0 _0102_
rlabel metal1 16698 25160 16698 25160 0 _0103_
rlabel metal1 16606 25466 16606 25466 0 _0104_
rlabel metal1 16100 26554 16100 26554 0 _0105_
rlabel metal2 16330 27268 16330 27268 0 _0106_
rlabel metal2 22770 36618 22770 36618 0 _0107_
rlabel metal1 23092 36006 23092 36006 0 _0108_
rlabel metal1 27186 33592 27186 33592 0 _0109_
rlabel metal1 27416 33626 27416 33626 0 _0110_
rlabel metal2 15778 36108 15778 36108 0 _0111_
rlabel metal1 16422 35666 16422 35666 0 _0112_
rlabel metal2 15226 20230 15226 20230 0 _0113_
rlabel metal1 15962 20570 15962 20570 0 _0114_
rlabel metal1 15870 34578 15870 34578 0 _0115_
rlabel metal2 16054 34170 16054 34170 0 _0116_
rlabel metal1 15824 27642 15824 27642 0 _0117_
rlabel metal1 16836 28050 16836 28050 0 _0118_
rlabel metal2 16790 13498 16790 13498 0 _0119_
rlabel metal2 16606 13702 16606 13702 0 _0120_
rlabel metal1 27278 17306 27278 17306 0 _0121_
rlabel metal1 27876 18258 27876 18258 0 _0122_
rlabel metal1 15548 17850 15548 17850 0 _0123_
rlabel metal2 16882 17612 16882 17612 0 _0124_
rlabel metal1 25484 15674 25484 15674 0 _0125_
rlabel metal1 24748 16082 24748 16082 0 _0126_
rlabel metal1 19412 22406 19412 22406 0 _0127_
rlabel metal1 19274 17170 19274 17170 0 _0128_
rlabel metal1 18768 17646 18768 17646 0 _0129_
rlabel metal1 19458 17680 19458 17680 0 _0130_
rlabel metal1 21344 18394 21344 18394 0 _0131_
rlabel metal2 19642 18292 19642 18292 0 _0132_
rlabel metal1 15962 33490 15962 33490 0 _0133_
rlabel metal2 17526 40188 17526 40188 0 _0134_
rlabel metal2 15502 38182 15502 38182 0 _0135_
rlabel metal1 20470 34170 20470 34170 0 _0136_
rlabel metal1 20746 31824 20746 31824 0 _0137_
rlabel metal2 19458 34323 19458 34323 0 _0138_
rlabel metal1 20424 37230 20424 37230 0 _0139_
rlabel metal1 19734 36346 19734 36346 0 _0140_
rlabel metal1 20700 39270 20700 39270 0 _0141_
rlabel metal2 20102 37604 20102 37604 0 _0142_
rlabel metal1 18538 37910 18538 37910 0 _0143_
rlabel metal1 16422 33014 16422 33014 0 _0144_
rlabel metal1 16468 37774 16468 37774 0 _0145_
rlabel metal1 18538 38998 18538 38998 0 _0146_
rlabel metal2 17158 37808 17158 37808 0 _0147_
rlabel metal2 18446 38012 18446 38012 0 _0148_
rlabel metal1 19136 37434 19136 37434 0 _0149_
rlabel metal1 16652 37842 16652 37842 0 _0150_
rlabel metal1 17404 37162 17404 37162 0 _0151_
rlabel metal2 17342 37638 17342 37638 0 _0152_
rlabel metal2 16054 38012 16054 38012 0 _0153_
rlabel metal1 16675 37910 16675 37910 0 _0154_
rlabel metal1 16836 19482 16836 19482 0 _0155_
rlabel metal2 17526 18428 17526 18428 0 _0156_
rlabel metal1 18216 17306 18216 17306 0 _0157_
rlabel metal1 17296 17578 17296 17578 0 _0158_
rlabel metal2 17710 23324 17710 23324 0 _0159_
rlabel metal1 17204 18734 17204 18734 0 _0160_
rlabel metal2 17250 18496 17250 18496 0 _0161_
rlabel metal1 17158 18292 17158 18292 0 _0162_
rlabel metal2 16882 18870 16882 18870 0 _0163_
rlabel metal2 17434 18598 17434 18598 0 _0164_
rlabel metal1 18262 19346 18262 19346 0 _0165_
rlabel metal2 19734 19142 19734 19142 0 _0166_
rlabel metal1 19274 30158 19274 30158 0 _0167_
rlabel metal1 25622 21522 25622 21522 0 _0168_
rlabel metal1 27002 25942 27002 25942 0 _0169_
rlabel metal1 23690 30022 23690 30022 0 _0170_
rlabel metal1 21758 19788 21758 19788 0 _0171_
rlabel metal1 22908 17646 22908 17646 0 _0172_
rlabel metal1 22448 12818 22448 12818 0 _0173_
rlabel metal1 23368 18870 23368 18870 0 _0174_
rlabel metal1 23506 18598 23506 18598 0 _0175_
rlabel metal2 23874 17374 23874 17374 0 _0176_
rlabel metal2 22494 28322 22494 28322 0 _0177_
rlabel metal1 23966 33932 23966 33932 0 _0178_
rlabel metal2 23230 29716 23230 29716 0 _0179_
rlabel metal1 22494 29274 22494 29274 0 _0180_
rlabel metal2 22954 26520 22954 26520 0 _0181_
rlabel metal1 22080 26962 22080 26962 0 _0182_
rlabel metal1 22678 22406 22678 22406 0 _0183_
rlabel metal2 22954 21828 22954 21828 0 _0184_
rlabel metal2 21758 25466 21758 25466 0 _0185_
rlabel metal2 22862 25024 22862 25024 0 _0186_
rlabel metal1 25116 11866 25116 11866 0 _0187_
rlabel metal2 25162 11764 25162 11764 0 _0188_
rlabel metal1 25070 12750 25070 12750 0 _0189_
rlabel metal1 24288 11866 24288 11866 0 _0190_
rlabel metal1 23138 12274 23138 12274 0 _0191_
rlabel metal1 23138 12614 23138 12614 0 _0192_
rlabel metal2 23598 11526 23598 11526 0 _0193_
rlabel metal1 22264 11118 22264 11118 0 _0194_
rlabel metal2 22402 11594 22402 11594 0 _0195_
rlabel metal1 22540 11730 22540 11730 0 _0196_
rlabel metal1 20654 19244 20654 19244 0 _0197_
rlabel metal1 19596 30226 19596 30226 0 _0198_
rlabel metal1 16928 31790 16928 31790 0 _0199_
rlabel metal1 20746 32538 20746 32538 0 _0200_
rlabel metal1 20562 32946 20562 32946 0 _0201_
rlabel metal1 16376 31790 16376 31790 0 _0202_
rlabel metal2 18906 32572 18906 32572 0 _0203_
rlabel metal2 20838 36482 20838 36482 0 _0204_
rlabel metal1 19918 38896 19918 38896 0 _0205_
rlabel metal2 20838 37060 20838 37060 0 _0206_
rlabel metal1 19918 39066 19918 39066 0 _0207_
rlabel metal1 19366 39814 19366 39814 0 _0208_
rlabel metal2 19274 38012 19274 38012 0 _0209_
rlabel metal1 18630 39542 18630 39542 0 _0210_
rlabel metal1 18860 39066 18860 39066 0 _0211_
rlabel metal1 18216 39270 18216 39270 0 _0212_
rlabel metal2 17342 39746 17342 39746 0 _0213_
rlabel metal1 16882 39950 16882 39950 0 _0214_
rlabel metal1 17112 36142 17112 36142 0 _0215_
rlabel metal1 16744 30090 16744 30090 0 _0216_
rlabel metal1 17112 30566 17112 30566 0 _0217_
rlabel metal2 16882 29818 16882 29818 0 _0218_
rlabel metal2 16652 31892 16652 31892 0 _0219_
rlabel metal1 16284 31178 16284 31178 0 _0220_
rlabel metal1 17434 31824 17434 31824 0 _0221_
rlabel metal1 17158 22644 17158 22644 0 _0222_
rlabel metal1 17526 23018 17526 23018 0 _0223_
rlabel metal1 16560 21998 16560 21998 0 _0224_
rlabel metal1 17940 23222 17940 23222 0 _0225_
rlabel metal2 17618 23324 17618 23324 0 _0226_
rlabel metal1 17296 23290 17296 23290 0 _0227_
rlabel metal1 19918 19142 19918 19142 0 _0228_
rlabel metal2 18906 23052 18906 23052 0 _0229_
rlabel metal1 18400 22746 18400 22746 0 _0230_
rlabel metal1 19182 19176 19182 19176 0 _0231_
rlabel metal1 18413 19482 18413 19482 0 _0232_
rlabel metal1 18906 14416 18906 14416 0 _0233_
rlabel metal2 23690 29954 23690 29954 0 _0234_
rlabel metal1 25392 30906 25392 30906 0 _0235_
rlabel metal1 24794 21590 24794 21590 0 _0236_
rlabel metal1 25292 32742 25292 32742 0 _0237_
rlabel metal1 23782 32878 23782 32878 0 _0238_
rlabel metal1 23736 31450 23736 31450 0 _0239_
rlabel metal1 24564 30226 24564 30226 0 _0240_
rlabel metal1 23874 31926 23874 31926 0 _0241_
rlabel metal1 25254 21556 25254 21556 0 _0242_
rlabel metal2 25162 20332 25162 20332 0 _0243_
rlabel metal1 23782 22474 23782 22474 0 _0244_
rlabel metal1 23966 24038 23966 24038 0 _0245_
rlabel metal1 24288 21454 24288 21454 0 _0246_
rlabel metal1 23782 22406 23782 22406 0 _0247_
rlabel metal1 24794 22032 24794 22032 0 _0248_
rlabel metal1 25622 25772 25622 25772 0 _0249_
rlabel metal1 25346 24922 25346 24922 0 _0250_
rlabel metal1 24058 26962 24058 26962 0 _0251_
rlabel metal2 24058 28118 24058 28118 0 _0252_
rlabel metal2 24702 24378 24702 24378 0 _0253_
rlabel metal1 24886 24378 24886 24378 0 _0254_
rlabel metal2 25530 26044 25530 26044 0 _0255_
rlabel metal1 25392 26010 25392 26010 0 _0256_
rlabel metal2 24978 29920 24978 29920 0 _0257_
rlabel metal1 25346 27404 25346 27404 0 _0258_
rlabel metal2 24702 27778 24702 27778 0 _0259_
rlabel metal2 23414 30974 23414 30974 0 _0260_
rlabel metal2 24518 28220 24518 28220 0 _0261_
rlabel metal2 25990 29750 25990 29750 0 _0262_
rlabel metal1 24610 28084 24610 28084 0 _0263_
rlabel metal2 24794 23834 24794 23834 0 _0264_
rlabel metal2 23138 31110 23138 31110 0 _0265_
rlabel metal1 22770 30906 22770 30906 0 _0266_
rlabel metal2 23230 31552 23230 31552 0 _0267_
rlabel metal2 23690 32028 23690 32028 0 _0268_
rlabel metal1 22816 31654 22816 31654 0 _0269_
rlabel metal2 23598 33354 23598 33354 0 _0270_
rlabel metal2 5934 3740 5934 3740 0 _0271_
rlabel metal2 1794 36380 1794 36380 0 _0272_
rlabel metal2 17066 3230 17066 3230 0 _0273_
rlabel metal1 2024 8058 2024 8058 0 _0274_
rlabel metal1 27002 6358 27002 6358 0 _0275_
rlabel metal1 2852 4114 2852 4114 0 _0276_
rlabel metal2 27370 28322 27370 28322 0 _0277_
rlabel metal2 1794 3740 1794 3740 0 _0278_
rlabel metal2 28198 40732 28198 40732 0 _0279_
rlabel metal1 26358 45866 26358 45866 0 _0280_
rlabel metal1 28060 16762 28060 16762 0 _0281_
rlabel metal2 19366 3230 19366 3230 0 _0282_
rlabel metal1 26864 45526 26864 45526 0 _0283_
rlabel metal2 3174 43486 3174 43486 0 _0284_
rlabel metal1 11178 45866 11178 45866 0 _0285_
rlabel metal2 1978 3774 1978 3774 0 _0286_
rlabel metal2 27278 22882 27278 22882 0 _0287_
rlabel metal1 27140 38998 27140 38998 0 _0288_
rlabel metal2 1794 42908 1794 42908 0 _0289_
rlabel metal1 27140 31246 27140 31246 0 _0290_
rlabel metal2 4094 9316 4094 9316 0 _0291_
rlabel metal2 26450 43996 26450 43996 0 _0292_
rlabel metal1 14352 44506 14352 44506 0 _0293_
rlabel metal2 9430 5712 9430 5712 0 _0294_
rlabel metal1 27002 24922 27002 24922 0 _0295_
rlabel metal2 4278 3876 4278 3876 0 _0296_
rlabel metal2 26726 14620 26726 14620 0 _0297_
rlabel metal1 4186 37910 4186 37910 0 _0298_
rlabel metal1 26542 5338 26542 5338 0 _0299_
rlabel metal2 4370 3502 4370 3502 0 _0300_
rlabel metal2 26726 20536 26726 20536 0 _0301_
rlabel metal1 25024 44438 25024 44438 0 _0302_
rlabel metal1 27002 36890 27002 36890 0 _0303_
rlabel metal2 16146 46172 16146 46172 0 _0304_
rlabel metal2 5474 4828 5474 4828 0 _0305_
rlabel metal1 2024 34170 2024 34170 0 _0306_
rlabel metal2 28106 33762 28106 33762 0 _0307_
rlabel metal2 7958 46308 7958 46308 0 _0308_
rlabel metal2 26450 46818 26450 46818 0 _0309_
rlabel metal2 1886 16286 1886 16286 0 _0310_
rlabel metal2 14214 3230 14214 3230 0 _0311_
rlabel metal1 10534 13498 10534 13498 0 _0312_
rlabel metal1 26956 30362 26956 30362 0 _0313_
rlabel metal2 9982 14110 9982 14110 0 _0314_
rlabel metal1 12236 13974 12236 13974 0 _0315_
rlabel metal2 26726 13532 26726 13532 0 _0316_
rlabel metal1 26036 36890 26036 36890 0 _0317_
rlabel metal2 12926 32164 12926 32164 0 _0318_
rlabel metal2 25990 32028 25990 32028 0 _0319_
rlabel metal1 4738 36890 4738 36890 0 _0320_
rlabel metal2 25806 9180 25806 9180 0 _0321_
rlabel metal2 22126 19074 22126 19074 0 _0322_
rlabel metal1 19596 43418 19596 43418 0 _0323_
rlabel metal1 14858 27574 14858 27574 0 _0324_
rlabel metal1 24380 6698 24380 6698 0 _0325_
rlabel metal2 27370 29410 27370 29410 0 _0326_
rlabel metal1 23046 4114 23046 4114 0 _0327_
rlabel metal2 22218 38692 22218 38692 0 _0328_
rlabel metal1 2806 6222 2806 6222 0 _0329_
rlabel metal2 20470 45730 20470 45730 0 _0330_
rlabel metal1 12972 3162 12972 3162 0 _0331_
rlabel metal2 26726 10268 26726 10268 0 _0332_
rlabel metal1 1978 7174 1978 7174 0 _0333_
rlabel metal2 2438 11492 2438 11492 0 _0334_
rlabel metal2 3266 37740 3266 37740 0 _0335_
rlabel metal2 28198 15708 28198 15708 0 _0336_
rlabel metal2 26726 42840 26726 42840 0 _0337_
rlabel metal2 27922 38658 27922 38658 0 _0338_
rlabel metal1 4140 45526 4140 45526 0 _0339_
rlabel metal2 27922 44642 27922 44642 0 _0340_
rlabel metal2 20562 3740 20562 3740 0 _0341_
rlabel metal2 27278 3298 27278 3298 0 _0342_
rlabel metal2 23138 46308 23138 46308 0 _0343_
rlabel metal2 19642 3196 19642 3196 0 _0344_
rlabel metal2 27738 10336 27738 10336 0 _0345_
rlabel metal1 2024 26214 2024 26214 0 _0346_
rlabel metal2 27370 23970 27370 23970 0 _0347_
rlabel metal1 2714 44506 2714 44506 0 _0348_
rlabel metal1 3450 2346 3450 2346 0 _0349_
rlabel metal2 7130 3230 7130 3230 0 _0350_
rlabel metal2 2070 13090 2070 13090 0 _0351_
rlabel metal2 28198 32402 28198 32402 0 _0352_
rlabel metal2 27922 21794 27922 21794 0 _0353_
rlabel metal2 27370 20162 27370 20162 0 _0354_
rlabel metal1 2116 5338 2116 5338 0 _0355_
rlabel metal2 2070 45220 2070 45220 0 _0356_
rlabel metal1 27048 12614 27048 12614 0 _0357_
rlabel metal2 10626 3740 10626 3740 0 _0358_
rlabel metal1 18308 46138 18308 46138 0 _0359_
rlabel metal1 2668 46614 2668 46614 0 _0360_
rlabel metal2 27830 27234 27830 27234 0 _0361_
rlabel metal2 3266 41820 3266 41820 0 _0362_
rlabel metal2 4186 8092 4186 8092 0 _0363_
rlabel metal2 9522 46546 9522 46546 0 _0364_
rlabel metal2 10166 46308 10166 46308 0 _0365_
rlabel metal1 27094 7310 27094 7310 0 _0366_
rlabel metal2 28198 41820 28198 41820 0 _0367_
rlabel metal1 13156 45594 13156 45594 0 _0368_
rlabel metal1 28014 4250 28014 4250 0 _0369_
rlabel metal1 27002 35802 27002 35802 0 _0370_
rlabel metal2 2346 40324 2346 40324 0 _0371_
rlabel metal1 27140 3094 27140 3094 0 _0372_
rlabel metal2 1794 20060 1794 20060 0 _0373_
rlabel metal2 28198 8092 28198 8092 0 _0374_
rlabel metal2 1886 40222 1886 40222 0 _0375_
rlabel metal2 1978 17442 1978 17442 0 _0376_
rlabel metal2 1794 9180 1794 9180 0 _0377_
rlabel metal2 1794 14620 1794 14620 0 _0378_
rlabel metal3 1786 36788 1786 36788 0 active
rlabel metal2 20838 28866 20838 28866 0 clknet_0_wb_clk_i
rlabel metal2 21298 14144 21298 14144 0 clknet_2_0__leaf_wb_clk_i
rlabel metal2 23506 20043 23506 20043 0 clknet_2_1__leaf_wb_clk_i
rlabel metal1 19136 32334 19136 32334 0 clknet_2_2__leaf_wb_clk_i
rlabel metal1 24058 34034 24058 34034 0 clknet_2_3__leaf_wb_clk_i
rlabel metal2 21206 33558 21206 33558 0 frequency_counter_0.clk_counter\[0\]
rlabel metal2 20286 27540 20286 27540 0 frequency_counter_0.clk_counter\[10\]
rlabel metal2 19596 11220 19596 11220 0 frequency_counter_0.clk_counter\[11\]
rlabel metal1 20700 33966 20700 33966 0 frequency_counter_0.clk_counter\[1\]
rlabel metal1 21160 36142 21160 36142 0 frequency_counter_0.clk_counter\[2\]
rlabel metal1 20884 39406 20884 39406 0 frequency_counter_0.clk_counter\[3\]
rlabel metal2 18262 37740 18262 37740 0 frequency_counter_0.clk_counter\[4\]
rlabel metal1 18216 40086 18216 40086 0 frequency_counter_0.clk_counter\[5\]
rlabel metal2 16698 30260 16698 30260 0 frequency_counter_0.clk_counter\[6\]
rlabel metal1 16974 32878 16974 32878 0 frequency_counter_0.clk_counter\[7\]
rlabel metal1 17250 21658 17250 21658 0 frequency_counter_0.clk_counter\[8\]
rlabel via2 18814 24667 18814 24667 0 frequency_counter_0.clk_counter\[9\]
rlabel metal2 24518 27472 24518 27472 0 frequency_counter_0.dbg_edge_count\[0\]
rlabel metal1 25530 17510 25530 17510 0 frequency_counter_0.dbg_edge_count\[1\]
rlabel metal1 22862 31994 22862 31994 0 frequency_counter_0.dbg_edge_count\[2\]
rlabel metal1 20792 18258 20792 18258 0 frequency_counter_0.dbg_state\[0\]
rlabel metal1 20838 19380 20838 19380 0 frequency_counter_0.dbg_state\[1\]
rlabel metal2 25806 32844 25806 32844 0 frequency_counter_0.digit
rlabel metal1 24058 32912 24058 32912 0 frequency_counter_0.edge_counter\[0\]
rlabel metal1 26910 20434 26910 20434 0 frequency_counter_0.edge_counter\[1\]
rlabel metal1 25576 21998 25576 21998 0 frequency_counter_0.edge_counter\[2\]
rlabel metal1 26220 25874 26220 25874 0 frequency_counter_0.edge_counter\[3\]
rlabel metal2 27738 34748 27738 34748 0 frequency_counter_0.edge_detect0.q0
rlabel metal1 25484 34714 25484 34714 0 frequency_counter_0.edge_detect0.q1
rlabel metal2 25898 33354 25898 33354 0 frequency_counter_0.edge_detect0.q2
rlabel metal1 11454 14518 11454 14518 0 frequency_counter_0.segments\[0\]
rlabel metal1 18170 14586 18170 14586 0 frequency_counter_0.segments\[1\]
rlabel metal1 10166 13974 10166 13974 0 frequency_counter_0.segments\[2\]
rlabel metal1 13938 13838 13938 13838 0 frequency_counter_0.segments\[3\]
rlabel metal1 14904 13906 14904 13906 0 frequency_counter_0.segments\[4\]
rlabel metal1 25346 37230 25346 37230 0 frequency_counter_0.segments\[5\]
rlabel metal1 13018 32266 13018 32266 0 frequency_counter_0.segments\[6\]
rlabel metal2 21022 11968 21022 11968 0 frequency_counter_0.seven_segment0.load
rlabel metal1 22678 15946 22678 15946 0 frequency_counter_0.seven_segment0.ten_count\[0\]
rlabel metal1 20930 11628 20930 11628 0 frequency_counter_0.seven_segment0.ten_count\[1\]
rlabel metal1 20838 12104 20838 12104 0 frequency_counter_0.seven_segment0.ten_count\[2\]
rlabel metal1 21827 11118 21827 11118 0 frequency_counter_0.seven_segment0.ten_count\[3\]
rlabel metal1 21620 16422 21620 16422 0 frequency_counter_0.seven_segment0.ten_count_reg\[0\]
rlabel metal1 20654 11866 20654 11866 0 frequency_counter_0.seven_segment0.ten_count_reg\[1\]
rlabel metal1 20792 12206 20792 12206 0 frequency_counter_0.seven_segment0.ten_count_reg\[2\]
rlabel metal2 22678 14790 22678 14790 0 frequency_counter_0.seven_segment0.ten_count_reg\[3\]
rlabel metal2 21298 26469 21298 26469 0 frequency_counter_0.seven_segment0.unit_count\[0\]
rlabel metal1 21482 26554 21482 26554 0 frequency_counter_0.seven_segment0.unit_count\[1\]
rlabel metal1 21390 20774 21390 20774 0 frequency_counter_0.seven_segment0.unit_count\[2\]
rlabel metal2 21666 24582 21666 24582 0 frequency_counter_0.seven_segment0.unit_count\[3\]
rlabel metal1 21574 21862 21574 21862 0 frequency_counter_0.seven_segment0.unit_count_reg\[0\]
rlabel metal1 20838 15538 20838 15538 0 frequency_counter_0.seven_segment0.unit_count_reg\[1\]
rlabel metal1 20516 20230 20516 20230 0 frequency_counter_0.seven_segment0.unit_count_reg\[2\]
rlabel metal1 21620 15470 21620 15470 0 frequency_counter_0.seven_segment0.unit_count_reg\[3\]
rlabel metal1 18998 26010 18998 26010 0 frequency_counter_0.update_period\[0\]
rlabel metal1 17848 17170 17848 17170 0 frequency_counter_0.update_period\[10\]
rlabel metal2 20470 16150 20470 16150 0 frequency_counter_0.update_period\[11\]
rlabel metal1 20010 36074 20010 36074 0 frequency_counter_0.update_period\[1\]
rlabel metal2 23414 37094 23414 37094 0 frequency_counter_0.update_period\[2\]
rlabel metal2 25070 34272 25070 34272 0 frequency_counter_0.update_period\[3\]
rlabel metal1 18124 38318 18124 38318 0 frequency_counter_0.update_period\[4\]
rlabel metal1 15456 19822 15456 19822 0 frequency_counter_0.update_period\[5\]
rlabel metal1 16606 33490 16606 33490 0 frequency_counter_0.update_period\[6\]
rlabel metal1 15962 33286 15962 33286 0 frequency_counter_0.update_period\[7\]
rlabel metal2 18078 18836 18078 18836 0 frequency_counter_0.update_period\[8\]
rlabel metal1 24909 18938 24909 18938 0 frequency_counter_0.update_period\[9\]
rlabel metal2 28382 37009 28382 37009 0 io_in[8]
rlabel metal2 21298 2166 21298 2166 0 io_oeb[0]
rlabel metal3 1142 13668 1142 13668 0 io_oeb[10]
rlabel via2 27554 32963 27554 32963 0 io_oeb[11]
rlabel metal2 27554 22015 27554 22015 0 io_oeb[12]
rlabel metal3 28850 21148 28850 21148 0 io_oeb[13]
rlabel metal3 1878 3468 1878 3468 0 io_oeb[14]
rlabel metal1 2162 45356 2162 45356 0 io_oeb[15]
rlabel metal3 28850 12308 28850 12308 0 io_oeb[16]
rlabel metal2 10994 2166 10994 2166 0 io_oeb[17]
rlabel metal2 18722 47882 18722 47882 0 io_oeb[18]
rlabel metal1 2392 46478 2392 46478 0 io_oeb[19]
rlabel metal3 28436 1428 28436 1428 0 io_oeb[1]
rlabel via2 27554 27523 27554 27523 0 io_oeb[20]
rlabel metal3 1142 41548 1142 41548 0 io_oeb[21]
rlabel metal2 3910 2200 3910 2200 0 io_oeb[22]
rlabel metal2 10350 48188 10350 48188 0 io_oeb[23]
rlabel metal2 10994 47882 10994 47882 0 io_oeb[24]
rlabel metal2 26174 7769 26174 7769 0 io_oeb[25]
rlabel metal2 27554 41599 27554 41599 0 io_oeb[26]
rlabel metal2 13570 47882 13570 47882 0 io_oeb[27]
rlabel metal2 27462 4063 27462 4063 0 io_oeb[28]
rlabel metal3 28850 36108 28850 36108 0 io_oeb[29]
rlabel metal1 23368 46478 23368 46478 0 io_oeb[2]
rlabel metal2 2806 41633 2806 41633 0 io_oeb[30]
rlabel metal2 26174 2873 26174 2873 0 io_oeb[31]
rlabel metal2 2806 19839 2806 19839 0 io_oeb[32]
rlabel metal2 27554 8415 27554 8415 0 io_oeb[33]
rlabel metal3 2108 49708 2108 49708 0 io_oeb[34]
rlabel via2 2806 17731 2806 17731 0 io_oeb[35]
rlabel metal3 1740 8908 1740 8908 0 io_oeb[36]
rlabel metal2 2806 14399 2806 14399 0 io_oeb[37]
rlabel metal2 20010 1622 20010 1622 0 io_oeb[3]
rlabel metal2 27554 10727 27554 10727 0 io_oeb[4]
rlabel metal3 1740 25908 1740 25908 0 io_oeb[5]
rlabel metal3 28850 24548 28850 24548 0 io_oeb[6]
rlabel metal2 881 49300 881 49300 0 io_oeb[7]
rlabel metal2 3266 1622 3266 1622 0 io_oeb[8]
rlabel metal2 8418 1860 8418 1860 0 io_oeb[9]
rlabel metal3 28804 47668 28804 47668 0 io_out[0]
rlabel metal3 28804 32028 28804 32028 0 io_out[10]
rlabel metal3 2108 2108 2108 2108 0 io_out[11]
rlabel metal3 2154 6188 2154 6188 0 io_out[12]
rlabel metal3 28727 2516 28727 2516 0 io_out[13]
rlabel metal2 26082 39797 26082 39797 0 io_out[14]
rlabel metal3 2108 33388 2108 33388 0 io_out[15]
rlabel metal3 28436 31348 28436 31348 0 io_out[16]
rlabel metal1 23414 37128 23414 37128 0 io_out[17]
rlabel metal3 29846 7548 29846 7548 0 io_out[18]
rlabel metal2 3358 18887 3358 18887 0 io_out[19]
rlabel metal2 16790 47644 16790 47644 0 io_out[1]
rlabel metal2 22586 47576 22586 47576 0 io_out[20]
rlabel metal3 1832 32028 1832 32028 0 io_out[21]
rlabel metal2 25162 3798 25162 3798 0 io_out[22]
rlabel metal3 28436 28628 28436 28628 0 io_out[23]
rlabel metal2 21942 1367 21942 1367 0 io_out[24]
rlabel metal2 23506 42874 23506 42874 0 io_out[25]
rlabel metal3 2384 4148 2384 4148 0 io_out[26]
rlabel metal2 21298 47644 21298 47644 0 io_out[27]
rlabel metal2 13570 1367 13570 1367 0 io_out[28]
rlabel metal3 29846 10948 29846 10948 0 io_out[29]
rlabel metal2 5842 2710 5842 2710 0 io_out[2]
rlabel metal3 1740 4828 1740 4828 0 io_out[30]
rlabel metal3 1740 11628 1740 11628 0 io_out[31]
rlabel metal3 1142 37468 1142 37468 0 io_out[32]
rlabel metal2 27554 15623 27554 15623 0 io_out[33]
rlabel metal3 28850 42908 28850 42908 0 io_out[34]
rlabel metal3 28988 40868 28988 40868 0 io_out[35]
rlabel metal1 3542 46002 3542 46002 0 io_out[36]
rlabel metal3 28436 46308 28436 46308 0 io_out[37]
rlabel metal2 2806 34629 2806 34629 0 io_out[3]
rlabel via2 27554 34051 27554 34051 0 io_out[4]
rlabel metal2 8418 47882 8418 47882 0 io_out[5]
rlabel metal2 28382 48188 28382 48188 0 io_out[6]
rlabel metal2 2806 15861 2806 15861 0 io_out[7]
rlabel metal2 14858 1231 14858 1231 0 io_out[8]
rlabel metal3 2154 12308 2154 12308 0 io_out[9]
rlabel via2 27370 16541 27370 16541 0 la1_data_in[0]
rlabel metal2 17434 1588 17434 1588 0 la1_data_in[10]
rlabel metal1 28428 13906 28428 13906 0 la1_data_in[11]
rlabel metal3 1142 29988 1142 29988 0 la1_data_in[12]
rlabel metal2 27094 1588 27094 1588 0 la1_data_in[13]
rlabel metal2 16146 1554 16146 1554 0 la1_data_in[1]
rlabel metal2 9062 1588 9062 1588 0 la1_data_in[2]
rlabel metal3 1142 25228 1142 25228 0 la1_data_in[3]
rlabel metal2 24058 48161 24058 48161 0 la1_data_in[4]
rlabel metal2 28382 30107 28382 30107 0 la1_data_in[5]
rlabel metal2 5842 48154 5842 48154 0 la1_data_in[6]
rlabel metal3 1142 18428 1142 18428 0 la1_data_in[7]
rlabel metal1 6532 47022 6532 47022 0 la1_data_in[8]
rlabel metal3 1142 27948 1142 27948 0 la1_data_in[9]
rlabel metal2 6486 2166 6486 2166 0 la1_data_out[0]
rlabel metal1 26358 17714 26358 17714 0 la1_data_out[10]
rlabel metal2 18078 1826 18078 1826 0 la1_data_out[11]
rlabel metal2 26082 46189 26082 46189 0 la1_data_out[12]
rlabel metal2 4186 43741 4186 43741 0 la1_data_out[13]
rlabel metal2 11822 46767 11822 46767 0 la1_data_out[14]
rlabel metal3 1740 1428 1740 1428 0 la1_data_out[15]
rlabel metal3 29846 23868 29846 23868 0 la1_data_out[16]
rlabel metal2 26174 39185 26174 39185 0 la1_data_out[17]
rlabel metal2 2806 43843 2806 43843 0 la1_data_out[18]
rlabel metal2 26174 30957 26174 30957 0 la1_data_out[19]
rlabel metal3 1740 36108 1740 36108 0 la1_data_out[1]
rlabel metal3 2384 8228 2384 8228 0 la1_data_out[20]
rlabel metal3 28712 44948 28712 44948 0 la1_data_out[21]
rlabel metal2 15226 46189 15226 46189 0 la1_data_out[22]
rlabel metal2 9706 1860 9706 1860 0 la1_data_out[23]
rlabel metal3 28850 25228 28850 25228 0 la1_data_out[24]
rlabel metal3 1786 2788 1786 2788 0 la1_data_out[25]
rlabel metal3 28850 14348 28850 14348 0 la1_data_out[26]
rlabel metal3 1740 38828 1740 38828 0 la1_data_out[27]
rlabel metal3 29846 5508 29846 5508 0 la1_data_out[28]
rlabel metal2 4554 1231 4554 1231 0 la1_data_out[29]
rlabel metal2 16790 1860 16790 1860 0 la1_data_out[2]
rlabel metal3 28850 20468 28850 20468 0 la1_data_out[30]
rlabel metal2 26174 46665 26174 46665 0 la1_data_out[31]
rlabel metal3 1740 7548 1740 7548 0 la1_data_out[3]
rlabel metal2 26174 6545 26174 6545 0 la1_data_out[4]
rlabel metal2 2622 1503 2622 1503 0 la1_data_out[5]
rlabel metal3 28390 26588 28390 26588 0 la1_data_out[6]
rlabel metal2 690 2200 690 2200 0 la1_data_out[7]
rlabel via2 27554 40579 27554 40579 0 la1_data_out[8]
rlabel metal2 27738 47644 27738 47644 0 la1_data_out[9]
rlabel metal1 3220 36822 3220 36822 0 net1
rlabel metal2 15778 25432 15778 25432 0 net10
rlabel metal2 1702 41548 1702 41548 0 net100
rlabel metal2 26634 4012 26634 4012 0 net101
rlabel metal1 1656 19346 1656 19346 0 net102
rlabel metal2 28382 8432 28382 8432 0 net103
rlabel metal1 2070 39950 2070 39950 0 net104
rlabel metal2 1610 17884 1610 17884 0 net105
rlabel metal2 1610 9180 1610 9180 0 net106
rlabel metal1 1656 13906 1656 13906 0 net107
rlabel metal1 26787 34646 26787 34646 0 net108
rlabel via1 24973 33966 24973 33966 0 net109
rlabel metal1 23598 37230 23598 37230 0 net11
rlabel metal1 27140 33422 27140 33422 0 net12
rlabel metal2 6026 41820 6026 41820 0 net13
rlabel metal2 15686 19142 15686 19142 0 net14
rlabel metal2 6762 41990 6762 41990 0 net15
rlabel metal2 1794 27608 1794 27608 0 net16
rlabel metal1 5520 3502 5520 3502 0 net17
rlabel metal1 1610 36244 1610 36244 0 net18
rlabel metal2 16238 3264 16238 3264 0 net19
rlabel metal1 28121 34986 28121 34986 0 net2
rlabel metal2 1702 9248 1702 9248 0 net20
rlabel metal2 26634 6528 26634 6528 0 net21
rlabel metal2 2990 4964 2990 4964 0 net22
rlabel metal2 26542 28798 26542 28798 0 net23
rlabel metal2 1610 4080 1610 4080 0 net24
rlabel metal2 28382 40732 28382 40732 0 net25
rlabel metal2 26542 46172 26542 46172 0 net26
rlabel metal2 28382 18224 28382 18224 0 net27
rlabel metal2 19182 3230 19182 3230 0 net28
rlabel metal1 27278 45458 27278 45458 0 net29
rlabel metal2 26450 16966 26450 16966 0 net3
rlabel metal2 2990 43724 2990 43724 0 net30
rlabel metal1 11546 46002 11546 46002 0 net31
rlabel metal1 1840 2618 1840 2618 0 net32
rlabel metal2 26542 23324 26542 23324 0 net33
rlabel metal1 27094 38930 27094 38930 0 net34
rlabel metal2 1610 43248 1610 43248 0 net35
rlabel metal1 27278 32198 27278 32198 0 net36
rlabel metal2 3082 9792 3082 9792 0 net37
rlabel metal2 26266 44336 26266 44336 0 net38
rlabel metal2 14214 45696 14214 45696 0 net39
rlabel metal1 17480 13906 17480 13906 0 net4
rlabel metal2 9246 3264 9246 3264 0 net40
rlabel metal1 27784 24786 27784 24786 0 net41
rlabel metal2 3726 4352 3726 4352 0 net42
rlabel metal1 26542 14484 26542 14484 0 net43
rlabel metal2 4002 38284 4002 38284 0 net44
rlabel metal1 26818 5202 26818 5202 0 net45
rlabel metal2 4186 4352 4186 4352 0 net46
rlabel metal1 27232 19890 27232 19890 0 net47
rlabel metal1 24886 44302 24886 44302 0 net48
rlabel metal1 26864 37842 26864 37842 0 net49
rlabel metal1 27922 14042 27922 14042 0 net5
rlabel metal2 15962 46240 15962 46240 0 net50
rlabel metal1 5060 4590 5060 4590 0 net51
rlabel metal2 1702 34816 1702 34816 0 net52
rlabel metal1 28198 34034 28198 34034 0 net53
rlabel metal2 7038 46784 7038 46784 0 net54
rlabel metal2 26634 46750 26634 46750 0 net55
rlabel metal2 1702 15844 1702 15844 0 net56
rlabel metal2 14030 3264 14030 3264 0 net57
rlabel metal1 3036 7174 3036 7174 0 net58
rlabel metal2 20286 46172 20286 46172 0 net59
rlabel metal2 1840 27268 1840 27268 0 net6
rlabel metal1 12880 3706 12880 3706 0 net60
rlabel metal1 26542 10132 26542 10132 0 net61
rlabel metal1 1656 6290 1656 6290 0 net62
rlabel metal2 1702 11492 1702 11492 0 net63
rlabel metal2 3450 38012 3450 38012 0 net64
rlabel metal2 28382 15708 28382 15708 0 net65
rlabel metal1 26864 42738 26864 42738 0 net66
rlabel metal2 26542 39644 26542 39644 0 net67
rlabel metal1 3680 45050 3680 45050 0 net68
rlabel metal2 28382 45084 28382 45084 0 net69
rlabel metal1 26174 2618 26174 2618 0 net7
rlabel metal2 20378 3740 20378 3740 0 net70
rlabel metal1 26312 3502 26312 3502 0 net71
rlabel metal2 22862 46784 22862 46784 0 net72
rlabel metal2 19458 2992 19458 2992 0 net73
rlabel metal1 28244 10642 28244 10642 0 net74
rlabel metal2 1702 25636 1702 25636 0 net75
rlabel metal1 27922 23732 27922 23732 0 net76
rlabel metal1 2990 43962 2990 43962 0 net77
rlabel metal1 3726 2414 3726 2414 0 net78
rlabel metal2 6946 3434 6946 3434 0 net79
rlabel metal1 16376 2550 16376 2550 0 net8
rlabel metal2 3450 13600 3450 13600 0 net80
rlabel metal1 27922 32402 27922 32402 0 net81
rlabel metal1 28244 22066 28244 22066 0 net82
rlabel metal1 27830 19278 27830 19278 0 net83
rlabel metal1 1656 5202 1656 5202 0 net84
rlabel metal2 1702 45900 1702 45900 0 net85
rlabel metal1 27232 12682 27232 12682 0 net86
rlabel metal1 10212 3502 10212 3502 0 net87
rlabel metal2 18262 46784 18262 46784 0 net88
rlabel metal1 2300 46546 2300 46546 0 net89
rlabel metal1 9476 2482 9476 2482 0 net9
rlabel metal1 28244 27506 28244 27506 0 net90
rlabel metal2 3450 41820 3450 41820 0 net91
rlabel metal2 4002 8092 4002 8092 0 net92
rlabel metal1 9522 45458 9522 45458 0 net93
rlabel metal1 9890 46410 9890 46410 0 net94
rlabel metal2 26634 7820 26634 7820 0 net95
rlabel metal1 28382 41684 28382 41684 0 net96
rlabel metal2 12926 46784 12926 46784 0 net97
rlabel metal1 28244 3026 28244 3026 0 net98
rlabel metal1 27232 36210 27232 36210 0 net99
rlabel metal1 24472 25262 24472 25262 0 wb_clk_i
<< properties >>
string FIXED_BBOX 0 0 30000 50000
<< end >>
