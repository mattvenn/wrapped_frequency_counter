magic
tech sky130A
magscale 1 2
timestamp 1647448632
<< obsli1 >>
rect 1104 2159 48852 17425
<< obsm1 >>
rect 658 1028 49666 17536
<< metal2 >>
rect -10 19200 102 20000
rect 634 19200 746 20000
rect 1278 19200 1390 20000
rect 1922 19200 2034 20000
rect 2566 19200 2678 20000
rect 3210 19200 3322 20000
rect 3854 19200 3966 20000
rect 4498 19200 4610 20000
rect 5142 19200 5254 20000
rect 5786 19200 5898 20000
rect 6430 19200 6542 20000
rect 7074 19200 7186 20000
rect 7718 19200 7830 20000
rect 8362 19200 8474 20000
rect 9006 19200 9118 20000
rect 9650 19200 9762 20000
rect 10294 19200 10406 20000
rect 10938 19200 11050 20000
rect 11582 19200 11694 20000
rect 12226 19200 12338 20000
rect 12870 19200 12982 20000
rect 13514 19200 13626 20000
rect 14158 19200 14270 20000
rect 14802 19200 14914 20000
rect 16090 19200 16202 20000
rect 16734 19200 16846 20000
rect 17378 19200 17490 20000
rect 18022 19200 18134 20000
rect 18666 19200 18778 20000
rect 19310 19200 19422 20000
rect 19954 19200 20066 20000
rect 20598 19200 20710 20000
rect 21242 19200 21354 20000
rect 21886 19200 21998 20000
rect 22530 19200 22642 20000
rect 23174 19200 23286 20000
rect 23818 19200 23930 20000
rect 24462 19200 24574 20000
rect 25106 19200 25218 20000
rect 25750 19200 25862 20000
rect 26394 19200 26506 20000
rect 27038 19200 27150 20000
rect 27682 19200 27794 20000
rect 28326 19200 28438 20000
rect 28970 19200 29082 20000
rect 29614 19200 29726 20000
rect 30258 19200 30370 20000
rect 30902 19200 31014 20000
rect 31546 19200 31658 20000
rect 32190 19200 32302 20000
rect 32834 19200 32946 20000
rect 33478 19200 33590 20000
rect 34122 19200 34234 20000
rect 34766 19200 34878 20000
rect 35410 19200 35522 20000
rect 36054 19200 36166 20000
rect 36698 19200 36810 20000
rect 37342 19200 37454 20000
rect 37986 19200 38098 20000
rect 38630 19200 38742 20000
rect 39274 19200 39386 20000
rect 39918 19200 40030 20000
rect 40562 19200 40674 20000
rect 41206 19200 41318 20000
rect 41850 19200 41962 20000
rect 42494 19200 42606 20000
rect 43138 19200 43250 20000
rect 43782 19200 43894 20000
rect 44426 19200 44538 20000
rect 45070 19200 45182 20000
rect 45714 19200 45826 20000
rect 46358 19200 46470 20000
rect 47002 19200 47114 20000
rect 47646 19200 47758 20000
rect 48290 19200 48402 20000
rect 48934 19200 49046 20000
rect 49578 19200 49690 20000
rect -10 0 102 800
rect 634 0 746 800
rect 1278 0 1390 800
rect 1922 0 2034 800
rect 2566 0 2678 800
rect 3210 0 3322 800
rect 3854 0 3966 800
rect 4498 0 4610 800
rect 5142 0 5254 800
rect 5786 0 5898 800
rect 6430 0 6542 800
rect 7074 0 7186 800
rect 7718 0 7830 800
rect 8362 0 8474 800
rect 9006 0 9118 800
rect 9650 0 9762 800
rect 10294 0 10406 800
rect 10938 0 11050 800
rect 11582 0 11694 800
rect 12226 0 12338 800
rect 12870 0 12982 800
rect 13514 0 13626 800
rect 14158 0 14270 800
rect 14802 0 14914 800
rect 15446 0 15558 800
rect 16090 0 16202 800
rect 16734 0 16846 800
rect 17378 0 17490 800
rect 18022 0 18134 800
rect 18666 0 18778 800
rect 19310 0 19422 800
rect 19954 0 20066 800
rect 20598 0 20710 800
rect 21242 0 21354 800
rect 21886 0 21998 800
rect 22530 0 22642 800
rect 23174 0 23286 800
rect 23818 0 23930 800
rect 24462 0 24574 800
rect 25106 0 25218 800
rect 25750 0 25862 800
rect 26394 0 26506 800
rect 27038 0 27150 800
rect 27682 0 27794 800
rect 28326 0 28438 800
rect 28970 0 29082 800
rect 29614 0 29726 800
rect 30258 0 30370 800
rect 30902 0 31014 800
rect 31546 0 31658 800
rect 32190 0 32302 800
rect 32834 0 32946 800
rect 33478 0 33590 800
rect 34766 0 34878 800
rect 35410 0 35522 800
rect 36054 0 36166 800
rect 36698 0 36810 800
rect 37342 0 37454 800
rect 37986 0 38098 800
rect 38630 0 38742 800
rect 39274 0 39386 800
rect 39918 0 40030 800
rect 40562 0 40674 800
rect 41206 0 41318 800
rect 41850 0 41962 800
rect 42494 0 42606 800
rect 43138 0 43250 800
rect 43782 0 43894 800
rect 44426 0 44538 800
rect 45070 0 45182 800
rect 45714 0 45826 800
rect 46358 0 46470 800
rect 47002 0 47114 800
rect 47646 0 47758 800
rect 48290 0 48402 800
rect 48934 0 49046 800
rect 49578 0 49690 800
<< obsm2 >>
rect 802 19144 1222 19200
rect 1446 19144 1866 19200
rect 2090 19144 2510 19200
rect 2734 19144 3154 19200
rect 3378 19144 3798 19200
rect 4022 19144 4442 19200
rect 4666 19144 5086 19200
rect 5310 19144 5730 19200
rect 5954 19144 6374 19200
rect 6598 19144 7018 19200
rect 7242 19144 7662 19200
rect 7886 19144 8306 19200
rect 8530 19144 8950 19200
rect 9174 19144 9594 19200
rect 9818 19144 10238 19200
rect 10462 19144 10882 19200
rect 11106 19144 11526 19200
rect 11750 19144 12170 19200
rect 12394 19144 12814 19200
rect 13038 19144 13458 19200
rect 13682 19144 14102 19200
rect 14326 19144 14746 19200
rect 14970 19144 16034 19200
rect 16258 19144 16678 19200
rect 16902 19144 17322 19200
rect 17546 19144 17966 19200
rect 18190 19144 18610 19200
rect 18834 19144 19254 19200
rect 19478 19144 19898 19200
rect 20122 19144 20542 19200
rect 20766 19144 21186 19200
rect 21410 19144 21830 19200
rect 22054 19144 22474 19200
rect 22698 19144 23118 19200
rect 23342 19144 23762 19200
rect 23986 19144 24406 19200
rect 24630 19144 25050 19200
rect 25274 19144 25694 19200
rect 25918 19144 26338 19200
rect 26562 19144 26982 19200
rect 27206 19144 27626 19200
rect 27850 19144 28270 19200
rect 28494 19144 28914 19200
rect 29138 19144 29558 19200
rect 29782 19144 30202 19200
rect 30426 19144 30846 19200
rect 31070 19144 31490 19200
rect 31714 19144 32134 19200
rect 32358 19144 32778 19200
rect 33002 19144 33422 19200
rect 33646 19144 34066 19200
rect 34290 19144 34710 19200
rect 34934 19144 35354 19200
rect 35578 19144 35998 19200
rect 36222 19144 36642 19200
rect 36866 19144 37286 19200
rect 37510 19144 37930 19200
rect 38154 19144 38574 19200
rect 38798 19144 39218 19200
rect 39442 19144 39862 19200
rect 40086 19144 40506 19200
rect 40730 19144 41150 19200
rect 41374 19144 41794 19200
rect 42018 19144 42438 19200
rect 42662 19144 43082 19200
rect 43306 19144 43726 19200
rect 43950 19144 44370 19200
rect 44594 19144 45014 19200
rect 45238 19144 45658 19200
rect 45882 19144 46302 19200
rect 46526 19144 46946 19200
rect 47170 19144 47590 19200
rect 47814 19144 48234 19200
rect 48458 19144 48878 19200
rect 49102 19144 49522 19200
rect 664 856 49660 19144
rect 802 31 1222 856
rect 1446 31 1866 856
rect 2090 31 2510 856
rect 2734 31 3154 856
rect 3378 31 3798 856
rect 4022 31 4442 856
rect 4666 31 5086 856
rect 5310 31 5730 856
rect 5954 31 6374 856
rect 6598 31 7018 856
rect 7242 31 7662 856
rect 7886 31 8306 856
rect 8530 31 8950 856
rect 9174 31 9594 856
rect 9818 31 10238 856
rect 10462 31 10882 856
rect 11106 31 11526 856
rect 11750 31 12170 856
rect 12394 31 12814 856
rect 13038 31 13458 856
rect 13682 31 14102 856
rect 14326 31 14746 856
rect 14970 31 15390 856
rect 15614 31 16034 856
rect 16258 31 16678 856
rect 16902 31 17322 856
rect 17546 31 17966 856
rect 18190 31 18610 856
rect 18834 31 19254 856
rect 19478 31 19898 856
rect 20122 31 20542 856
rect 20766 31 21186 856
rect 21410 31 21830 856
rect 22054 31 22474 856
rect 22698 31 23118 856
rect 23342 31 23762 856
rect 23986 31 24406 856
rect 24630 31 25050 856
rect 25274 31 25694 856
rect 25918 31 26338 856
rect 26562 31 26982 856
rect 27206 31 27626 856
rect 27850 31 28270 856
rect 28494 31 28914 856
rect 29138 31 29558 856
rect 29782 31 30202 856
rect 30426 31 30846 856
rect 31070 31 31490 856
rect 31714 31 32134 856
rect 32358 31 32778 856
rect 33002 31 33422 856
rect 33646 31 34710 856
rect 34934 31 35354 856
rect 35578 31 35998 856
rect 36222 31 36642 856
rect 36866 31 37286 856
rect 37510 31 37930 856
rect 38154 31 38574 856
rect 38798 31 39218 856
rect 39442 31 39862 856
rect 40086 31 40506 856
rect 40730 31 41150 856
rect 41374 31 41794 856
rect 42018 31 42438 856
rect 42662 31 43082 856
rect 43306 31 43726 856
rect 43950 31 44370 856
rect 44594 31 45014 856
rect 45238 31 45658 856
rect 45882 31 46302 856
rect 46526 31 46946 856
rect 47170 31 47590 856
rect 47814 31 48234 856
rect 48458 31 48878 856
rect 49102 31 49522 856
<< metal3 >>
rect 0 19668 800 19908
rect 0 18988 800 19228
rect 49200 18988 50000 19228
rect 0 18308 800 18548
rect 49200 18308 50000 18548
rect 0 17628 800 17868
rect 49200 17628 50000 17868
rect 0 16948 800 17188
rect 49200 16948 50000 17188
rect 0 16268 800 16508
rect 49200 16268 50000 16508
rect 0 15588 800 15828
rect 49200 15588 50000 15828
rect 0 14908 800 15148
rect 49200 14908 50000 15148
rect 0 14228 800 14468
rect 49200 14228 50000 14468
rect 0 13548 800 13788
rect 49200 13548 50000 13788
rect 0 12868 800 13108
rect 49200 12868 50000 13108
rect 0 12188 800 12428
rect 49200 12188 50000 12428
rect 0 11508 800 11748
rect 49200 11508 50000 11748
rect 0 10828 800 11068
rect 49200 10828 50000 11068
rect 0 10148 800 10388
rect 49200 10148 50000 10388
rect 0 9468 800 9708
rect 49200 9468 50000 9708
rect 0 8788 800 9028
rect 49200 8788 50000 9028
rect 0 8108 800 8348
rect 49200 8108 50000 8348
rect 0 7428 800 7668
rect 49200 7428 50000 7668
rect 0 6748 800 6988
rect 49200 6748 50000 6988
rect 0 6068 800 6308
rect 49200 6068 50000 6308
rect 0 5388 800 5628
rect 49200 5388 50000 5628
rect 0 4708 800 4948
rect 49200 4708 50000 4948
rect 0 4028 800 4268
rect 49200 4028 50000 4268
rect 0 3348 800 3588
rect 49200 3348 50000 3588
rect 0 2668 800 2908
rect 49200 2668 50000 2908
rect 0 1988 800 2228
rect 49200 1988 50000 2228
rect 0 1308 800 1548
rect 49200 1308 50000 1548
rect 0 628 800 868
rect 49200 628 50000 868
rect 49200 -52 50000 188
<< obsm3 >>
rect 880 18908 49120 19141
rect 800 18628 49200 18908
rect 880 18228 49120 18628
rect 800 17948 49200 18228
rect 880 17548 49120 17948
rect 800 17268 49200 17548
rect 880 16868 49120 17268
rect 800 16588 49200 16868
rect 880 16188 49120 16588
rect 800 15908 49200 16188
rect 880 15508 49120 15908
rect 800 15228 49200 15508
rect 880 14828 49120 15228
rect 800 14548 49200 14828
rect 880 14148 49120 14548
rect 800 13868 49200 14148
rect 880 13468 49120 13868
rect 800 13188 49200 13468
rect 880 12788 49120 13188
rect 800 12508 49200 12788
rect 880 12108 49120 12508
rect 800 11828 49200 12108
rect 880 11428 49120 11828
rect 800 11148 49200 11428
rect 880 10748 49120 11148
rect 800 10468 49200 10748
rect 880 10068 49120 10468
rect 800 9788 49200 10068
rect 880 9388 49120 9788
rect 800 9108 49200 9388
rect 880 8708 49120 9108
rect 800 8428 49200 8708
rect 880 8028 49120 8428
rect 800 7748 49200 8028
rect 880 7348 49120 7748
rect 800 7068 49200 7348
rect 880 6668 49120 7068
rect 800 6388 49200 6668
rect 880 5988 49120 6388
rect 800 5708 49200 5988
rect 880 5308 49120 5708
rect 800 5028 49200 5308
rect 880 4628 49120 5028
rect 800 4348 49200 4628
rect 880 3948 49120 4348
rect 800 3668 49200 3948
rect 880 3268 49120 3668
rect 800 2988 49200 3268
rect 880 2588 49120 2988
rect 800 2308 49200 2588
rect 880 1908 49120 2308
rect 800 1628 49200 1908
rect 880 1228 49120 1628
rect 800 948 49200 1228
rect 880 548 49120 948
rect 800 268 49200 548
rect 800 35 49120 268
<< metal4 >>
rect 8910 2128 9230 17456
rect 16874 2128 17194 17456
rect 24840 2128 25160 17456
rect 32805 2128 33125 17456
rect 40771 2128 41091 17456
<< obsm4 >>
rect 9310 2128 16794 17456
rect 17274 2128 24760 17456
rect 25240 2128 32725 17456
rect 33205 2128 40691 17456
<< labels >>
rlabel metal2 s 11582 19200 11694 20000 6 active
port 1 nsew signal input
rlabel metal2 s 10938 0 11050 800 6 io_in[0]
port 2 nsew signal input
rlabel metal2 s 34122 19200 34234 20000 6 io_in[10]
port 3 nsew signal input
rlabel metal2 s 14158 19200 14270 20000 6 io_in[11]
port 4 nsew signal input
rlabel metal3 s 49200 14228 50000 14468 6 io_in[12]
port 5 nsew signal input
rlabel metal2 s 16734 0 16846 800 6 io_in[13]
port 6 nsew signal input
rlabel metal2 s 27682 19200 27794 20000 6 io_in[14]
port 7 nsew signal input
rlabel metal3 s 49200 15588 50000 15828 6 io_in[15]
port 8 nsew signal input
rlabel metal2 s 38630 0 38742 800 6 io_in[16]
port 9 nsew signal input
rlabel metal2 s 21886 19200 21998 20000 6 io_in[17]
port 10 nsew signal input
rlabel metal2 s 23174 19200 23286 20000 6 io_in[18]
port 11 nsew signal input
rlabel metal2 s 30258 0 30370 800 6 io_in[19]
port 12 nsew signal input
rlabel metal3 s 0 11508 800 11748 6 io_in[1]
port 13 nsew signal input
rlabel metal2 s -10 19200 102 20000 6 io_in[20]
port 14 nsew signal input
rlabel metal3 s 0 13548 800 13788 6 io_in[21]
port 15 nsew signal input
rlabel metal2 s 46358 0 46470 800 6 io_in[22]
port 16 nsew signal input
rlabel metal2 s 21242 19200 21354 20000 6 io_in[23]
port 17 nsew signal input
rlabel metal2 s 19310 19200 19422 20000 6 io_in[24]
port 18 nsew signal input
rlabel metal2 s 26394 0 26506 800 6 io_in[25]
port 19 nsew signal input
rlabel metal2 s 25750 0 25862 800 6 io_in[26]
port 20 nsew signal input
rlabel metal2 s 43138 0 43250 800 6 io_in[27]
port 21 nsew signal input
rlabel metal2 s 23174 0 23286 800 6 io_in[28]
port 22 nsew signal input
rlabel metal2 s 49578 19200 49690 20000 6 io_in[29]
port 23 nsew signal input
rlabel metal2 s 11582 0 11694 800 6 io_in[2]
port 24 nsew signal input
rlabel metal2 s 48934 0 49046 800 6 io_in[30]
port 25 nsew signal input
rlabel metal2 s 10294 19200 10406 20000 6 io_in[31]
port 26 nsew signal input
rlabel metal2 s 21886 0 21998 800 6 io_in[32]
port 27 nsew signal input
rlabel metal3 s 0 18308 800 18548 6 io_in[33]
port 28 nsew signal input
rlabel metal2 s 41206 19200 41318 20000 6 io_in[34]
port 29 nsew signal input
rlabel metal2 s 45070 19200 45182 20000 6 io_in[35]
port 30 nsew signal input
rlabel metal3 s 49200 6748 50000 6988 6 io_in[36]
port 31 nsew signal input
rlabel metal2 s 45714 19200 45826 20000 6 io_in[37]
port 32 nsew signal input
rlabel metal2 s 34766 19200 34878 20000 6 io_in[3]
port 33 nsew signal input
rlabel metal3 s 49200 6068 50000 6308 6 io_in[4]
port 34 nsew signal input
rlabel metal3 s 49200 18308 50000 18548 6 io_in[5]
port 35 nsew signal input
rlabel metal2 s 1278 19200 1390 20000 6 io_in[6]
port 36 nsew signal input
rlabel metal3 s 0 14908 800 15148 6 io_in[7]
port 37 nsew signal input
rlabel metal3 s 49200 8108 50000 8348 6 io_in[8]
port 38 nsew signal input
rlabel metal2 s 20598 19200 20710 20000 6 io_in[9]
port 39 nsew signal input
rlabel metal2 s 18666 0 18778 800 6 io_oeb[0]
port 40 nsew signal output
rlabel metal3 s 0 12188 800 12428 6 io_oeb[10]
port 41 nsew signal output
rlabel metal3 s 49200 4708 50000 4948 6 io_oeb[11]
port 42 nsew signal output
rlabel metal2 s 45714 0 45826 800 6 io_oeb[12]
port 43 nsew signal output
rlabel metal2 s 45070 0 45182 800 6 io_oeb[13]
port 44 nsew signal output
rlabel metal3 s 0 3348 800 3588 6 io_oeb[14]
port 45 nsew signal output
rlabel metal2 s 24462 19200 24574 20000 6 io_oeb[15]
port 46 nsew signal output
rlabel metal2 s 37342 0 37454 800 6 io_oeb[16]
port 47 nsew signal output
rlabel metal2 s 9650 0 9762 800 6 io_oeb[17]
port 48 nsew signal output
rlabel metal2 s 39918 19200 40030 20000 6 io_oeb[18]
port 49 nsew signal output
rlabel metal2 s 25106 19200 25218 20000 6 io_oeb[19]
port 50 nsew signal output
rlabel metal2 s 27682 0 27794 800 6 io_oeb[1]
port 51 nsew signal output
rlabel metal3 s 49200 -52 50000 188 6 io_oeb[20]
port 52 nsew signal output
rlabel metal2 s 16090 19200 16202 20000 6 io_oeb[21]
port 53 nsew signal output
rlabel metal2 s 3854 0 3966 800 6 io_oeb[22]
port 54 nsew signal output
rlabel metal2 s 32190 19200 32302 20000 6 io_oeb[23]
port 55 nsew signal output
rlabel metal2 s 32834 19200 32946 20000 6 io_oeb[24]
port 56 nsew signal output
rlabel metal2 s 33478 0 33590 800 6 io_oeb[25]
port 57 nsew signal output
rlabel metal3 s 49200 12188 50000 12428 6 io_oeb[26]
port 58 nsew signal output
rlabel metal2 s 35410 19200 35522 20000 6 io_oeb[27]
port 59 nsew signal output
rlabel metal2 s 29614 0 29726 800 6 io_oeb[28]
port 60 nsew signal output
rlabel metal3 s 49200 7428 50000 7668 6 io_oeb[29]
port 61 nsew signal output
rlabel metal2 s 43782 19200 43894 20000 6 io_oeb[2]
port 62 nsew signal output
rlabel metal2 s 16734 19200 16846 20000 6 io_oeb[30]
port 63 nsew signal output
rlabel metal2 s 28970 0 29082 800 6 io_oeb[31]
port 64 nsew signal output
rlabel metal3 s 0 17628 800 17868 6 io_oeb[32]
port 65 nsew signal output
rlabel metal2 s 34766 0 34878 800 6 io_oeb[33]
port 66 nsew signal output
rlabel metal2 s 22530 19200 22642 20000 6 io_oeb[34]
port 67 nsew signal output
rlabel metal3 s 0 15588 800 15828 6 io_oeb[35]
port 68 nsew signal output
rlabel metal3 s 0 8108 800 8348 6 io_oeb[36]
port 69 nsew signal output
rlabel metal3 s 0 12868 800 13108 6 io_oeb[37]
port 70 nsew signal output
rlabel metal2 s 18022 0 18134 800 6 io_oeb[3]
port 71 nsew signal output
rlabel metal2 s 36054 0 36166 800 6 io_oeb[4]
port 72 nsew signal output
rlabel metal2 s 2566 19200 2678 20000 6 io_oeb[5]
port 73 nsew signal output
rlabel metal2 s 47646 0 47758 800 6 io_oeb[6]
port 74 nsew signal output
rlabel metal2 s 23818 19200 23930 20000 6 io_oeb[7]
port 75 nsew signal output
rlabel metal2 s 3210 0 3322 800 6 io_oeb[8]
port 76 nsew signal output
rlabel metal2 s 7718 0 7830 800 6 io_oeb[9]
port 77 nsew signal output
rlabel metal3 s 49200 17628 50000 17868 6 io_out[0]
port 78 nsew signal output
rlabel metal3 s 49200 4028 50000 4268 6 io_out[10]
port 79 nsew signal output
rlabel metal3 s 0 1988 800 2228 6 io_out[11]
port 80 nsew signal output
rlabel metal3 s 0 5388 800 5628 6 io_out[12]
port 81 nsew signal output
rlabel metal2 s 28326 0 28438 800 6 io_out[13]
port 82 nsew signal output
rlabel metal3 s 49200 12868 50000 13108 6 io_out[14]
port 83 nsew signal output
rlabel metal2 s 8362 19200 8474 20000 6 io_out[15]
port 84 nsew signal output
rlabel metal3 s 49200 3348 50000 3588 6 io_out[16]
port 85 nsew signal output
rlabel metal2 s 47002 19200 47114 20000 6 io_out[17]
port 86 nsew signal output
rlabel metal2 s 32834 0 32946 800 6 io_out[18]
port 87 nsew signal output
rlabel metal3 s 0 16948 800 17188 6 io_out[19]
port 88 nsew signal output
rlabel metal2 s 37986 19200 38098 20000 6 io_out[1]
port 89 nsew signal output
rlabel metal2 s 43138 19200 43250 20000 6 io_out[20]
port 90 nsew signal output
rlabel metal2 s 7718 19200 7830 20000 6 io_out[21]
port 91 nsew signal output
rlabel metal2 s 22530 0 22642 800 6 io_out[22]
port 92 nsew signal output
rlabel metal3 s 49200 628 50000 868 6 io_out[23]
port 93 nsew signal output
rlabel metal2 s 19310 0 19422 800 6 io_out[24]
port 94 nsew signal output
rlabel metal2 s 40562 19200 40674 20000 6 io_out[25]
port 95 nsew signal output
rlabel metal3 s 0 4028 800 4268 6 io_out[26]
port 96 nsew signal output
rlabel metal2 s 41850 19200 41962 20000 6 io_out[27]
port 97 nsew signal output
rlabel metal2 s 12226 0 12338 800 6 io_out[28]
port 98 nsew signal output
rlabel metal2 s 36698 0 36810 800 6 io_out[29]
port 99 nsew signal output
rlabel metal2 s 5142 0 5254 800 6 io_out[2]
port 100 nsew signal output
rlabel metal3 s 0 4708 800 4948 6 io_out[30]
port 101 nsew signal output
rlabel metal3 s 0 10148 800 10388 6 io_out[31]
port 102 nsew signal output
rlabel metal2 s 12226 19200 12338 20000 6 io_out[32]
port 103 nsew signal output
rlabel metal2 s 40562 0 40674 800 6 io_out[33]
port 104 nsew signal output
rlabel metal3 s 49200 13548 50000 13788 6 io_out[34]
port 105 nsew signal output
rlabel metal3 s 49200 11508 50000 11748 6 io_out[35]
port 106 nsew signal output
rlabel metal2 s 25750 19200 25862 20000 6 io_out[36]
port 107 nsew signal output
rlabel metal3 s 49200 16268 50000 16508 6 io_out[37]
port 108 nsew signal output
rlabel metal2 s 9650 19200 9762 20000 6 io_out[3]
port 109 nsew signal output
rlabel metal3 s 49200 5388 50000 5628 6 io_out[4]
port 110 nsew signal output
rlabel metal2 s 30902 19200 31014 20000 6 io_out[5]
port 111 nsew signal output
rlabel metal2 s 48290 19200 48402 20000 6 io_out[6]
port 112 nsew signal output
rlabel metal3 s 0 14228 800 14468 6 io_out[7]
port 113 nsew signal output
rlabel metal2 s 13514 0 13626 800 6 io_out[8]
port 114 nsew signal output
rlabel metal3 s 0 10828 800 11068 6 io_out[9]
port 115 nsew signal output
rlabel metal2 s 41206 0 41318 800 6 la1_data_in[0]
port 116 nsew signal input
rlabel metal2 s 15446 0 15558 800 6 la1_data_in[10]
port 117 nsew signal input
rlabel metal2 s 39918 0 40030 800 6 la1_data_in[11]
port 118 nsew signal input
rlabel metal2 s 5786 19200 5898 20000 6 la1_data_in[12]
port 119 nsew signal input
rlabel metal2 s 23818 0 23930 800 6 la1_data_in[13]
port 120 nsew signal input
rlabel metal3 s 0 9468 800 9708 6 la1_data_in[14]
port 121 nsew signal input
rlabel metal2 s 26394 19200 26506 20000 6 la1_data_in[15]
port 122 nsew signal input
rlabel metal2 s 36698 19200 36810 20000 6 la1_data_in[16]
port 123 nsew signal input
rlabel metal2 s 31546 19200 31658 20000 6 la1_data_in[17]
port 124 nsew signal input
rlabel metal2 s 30902 0 31014 800 6 la1_data_in[18]
port 125 nsew signal input
rlabel metal2 s 27038 19200 27150 20000 6 la1_data_in[19]
port 126 nsew signal input
rlabel metal2 s 14158 0 14270 800 6 la1_data_in[1]
port 127 nsew signal input
rlabel metal2 s 5142 19200 5254 20000 6 la1_data_in[20]
port 128 nsew signal input
rlabel metal2 s 48934 19200 49046 20000 6 la1_data_in[21]
port 129 nsew signal input
rlabel metal2 s 41850 0 41962 800 6 la1_data_in[22]
port 130 nsew signal input
rlabel metal3 s 0 628 800 868 6 la1_data_in[23]
port 131 nsew signal input
rlabel metal2 s 10294 0 10406 800 6 la1_data_in[24]
port 132 nsew signal input
rlabel metal2 s 6430 19200 6542 20000 6 la1_data_in[25]
port 133 nsew signal input
rlabel metal2 s 37986 0 38098 800 6 la1_data_in[26]
port 134 nsew signal input
rlabel metal2 s 20598 0 20710 800 6 la1_data_in[27]
port 135 nsew signal input
rlabel metal2 s 3210 19200 3322 20000 6 la1_data_in[28]
port 136 nsew signal input
rlabel metal2 s 14802 19200 14914 20000 6 la1_data_in[29]
port 137 nsew signal input
rlabel metal2 s 8362 0 8474 800 6 la1_data_in[2]
port 138 nsew signal input
rlabel metal2 s 1278 0 1390 800 6 la1_data_in[30]
port 139 nsew signal input
rlabel metal2 s 27038 0 27150 800 6 la1_data_in[31]
port 140 nsew signal input
rlabel metal2 s 1922 19200 2034 20000 6 la1_data_in[3]
port 141 nsew signal input
rlabel metal2 s 44426 19200 44538 20000 6 la1_data_in[4]
port 142 nsew signal input
rlabel metal3 s 49200 1988 50000 2228 6 la1_data_in[5]
port 143 nsew signal input
rlabel metal2 s 28326 19200 28438 20000 6 la1_data_in[6]
port 144 nsew signal input
rlabel metal3 s 0 16268 800 16508 6 la1_data_in[7]
port 145 nsew signal input
rlabel metal2 s 28970 19200 29082 20000 6 la1_data_in[8]
port 146 nsew signal input
rlabel metal2 s 3854 19200 3966 20000 6 la1_data_in[9]
port 147 nsew signal input
rlabel metal2 s 5786 0 5898 800 6 la1_data_out[0]
port 148 nsew signal output
rlabel metal2 s 43782 0 43894 800 6 la1_data_out[10]
port 149 nsew signal output
rlabel metal2 s 16090 0 16202 800 6 la1_data_out[11]
port 150 nsew signal output
rlabel metal3 s 49200 16948 50000 17188 6 la1_data_out[12]
port 151 nsew signal output
rlabel metal2 s 18022 19200 18134 20000 6 la1_data_out[13]
port 152 nsew signal output
rlabel metal2 s 33478 19200 33590 20000 6 la1_data_out[14]
port 153 nsew signal output
rlabel metal3 s 0 1308 800 1548 6 la1_data_out[15]
port 154 nsew signal output
rlabel metal2 s 47002 0 47114 800 6 la1_data_out[16]
port 155 nsew signal output
rlabel metal3 s 49200 10148 50000 10388 6 la1_data_out[17]
port 156 nsew signal output
rlabel metal2 s 18666 19200 18778 20000 6 la1_data_out[18]
port 157 nsew signal output
rlabel metal3 s 49200 2668 50000 2908 6 la1_data_out[19]
port 158 nsew signal output
rlabel metal2 s 10938 19200 11050 20000 6 la1_data_out[1]
port 159 nsew signal output
rlabel metal3 s 0 7428 800 7668 6 la1_data_out[20]
port 160 nsew signal output
rlabel metal3 s 49200 14908 50000 15148 6 la1_data_out[21]
port 161 nsew signal output
rlabel metal2 s 36054 19200 36166 20000 6 la1_data_out[22]
port 162 nsew signal output
rlabel metal2 s 9006 0 9118 800 6 la1_data_out[23]
port 163 nsew signal output
rlabel metal2 s 48290 0 48402 800 6 la1_data_out[24]
port 164 nsew signal output
rlabel metal3 s 0 2668 800 2908 6 la1_data_out[25]
port 165 nsew signal output
rlabel metal2 s 39274 0 39386 800 6 la1_data_out[26]
port 166 nsew signal output
rlabel metal2 s 12870 19200 12982 20000 6 la1_data_out[27]
port 167 nsew signal output
rlabel metal2 s 31546 0 31658 800 6 la1_data_out[28]
port 168 nsew signal output
rlabel metal2 s 4498 0 4610 800 6 la1_data_out[29]
port 169 nsew signal output
rlabel metal2 s 14802 0 14914 800 6 la1_data_out[2]
port 170 nsew signal output
rlabel metal2 s 44426 0 44538 800 6 la1_data_out[30]
port 171 nsew signal output
rlabel metal3 s 49200 18988 50000 19228 6 la1_data_out[31]
port 172 nsew signal output
rlabel metal3 s 0 6748 800 6988 6 la1_data_out[3]
port 173 nsew signal output
rlabel metal2 s 32190 0 32302 800 6 la1_data_out[4]
port 174 nsew signal output
rlabel metal2 s 2566 0 2678 800 6 la1_data_out[5]
port 175 nsew signal output
rlabel metal2 s 49578 0 49690 800 6 la1_data_out[6]
port 176 nsew signal output
rlabel metal2 s 634 0 746 800 6 la1_data_out[7]
port 177 nsew signal output
rlabel metal3 s 49200 10828 50000 11068 6 la1_data_out[8]
port 178 nsew signal output
rlabel metal2 s 47646 19200 47758 20000 6 la1_data_out[9]
port 179 nsew signal output
rlabel metal2 s 35410 0 35522 800 6 la1_oenb[0]
port 180 nsew signal input
rlabel metal2 s 46358 19200 46470 20000 6 la1_oenb[10]
port 181 nsew signal input
rlabel metal3 s 0 19668 800 19908 6 la1_oenb[11]
port 182 nsew signal input
rlabel metal2 s 634 19200 746 20000 6 la1_oenb[12]
port 183 nsew signal input
rlabel metal2 s 21242 0 21354 800 6 la1_oenb[13]
port 184 nsew signal input
rlabel metal2 s -10 0 102 800 6 la1_oenb[14]
port 185 nsew signal input
rlabel metal2 s 25106 0 25218 800 6 la1_oenb[15]
port 186 nsew signal input
rlabel metal2 s 4498 19200 4610 20000 6 la1_oenb[16]
port 187 nsew signal input
rlabel metal2 s 17378 19200 17490 20000 6 la1_oenb[17]
port 188 nsew signal input
rlabel metal2 s 30258 19200 30370 20000 6 la1_oenb[18]
port 189 nsew signal input
rlabel metal3 s 0 18988 800 19228 6 la1_oenb[19]
port 190 nsew signal input
rlabel metal2 s 6430 0 6542 800 6 la1_oenb[1]
port 191 nsew signal input
rlabel metal2 s 1922 0 2034 800 6 la1_oenb[20]
port 192 nsew signal input
rlabel metal2 s 37342 19200 37454 20000 6 la1_oenb[21]
port 193 nsew signal input
rlabel metal2 s 29614 19200 29726 20000 6 la1_oenb[22]
port 194 nsew signal input
rlabel metal2 s 17378 0 17490 800 6 la1_oenb[23]
port 195 nsew signal input
rlabel metal2 s 42494 19200 42606 20000 6 la1_oenb[24]
port 196 nsew signal input
rlabel metal2 s 42494 0 42606 800 6 la1_oenb[25]
port 197 nsew signal input
rlabel metal2 s 7074 19200 7186 20000 6 la1_oenb[26]
port 198 nsew signal input
rlabel metal3 s 49200 9468 50000 9708 6 la1_oenb[27]
port 199 nsew signal input
rlabel metal2 s 7074 0 7186 800 6 la1_oenb[28]
port 200 nsew signal input
rlabel metal2 s 12870 0 12982 800 6 la1_oenb[29]
port 201 nsew signal input
rlabel metal3 s 0 6068 800 6308 6 la1_oenb[2]
port 202 nsew signal input
rlabel metal3 s 49200 8788 50000 9028 6 la1_oenb[30]
port 203 nsew signal input
rlabel metal2 s 19954 0 20066 800 6 la1_oenb[31]
port 204 nsew signal input
rlabel metal2 s 39274 19200 39386 20000 6 la1_oenb[3]
port 205 nsew signal input
rlabel metal2 s 38630 19200 38742 20000 6 la1_oenb[4]
port 206 nsew signal input
rlabel metal2 s 13514 19200 13626 20000 6 la1_oenb[5]
port 207 nsew signal input
rlabel metal2 s 19954 19200 20066 20000 6 la1_oenb[6]
port 208 nsew signal input
rlabel metal2 s 24462 0 24574 800 6 la1_oenb[7]
port 209 nsew signal input
rlabel metal3 s 0 8788 800 9028 6 la1_oenb[8]
port 210 nsew signal input
rlabel metal2 s 9006 19200 9118 20000 6 la1_oenb[9]
port 211 nsew signal input
rlabel metal4 s 8910 2128 9230 17456 6 vccd1
port 212 nsew power input
rlabel metal4 s 24840 2128 25160 17456 6 vccd1
port 212 nsew power input
rlabel metal4 s 40771 2128 41091 17456 6 vccd1
port 212 nsew power input
rlabel metal4 s 16874 2128 17194 17456 6 vssd1
port 213 nsew ground input
rlabel metal4 s 32805 2128 33125 17456 6 vssd1
port 213 nsew ground input
rlabel metal3 s 49200 1308 50000 1548 6 wb_clk_i
port 214 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 50000 20000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 787908
string GDS_FILE /openlane/designs/wrapped_frequency_counter/runs/RUN_2022.03.16_16.36.24/results/finishing/wrapped_frequency_counter.magic.gds
string GDS_START 88388
<< end >>

