// This is the unpowered netlist.
module wrapped_frequency_counter (active,
    wb_clk_i,
    io_in,
    io_oeb,
    io_out,
    la1_data_in,
    la1_data_out,
    la1_oenb);
 input active;
 input wb_clk_i;
 input [37:0] io_in;
 output [37:0] io_oeb;
 output [37:0] io_out;
 input [31:0] la1_data_in;
 output [31:0] la1_data_out;
 input [31:0] la1_oenb;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire clknet_0_wb_clk_i;
 wire \frequency_counter_0.clk_counter[0] ;
 wire \frequency_counter_0.clk_counter[10] ;
 wire \frequency_counter_0.clk_counter[11] ;
 wire \frequency_counter_0.clk_counter[1] ;
 wire \frequency_counter_0.clk_counter[2] ;
 wire \frequency_counter_0.clk_counter[3] ;
 wire \frequency_counter_0.clk_counter[4] ;
 wire \frequency_counter_0.clk_counter[5] ;
 wire \frequency_counter_0.clk_counter[6] ;
 wire \frequency_counter_0.clk_counter[7] ;
 wire \frequency_counter_0.clk_counter[8] ;
 wire \frequency_counter_0.clk_counter[9] ;
 wire \frequency_counter_0.dbg_edge_count[0] ;
 wire \frequency_counter_0.dbg_edge_count[1] ;
 wire \frequency_counter_0.dbg_edge_count[2] ;
 wire \frequency_counter_0.dbg_state[0] ;
 wire \frequency_counter_0.dbg_state[1] ;
 wire \frequency_counter_0.digit ;
 wire \frequency_counter_0.edge_counter[0] ;
 wire \frequency_counter_0.edge_counter[1] ;
 wire \frequency_counter_0.edge_counter[2] ;
 wire \frequency_counter_0.edge_counter[3] ;
 wire \frequency_counter_0.edge_detect0.q0 ;
 wire \frequency_counter_0.edge_detect0.q1 ;
 wire \frequency_counter_0.edge_detect0.q2 ;
 wire \frequency_counter_0.segments[0] ;
 wire \frequency_counter_0.segments[1] ;
 wire \frequency_counter_0.segments[2] ;
 wire \frequency_counter_0.segments[3] ;
 wire \frequency_counter_0.segments[4] ;
 wire \frequency_counter_0.segments[5] ;
 wire \frequency_counter_0.segments[6] ;
 wire \frequency_counter_0.seven_segment0.load ;
 wire \frequency_counter_0.seven_segment0.ten_count[0] ;
 wire \frequency_counter_0.seven_segment0.ten_count[1] ;
 wire \frequency_counter_0.seven_segment0.ten_count[2] ;
 wire \frequency_counter_0.seven_segment0.ten_count[3] ;
 wire \frequency_counter_0.seven_segment0.ten_count_reg[0] ;
 wire \frequency_counter_0.seven_segment0.ten_count_reg[1] ;
 wire \frequency_counter_0.seven_segment0.ten_count_reg[2] ;
 wire \frequency_counter_0.seven_segment0.ten_count_reg[3] ;
 wire \frequency_counter_0.seven_segment0.unit_count[0] ;
 wire \frequency_counter_0.seven_segment0.unit_count[1] ;
 wire \frequency_counter_0.seven_segment0.unit_count[2] ;
 wire \frequency_counter_0.seven_segment0.unit_count[3] ;
 wire \frequency_counter_0.seven_segment0.unit_count_reg[0] ;
 wire \frequency_counter_0.seven_segment0.unit_count_reg[1] ;
 wire \frequency_counter_0.seven_segment0.unit_count_reg[2] ;
 wire \frequency_counter_0.seven_segment0.unit_count_reg[3] ;
 wire \frequency_counter_0.update_period[0] ;
 wire \frequency_counter_0.update_period[10] ;
 wire \frequency_counter_0.update_period[11] ;
 wire \frequency_counter_0.update_period[1] ;
 wire \frequency_counter_0.update_period[2] ;
 wire \frequency_counter_0.update_period[3] ;
 wire \frequency_counter_0.update_period[4] ;
 wire \frequency_counter_0.update_period[5] ;
 wire \frequency_counter_0.update_period[6] ;
 wire \frequency_counter_0.update_period[7] ;
 wire \frequency_counter_0.update_period[8] ;
 wire \frequency_counter_0.update_period[9] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire clknet_2_0__leaf_wb_clk_i;
 wire clknet_2_1__leaf_wb_clk_i;
 wire clknet_2_2__leaf_wb_clk_i;
 wire clknet_2_3__leaf_wb_clk_i;
 wire net108;
 wire net109;

 sky130_fd_sc_hd__clkbuf_8 _0470_ (.A(net1),
    .X(_0051_));
 sky130_fd_sc_hd__buf_8 _0471_ (.A(_0051_),
    .X(_0052_));
 sky130_fd_sc_hd__buf_6 _0472_ (.A(_0052_),
    .X(_0053_));
 sky130_fd_sc_hd__inv_2 _0473_ (.A(_0053_),
    .Y(_0378_));
 sky130_fd_sc_hd__inv_2 _0474_ (.A(_0053_),
    .Y(_0377_));
 sky130_fd_sc_hd__inv_2 _0475_ (.A(_0053_),
    .Y(_0376_));
 sky130_fd_sc_hd__inv_2 _0476_ (.A(_0053_),
    .Y(_0375_));
 sky130_fd_sc_hd__inv_2 _0477_ (.A(_0053_),
    .Y(_0374_));
 sky130_fd_sc_hd__inv_2 _0478_ (.A(_0053_),
    .Y(_0373_));
 sky130_fd_sc_hd__inv_2 _0479_ (.A(_0053_),
    .Y(_0372_));
 sky130_fd_sc_hd__inv_2 _0480_ (.A(_0053_),
    .Y(_0371_));
 sky130_fd_sc_hd__inv_2 _0481_ (.A(_0053_),
    .Y(_0370_));
 sky130_fd_sc_hd__inv_2 _0482_ (.A(_0053_),
    .Y(_0369_));
 sky130_fd_sc_hd__buf_8 _0483_ (.A(_0052_),
    .X(_0054_));
 sky130_fd_sc_hd__inv_2 _0484_ (.A(_0054_),
    .Y(_0368_));
 sky130_fd_sc_hd__inv_2 _0485_ (.A(_0054_),
    .Y(_0367_));
 sky130_fd_sc_hd__inv_2 _0486_ (.A(_0054_),
    .Y(_0366_));
 sky130_fd_sc_hd__inv_2 _0487_ (.A(_0054_),
    .Y(_0365_));
 sky130_fd_sc_hd__inv_2 _0488_ (.A(_0054_),
    .Y(_0364_));
 sky130_fd_sc_hd__inv_2 _0489_ (.A(_0054_),
    .Y(_0363_));
 sky130_fd_sc_hd__inv_2 _0490_ (.A(_0054_),
    .Y(_0362_));
 sky130_fd_sc_hd__inv_2 _0491_ (.A(_0054_),
    .Y(_0361_));
 sky130_fd_sc_hd__inv_2 _0492_ (.A(_0054_),
    .Y(_0360_));
 sky130_fd_sc_hd__inv_2 _0493_ (.A(_0054_),
    .Y(_0359_));
 sky130_fd_sc_hd__buf_8 _0494_ (.A(_0051_),
    .X(_0055_));
 sky130_fd_sc_hd__inv_2 _0495_ (.A(_0055_),
    .Y(_0358_));
 sky130_fd_sc_hd__inv_2 _0496_ (.A(_0055_),
    .Y(_0357_));
 sky130_fd_sc_hd__inv_2 _0497_ (.A(_0055_),
    .Y(_0356_));
 sky130_fd_sc_hd__inv_2 _0498_ (.A(_0055_),
    .Y(_0355_));
 sky130_fd_sc_hd__inv_2 _0499_ (.A(_0055_),
    .Y(_0354_));
 sky130_fd_sc_hd__inv_2 _0500_ (.A(_0055_),
    .Y(_0353_));
 sky130_fd_sc_hd__inv_2 _0501_ (.A(_0055_),
    .Y(_0352_));
 sky130_fd_sc_hd__inv_2 _0502_ (.A(_0055_),
    .Y(_0351_));
 sky130_fd_sc_hd__inv_2 _0503_ (.A(_0055_),
    .Y(_0339_));
 sky130_fd_sc_hd__inv_2 _0504_ (.A(_0055_),
    .Y(_0340_));
 sky130_fd_sc_hd__buf_8 _0505_ (.A(_0051_),
    .X(_0056_));
 sky130_fd_sc_hd__inv_2 _0506_ (.A(_0056_),
    .Y(_0342_));
 sky130_fd_sc_hd__inv_2 _0507_ (.A(_0056_),
    .Y(_0343_));
 sky130_fd_sc_hd__inv_2 _0508_ (.A(_0056_),
    .Y(_0344_));
 sky130_fd_sc_hd__inv_2 _0509_ (.A(_0056_),
    .Y(_0345_));
 sky130_fd_sc_hd__inv_2 _0510_ (.A(_0056_),
    .Y(_0346_));
 sky130_fd_sc_hd__inv_2 _0511_ (.A(_0056_),
    .Y(_0347_));
 sky130_fd_sc_hd__inv_2 _0512_ (.A(_0056_),
    .Y(_0348_));
 sky130_fd_sc_hd__inv_2 _0513_ (.A(_0056_),
    .Y(_0349_));
 sky130_fd_sc_hd__inv_2 _0514_ (.A(_0056_),
    .Y(_0290_));
 sky130_fd_sc_hd__inv_2 _0515_ (.A(_0056_),
    .Y(_0297_));
 sky130_fd_sc_hd__buf_8 _0516_ (.A(_0051_),
    .X(_0057_));
 sky130_fd_sc_hd__inv_2 _0517_ (.A(_0057_),
    .Y(_0301_));
 sky130_fd_sc_hd__inv_2 _0518_ (.A(_0057_),
    .Y(_0325_));
 sky130_fd_sc_hd__inv_2 _0519_ (.A(_0057_),
    .Y(_0326_));
 sky130_fd_sc_hd__inv_2 _0520_ (.A(_0057_),
    .Y(_0327_));
 sky130_fd_sc_hd__inv_2 _0521_ (.A(_0057_),
    .Y(_0271_));
 sky130_fd_sc_hd__inv_2 _0522_ (.A(_0057_),
    .Y(_0272_));
 sky130_fd_sc_hd__inv_2 _0523_ (.A(_0057_),
    .Y(_0273_));
 sky130_fd_sc_hd__inv_2 _0524_ (.A(_0057_),
    .Y(_0274_));
 sky130_fd_sc_hd__inv_2 _0525_ (.A(_0057_),
    .Y(_0275_));
 sky130_fd_sc_hd__inv_2 _0526_ (.A(_0057_),
    .Y(_0276_));
 sky130_fd_sc_hd__buf_8 _0527_ (.A(_0051_),
    .X(_0058_));
 sky130_fd_sc_hd__inv_2 _0528_ (.A(_0058_),
    .Y(_0277_));
 sky130_fd_sc_hd__inv_2 _0529_ (.A(_0058_),
    .Y(_0278_));
 sky130_fd_sc_hd__inv_2 _0530_ (.A(_0058_),
    .Y(_0279_));
 sky130_fd_sc_hd__inv_2 _0531_ (.A(_0058_),
    .Y(_0280_));
 sky130_fd_sc_hd__inv_2 _0532_ (.A(_0058_),
    .Y(_0281_));
 sky130_fd_sc_hd__inv_2 _0533_ (.A(_0058_),
    .Y(_0282_));
 sky130_fd_sc_hd__inv_2 _0534_ (.A(_0058_),
    .Y(_0283_));
 sky130_fd_sc_hd__inv_2 _0535_ (.A(_0058_),
    .Y(_0284_));
 sky130_fd_sc_hd__inv_2 _0536_ (.A(_0058_),
    .Y(_0285_));
 sky130_fd_sc_hd__inv_2 _0537_ (.A(_0058_),
    .Y(_0286_));
 sky130_fd_sc_hd__buf_8 _0538_ (.A(_0051_),
    .X(_0059_));
 sky130_fd_sc_hd__inv_2 _0539_ (.A(_0059_),
    .Y(_0287_));
 sky130_fd_sc_hd__inv_2 _0540_ (.A(_0059_),
    .Y(_0288_));
 sky130_fd_sc_hd__inv_2 _0541_ (.A(_0059_),
    .Y(_0289_));
 sky130_fd_sc_hd__inv_2 _0542_ (.A(_0059_),
    .Y(_0328_));
 sky130_fd_sc_hd__inv_2 _0543_ (.A(_0059_),
    .Y(_0302_));
 sky130_fd_sc_hd__inv_2 _0544_ (.A(_0059_),
    .Y(_0304_));
 sky130_fd_sc_hd__inv_2 _0545_ (.A(_0059_),
    .Y(_0329_));
 sky130_fd_sc_hd__inv_2 _0546_ (.A(_0059_),
    .Y(_0305_));
 sky130_fd_sc_hd__inv_2 _0547_ (.A(_0059_),
    .Y(_0306_));
 sky130_fd_sc_hd__inv_2 _0548_ (.A(_0059_),
    .Y(_0330_));
 sky130_fd_sc_hd__buf_8 _0549_ (.A(_0051_),
    .X(_0060_));
 sky130_fd_sc_hd__inv_2 _0550_ (.A(_0060_),
    .Y(_0307_));
 sky130_fd_sc_hd__inv_2 _0551_ (.A(_0060_),
    .Y(_0308_));
 sky130_fd_sc_hd__inv_2 _0552_ (.A(_0060_),
    .Y(_0331_));
 sky130_fd_sc_hd__inv_2 _0553_ (.A(_0060_),
    .Y(_0309_));
 sky130_fd_sc_hd__inv_2 _0554_ (.A(_0060_),
    .Y(_0310_));
 sky130_fd_sc_hd__inv_2 _0555_ (.A(_0060_),
    .Y(_0332_));
 sky130_fd_sc_hd__inv_2 _0556_ (.A(_0060_),
    .Y(_0311_));
 sky130_fd_sc_hd__inv_2 _0557_ (.A(_0060_),
    .Y(_0312_));
 sky130_fd_sc_hd__inv_2 _0558_ (.A(_0060_),
    .Y(_0333_));
 sky130_fd_sc_hd__inv_2 _0559_ (.A(_0060_),
    .Y(_0334_));
 sky130_fd_sc_hd__buf_6 _0560_ (.A(_0051_),
    .X(_0061_));
 sky130_fd_sc_hd__inv_2 _0561_ (.A(_0061_),
    .Y(_0338_));
 sky130_fd_sc_hd__inv_2 _0562_ (.A(_0061_),
    .Y(_0313_));
 sky130_fd_sc_hd__inv_2 _0563_ (.A(_0061_),
    .Y(_0314_));
 sky130_fd_sc_hd__inv_2 _0564_ (.A(_0061_),
    .Y(_0315_));
 sky130_fd_sc_hd__inv_2 _0565_ (.A(_0061_),
    .Y(_0316_));
 sky130_fd_sc_hd__inv_2 _0566_ (.A(_0061_),
    .Y(_0335_));
 sky130_fd_sc_hd__inv_2 _0567_ (.A(_0061_),
    .Y(_0317_));
 sky130_fd_sc_hd__inv_2 _0568_ (.A(_0061_),
    .Y(_0336_));
 sky130_fd_sc_hd__inv_2 _0569_ (.A(_0061_),
    .Y(_0318_));
 sky130_fd_sc_hd__inv_2 _0570_ (.A(_0061_),
    .Y(_0319_));
 sky130_fd_sc_hd__buf_8 _0571_ (.A(_0051_),
    .X(_0062_));
 sky130_fd_sc_hd__inv_2 _0572_ (.A(_0062_),
    .Y(_0320_));
 sky130_fd_sc_hd__inv_2 _0573_ (.A(_0062_),
    .Y(_0321_));
 sky130_fd_sc_hd__inv_2 _0574_ (.A(_0062_),
    .Y(_0322_));
 sky130_fd_sc_hd__inv_2 _0575_ (.A(_0062_),
    .Y(_0323_));
 sky130_fd_sc_hd__inv_2 _0576_ (.A(_0062_),
    .Y(_0324_));
 sky130_fd_sc_hd__inv_2 _0577_ (.A(_0062_),
    .Y(_0337_));
 sky130_fd_sc_hd__inv_2 _0578_ (.A(_0062_),
    .Y(_0291_));
 sky130_fd_sc_hd__inv_2 _0579_ (.A(_0062_),
    .Y(_0292_));
 sky130_fd_sc_hd__inv_2 _0580_ (.A(_0062_),
    .Y(_0293_));
 sky130_fd_sc_hd__inv_2 _0581_ (.A(_0062_),
    .Y(_0294_));
 sky130_fd_sc_hd__inv_2 _0582_ (.A(_0052_),
    .Y(_0295_));
 sky130_fd_sc_hd__inv_2 _0583_ (.A(_0052_),
    .Y(_0296_));
 sky130_fd_sc_hd__inv_2 _0584_ (.A(_0052_),
    .Y(_0299_));
 sky130_fd_sc_hd__inv_2 _0585_ (.A(_0052_),
    .Y(_0300_));
 sky130_fd_sc_hd__inv_2 _0586_ (.A(_0052_),
    .Y(_0298_));
 sky130_fd_sc_hd__inv_2 _0587_ (.A(_0052_),
    .Y(_0350_));
 sky130_fd_sc_hd__inv_2 _0588_ (.A(_0052_),
    .Y(_0341_));
 sky130_fd_sc_hd__inv_2 _0589_ (.A(_0052_),
    .Y(_0303_));
 sky130_fd_sc_hd__mux2_2 _0590_ (.A0(\frequency_counter_0.seven_segment0.unit_count_reg[3] ),
    .A1(\frequency_counter_0.seven_segment0.ten_count_reg[3] ),
    .S(\frequency_counter_0.digit ),
    .X(_0063_));
 sky130_fd_sc_hd__inv_2 _0591_ (.A(_0063_),
    .Y(_0064_));
 sky130_fd_sc_hd__mux2_1 _0592_ (.A0(\frequency_counter_0.seven_segment0.unit_count_reg[2] ),
    .A1(\frequency_counter_0.seven_segment0.ten_count_reg[2] ),
    .S(\frequency_counter_0.digit ),
    .X(_0065_));
 sky130_fd_sc_hd__mux2_2 _0593_ (.A0(\frequency_counter_0.seven_segment0.unit_count_reg[0] ),
    .A1(\frequency_counter_0.seven_segment0.ten_count_reg[0] ),
    .S(\frequency_counter_0.digit ),
    .X(_0066_));
 sky130_fd_sc_hd__nor2_1 _0594_ (.A(_0065_),
    .B(_0066_),
    .Y(_0067_));
 sky130_fd_sc_hd__mux2_2 _0595_ (.A0(\frequency_counter_0.seven_segment0.unit_count_reg[1] ),
    .A1(\frequency_counter_0.seven_segment0.ten_count_reg[1] ),
    .S(\frequency_counter_0.digit ),
    .X(_0068_));
 sky130_fd_sc_hd__nor2_1 _0596_ (.A(_0065_),
    .B(_0068_),
    .Y(_0069_));
 sky130_fd_sc_hd__nor2_1 _0597_ (.A(_0069_),
    .B(_0063_),
    .Y(_0070_));
 sky130_fd_sc_hd__and2_1 _0598_ (.A(_0069_),
    .B(_0063_),
    .X(_0071_));
 sky130_fd_sc_hd__a221o_1 _0599_ (.A1(_0064_),
    .A2(_0067_),
    .B1(_0070_),
    .B2(_0066_),
    .C1(_0071_),
    .X(\frequency_counter_0.segments[0] ));
 sky130_fd_sc_hd__a21bo_1 _0600_ (.A1(_0068_),
    .A2(_0066_),
    .B1_N(_0065_),
    .X(_0072_));
 sky130_fd_sc_hd__or2_1 _0601_ (.A(_0068_),
    .B(_0066_),
    .X(_0073_));
 sky130_fd_sc_hd__or2b_1 _0602_ (.A(_0072_),
    .B_N(_0073_),
    .X(_0074_));
 sky130_fd_sc_hd__a21o_1 _0603_ (.A1(_0064_),
    .A2(_0074_),
    .B1(_0071_),
    .X(\frequency_counter_0.segments[1] ));
 sky130_fd_sc_hd__o21bai_1 _0604_ (.A1(_0063_),
    .A2(_0067_),
    .B1_N(_0069_),
    .Y(\frequency_counter_0.segments[2] ));
 sky130_fd_sc_hd__nand2_1 _0605_ (.A(_0065_),
    .B(_0068_),
    .Y(_0075_));
 sky130_fd_sc_hd__a21oi_1 _0606_ (.A1(_0068_),
    .A2(_0064_),
    .B1(_0069_),
    .Y(_0076_));
 sky130_fd_sc_hd__nor2_1 _0607_ (.A(_0066_),
    .B(_0076_),
    .Y(\frequency_counter_0.segments[4] ));
 sky130_fd_sc_hd__a31o_1 _0608_ (.A1(_0070_),
    .A2(_0073_),
    .A3(_0075_),
    .B1(\frequency_counter_0.segments[4] ),
    .X(\frequency_counter_0.segments[3] ));
 sky130_fd_sc_hd__a21oi_1 _0609_ (.A1(_0072_),
    .A2(_0073_),
    .B1(_0063_),
    .Y(_0077_));
 sky130_fd_sc_hd__or2_1 _0610_ (.A(_0071_),
    .B(_0077_),
    .X(_0078_));
 sky130_fd_sc_hd__clkbuf_1 _0611_ (.A(_0078_),
    .X(\frequency_counter_0.segments[5] ));
 sky130_fd_sc_hd__nand3_1 _0612_ (.A(_0065_),
    .B(_0068_),
    .C(_0066_),
    .Y(_0079_));
 sky130_fd_sc_hd__a21o_1 _0613_ (.A1(_0070_),
    .A2(_0079_),
    .B1(_0071_),
    .X(\frequency_counter_0.segments[6] ));
 sky130_fd_sc_hd__clkbuf_4 _0614_ (.A(net3),
    .X(_0080_));
 sky130_fd_sc_hd__clkbuf_4 _0615_ (.A(_0080_),
    .X(_0081_));
 sky130_fd_sc_hd__nor2_1 _0616_ (.A(\frequency_counter_0.digit ),
    .B(_0081_),
    .Y(_0000_));
 sky130_fd_sc_hd__inv_2 _0617_ (.A(net3),
    .Y(_0082_));
 sky130_fd_sc_hd__buf_2 _0618_ (.A(_0082_),
    .X(_0083_));
 sky130_fd_sc_hd__mux2_1 _0619_ (.A0(\frequency_counter_0.seven_segment0.ten_count_reg[0] ),
    .A1(\frequency_counter_0.seven_segment0.ten_count[0] ),
    .S(\frequency_counter_0.seven_segment0.load ),
    .X(_0084_));
 sky130_fd_sc_hd__and2_1 _0620_ (.A(_0083_),
    .B(_0084_),
    .X(_0085_));
 sky130_fd_sc_hd__clkbuf_1 _0621_ (.A(_0085_),
    .X(_0001_));
 sky130_fd_sc_hd__buf_2 _0622_ (.A(_0082_),
    .X(_0086_));
 sky130_fd_sc_hd__mux2_1 _0623_ (.A0(\frequency_counter_0.seven_segment0.ten_count_reg[1] ),
    .A1(\frequency_counter_0.seven_segment0.ten_count[1] ),
    .S(\frequency_counter_0.seven_segment0.load ),
    .X(_0087_));
 sky130_fd_sc_hd__and2_1 _0624_ (.A(_0086_),
    .B(_0087_),
    .X(_0088_));
 sky130_fd_sc_hd__clkbuf_1 _0625_ (.A(_0088_),
    .X(_0002_));
 sky130_fd_sc_hd__mux2_1 _0626_ (.A0(\frequency_counter_0.seven_segment0.ten_count_reg[2] ),
    .A1(\frequency_counter_0.seven_segment0.ten_count[2] ),
    .S(\frequency_counter_0.seven_segment0.load ),
    .X(_0089_));
 sky130_fd_sc_hd__and2_1 _0627_ (.A(_0086_),
    .B(_0089_),
    .X(_0090_));
 sky130_fd_sc_hd__clkbuf_1 _0628_ (.A(_0090_),
    .X(_0003_));
 sky130_fd_sc_hd__mux2_1 _0629_ (.A0(\frequency_counter_0.seven_segment0.ten_count_reg[3] ),
    .A1(\frequency_counter_0.seven_segment0.ten_count[3] ),
    .S(\frequency_counter_0.seven_segment0.load ),
    .X(_0091_));
 sky130_fd_sc_hd__and2_1 _0630_ (.A(_0086_),
    .B(_0091_),
    .X(_0092_));
 sky130_fd_sc_hd__clkbuf_1 _0631_ (.A(_0092_),
    .X(_0004_));
 sky130_fd_sc_hd__mux2_1 _0632_ (.A0(\frequency_counter_0.seven_segment0.unit_count_reg[0] ),
    .A1(\frequency_counter_0.seven_segment0.unit_count[0] ),
    .S(\frequency_counter_0.seven_segment0.load ),
    .X(_0093_));
 sky130_fd_sc_hd__and2_1 _0633_ (.A(_0086_),
    .B(_0093_),
    .X(_0094_));
 sky130_fd_sc_hd__clkbuf_1 _0634_ (.A(_0094_),
    .X(_0005_));
 sky130_fd_sc_hd__mux2_1 _0635_ (.A0(\frequency_counter_0.seven_segment0.unit_count_reg[1] ),
    .A1(\frequency_counter_0.seven_segment0.unit_count[1] ),
    .S(\frequency_counter_0.seven_segment0.load ),
    .X(_0095_));
 sky130_fd_sc_hd__and2_1 _0636_ (.A(_0086_),
    .B(_0095_),
    .X(_0096_));
 sky130_fd_sc_hd__clkbuf_1 _0637_ (.A(_0096_),
    .X(_0006_));
 sky130_fd_sc_hd__mux2_1 _0638_ (.A0(\frequency_counter_0.seven_segment0.unit_count_reg[2] ),
    .A1(\frequency_counter_0.seven_segment0.unit_count[2] ),
    .S(\frequency_counter_0.seven_segment0.load ),
    .X(_0097_));
 sky130_fd_sc_hd__and2_1 _0639_ (.A(_0086_),
    .B(_0097_),
    .X(_0098_));
 sky130_fd_sc_hd__clkbuf_1 _0640_ (.A(_0098_),
    .X(_0007_));
 sky130_fd_sc_hd__mux2_1 _0641_ (.A0(\frequency_counter_0.seven_segment0.unit_count_reg[3] ),
    .A1(\frequency_counter_0.seven_segment0.unit_count[3] ),
    .S(\frequency_counter_0.seven_segment0.load ),
    .X(_0099_));
 sky130_fd_sc_hd__and2_1 _0642_ (.A(_0086_),
    .B(_0099_),
    .X(_0100_));
 sky130_fd_sc_hd__clkbuf_1 _0643_ (.A(_0100_),
    .X(_0008_));
 sky130_fd_sc_hd__clkbuf_4 _0644_ (.A(_0080_),
    .X(_0101_));
 sky130_fd_sc_hd__buf_4 _0645_ (.A(net8),
    .X(_0102_));
 sky130_fd_sc_hd__mux2_1 _0646_ (.A0(\frequency_counter_0.update_period[0] ),
    .A1(net9),
    .S(_0102_),
    .X(_0103_));
 sky130_fd_sc_hd__or2_1 _0647_ (.A(_0101_),
    .B(_0103_),
    .X(_0104_));
 sky130_fd_sc_hd__clkbuf_1 _0648_ (.A(_0104_),
    .X(_0009_));
 sky130_fd_sc_hd__mux2_1 _0649_ (.A0(\frequency_counter_0.update_period[1] ),
    .A1(net10),
    .S(_0102_),
    .X(_0105_));
 sky130_fd_sc_hd__or2_1 _0650_ (.A(_0101_),
    .B(_0105_),
    .X(_0106_));
 sky130_fd_sc_hd__clkbuf_1 _0651_ (.A(_0106_),
    .X(_0010_));
 sky130_fd_sc_hd__mux2_1 _0652_ (.A0(\frequency_counter_0.update_period[2] ),
    .A1(net11),
    .S(_0102_),
    .X(_0107_));
 sky130_fd_sc_hd__or2_1 _0653_ (.A(_0080_),
    .B(_0107_),
    .X(_0108_));
 sky130_fd_sc_hd__clkbuf_1 _0654_ (.A(_0108_),
    .X(_0011_));
 sky130_fd_sc_hd__mux2_1 _0655_ (.A0(\frequency_counter_0.update_period[3] ),
    .A1(net12),
    .S(_0102_),
    .X(_0109_));
 sky130_fd_sc_hd__or2_1 _0656_ (.A(_0080_),
    .B(_0109_),
    .X(_0110_));
 sky130_fd_sc_hd__clkbuf_1 _0657_ (.A(_0110_),
    .X(_0012_));
 sky130_fd_sc_hd__mux2_1 _0658_ (.A0(\frequency_counter_0.update_period[4] ),
    .A1(net13),
    .S(_0102_),
    .X(_0111_));
 sky130_fd_sc_hd__and2_1 _0659_ (.A(_0086_),
    .B(_0111_),
    .X(_0112_));
 sky130_fd_sc_hd__clkbuf_1 _0660_ (.A(_0112_),
    .X(_0013_));
 sky130_fd_sc_hd__mux2_1 _0661_ (.A0(\frequency_counter_0.update_period[5] ),
    .A1(net14),
    .S(_0102_),
    .X(_0113_));
 sky130_fd_sc_hd__or2_1 _0662_ (.A(_0080_),
    .B(_0113_),
    .X(_0114_));
 sky130_fd_sc_hd__clkbuf_1 _0663_ (.A(_0114_),
    .X(_0014_));
 sky130_fd_sc_hd__mux2_1 _0664_ (.A0(\frequency_counter_0.update_period[6] ),
    .A1(net15),
    .S(_0102_),
    .X(_0115_));
 sky130_fd_sc_hd__and2_1 _0665_ (.A(_0086_),
    .B(_0115_),
    .X(_0116_));
 sky130_fd_sc_hd__clkbuf_1 _0666_ (.A(_0116_),
    .X(_0015_));
 sky130_fd_sc_hd__mux2_1 _0667_ (.A0(\frequency_counter_0.update_period[7] ),
    .A1(net16),
    .S(net8),
    .X(_0117_));
 sky130_fd_sc_hd__or2_1 _0668_ (.A(_0080_),
    .B(_0117_),
    .X(_0118_));
 sky130_fd_sc_hd__clkbuf_1 _0669_ (.A(_0118_),
    .X(_0016_));
 sky130_fd_sc_hd__mux2_1 _0670_ (.A0(\frequency_counter_0.update_period[8] ),
    .A1(net4),
    .S(_0102_),
    .X(_0119_));
 sky130_fd_sc_hd__and2_1 _0671_ (.A(_0086_),
    .B(_0119_),
    .X(_0120_));
 sky130_fd_sc_hd__clkbuf_1 _0672_ (.A(_0120_),
    .X(_0017_));
 sky130_fd_sc_hd__mux2_1 _0673_ (.A0(\frequency_counter_0.update_period[9] ),
    .A1(net5),
    .S(_0102_),
    .X(_0121_));
 sky130_fd_sc_hd__and2_1 _0674_ (.A(_0082_),
    .B(_0121_),
    .X(_0122_));
 sky130_fd_sc_hd__clkbuf_1 _0675_ (.A(_0122_),
    .X(_0018_));
 sky130_fd_sc_hd__mux2_1 _0676_ (.A0(\frequency_counter_0.update_period[10] ),
    .A1(net6),
    .S(net8),
    .X(_0123_));
 sky130_fd_sc_hd__or2_1 _0677_ (.A(_0080_),
    .B(_0123_),
    .X(_0124_));
 sky130_fd_sc_hd__clkbuf_1 _0678_ (.A(_0124_),
    .X(_0019_));
 sky130_fd_sc_hd__mux2_1 _0679_ (.A0(\frequency_counter_0.update_period[11] ),
    .A1(net7),
    .S(_0102_),
    .X(_0125_));
 sky130_fd_sc_hd__and2_1 _0680_ (.A(_0082_),
    .B(_0125_),
    .X(_0126_));
 sky130_fd_sc_hd__clkbuf_1 _0681_ (.A(_0126_),
    .X(_0020_));
 sky130_fd_sc_hd__inv_2 _0682_ (.A(\frequency_counter_0.clk_counter[10] ),
    .Y(_0127_));
 sky130_fd_sc_hd__inv_2 _0683_ (.A(\frequency_counter_0.update_period[11] ),
    .Y(_0128_));
 sky130_fd_sc_hd__a2bb2o_1 _0684_ (.A1_N(\frequency_counter_0.update_period[10] ),
    .A2_N(_0127_),
    .B1(\frequency_counter_0.clk_counter[11] ),
    .B2(_0128_),
    .X(_0129_));
 sky130_fd_sc_hd__or2_1 _0685_ (.A(\frequency_counter_0.clk_counter[11] ),
    .B(_0128_),
    .X(_0130_));
 sky130_fd_sc_hd__or2_1 _0686_ (.A(\frequency_counter_0.dbg_state[1] ),
    .B(\frequency_counter_0.dbg_state[0] ),
    .X(_0131_));
 sky130_fd_sc_hd__a21oi_1 _0687_ (.A1(_0129_),
    .A2(_0130_),
    .B1(_0131_),
    .Y(_0132_));
 sky130_fd_sc_hd__inv_2 _0688_ (.A(\frequency_counter_0.clk_counter[6] ),
    .Y(_0133_));
 sky130_fd_sc_hd__inv_2 _0689_ (.A(\frequency_counter_0.clk_counter[5] ),
    .Y(_0134_));
 sky130_fd_sc_hd__a22oi_1 _0690_ (.A1(_0133_),
    .A2(\frequency_counter_0.update_period[6] ),
    .B1(\frequency_counter_0.update_period[5] ),
    .B2(_0134_),
    .Y(_0135_));
 sky130_fd_sc_hd__inv_2 _0691_ (.A(\frequency_counter_0.clk_counter[1] ),
    .Y(_0136_));
 sky130_fd_sc_hd__inv_2 _0692_ (.A(\frequency_counter_0.clk_counter[0] ),
    .Y(_0137_));
 sky130_fd_sc_hd__o211a_1 _0693_ (.A1(_0136_),
    .A2(\frequency_counter_0.update_period[1] ),
    .B1(\frequency_counter_0.update_period[0] ),
    .C1(_0137_),
    .X(_0138_));
 sky130_fd_sc_hd__inv_2 _0694_ (.A(\frequency_counter_0.clk_counter[2] ),
    .Y(_0139_));
 sky130_fd_sc_hd__a22o_1 _0695_ (.A1(_0139_),
    .A2(\frequency_counter_0.update_period[2] ),
    .B1(\frequency_counter_0.update_period[1] ),
    .B2(_0136_),
    .X(_0140_));
 sky130_fd_sc_hd__inv_2 _0696_ (.A(\frequency_counter_0.clk_counter[3] ),
    .Y(_0141_));
 sky130_fd_sc_hd__o22a_1 _0697_ (.A1(_0141_),
    .A2(\frequency_counter_0.update_period[3] ),
    .B1(\frequency_counter_0.update_period[2] ),
    .B2(_0139_),
    .X(_0142_));
 sky130_fd_sc_hd__o21ai_1 _0698_ (.A1(_0138_),
    .A2(_0140_),
    .B1(_0142_),
    .Y(_0143_));
 sky130_fd_sc_hd__inv_2 _0699_ (.A(\frequency_counter_0.clk_counter[7] ),
    .Y(_0144_));
 sky130_fd_sc_hd__o22a_1 _0700_ (.A1(_0144_),
    .A2(\frequency_counter_0.update_period[7] ),
    .B1(\frequency_counter_0.update_period[6] ),
    .B2(_0133_),
    .X(_0145_));
 sky130_fd_sc_hd__inv_2 _0701_ (.A(\frequency_counter_0.clk_counter[4] ),
    .Y(_0146_));
 sky130_fd_sc_hd__o22a_1 _0702_ (.A1(_0134_),
    .A2(\frequency_counter_0.update_period[5] ),
    .B1(\frequency_counter_0.update_period[4] ),
    .B2(_0146_),
    .X(_0147_));
 sky130_fd_sc_hd__inv_2 _0703_ (.A(\frequency_counter_0.update_period[4] ),
    .Y(_0148_));
 sky130_fd_sc_hd__inv_2 _0704_ (.A(\frequency_counter_0.update_period[3] ),
    .Y(_0149_));
 sky130_fd_sc_hd__or2b_1 _0705_ (.A(\frequency_counter_0.clk_counter[7] ),
    .B_N(\frequency_counter_0.update_period[7] ),
    .X(_0150_));
 sky130_fd_sc_hd__o221a_1 _0706_ (.A1(\frequency_counter_0.clk_counter[4] ),
    .A2(_0148_),
    .B1(_0149_),
    .B2(\frequency_counter_0.clk_counter[3] ),
    .C1(_0150_),
    .X(_0151_));
 sky130_fd_sc_hd__and3_1 _0707_ (.A(_0145_),
    .B(_0147_),
    .C(_0151_),
    .X(_0152_));
 sky130_fd_sc_hd__a22o_1 _0708_ (.A1(_0133_),
    .A2(\frequency_counter_0.update_period[6] ),
    .B1(\frequency_counter_0.update_period[5] ),
    .B2(_0134_),
    .X(_0153_));
 sky130_fd_sc_hd__o21ai_1 _0709_ (.A1(_0153_),
    .A2(_0147_),
    .B1(_0145_),
    .Y(_0154_));
 sky130_fd_sc_hd__a32o_1 _0710_ (.A1(_0135_),
    .A2(_0143_),
    .A3(_0152_),
    .B1(_0154_),
    .B2(_0150_),
    .X(_0155_));
 sky130_fd_sc_hd__inv_2 _0711_ (.A(\frequency_counter_0.update_period[8] ),
    .Y(_0156_));
 sky130_fd_sc_hd__nand2_1 _0712_ (.A(_0127_),
    .B(\frequency_counter_0.update_period[10] ),
    .Y(_0157_));
 sky130_fd_sc_hd__and3b_1 _0713_ (.A_N(_0129_),
    .B(_0130_),
    .C(_0157_),
    .X(_0158_));
 sky130_fd_sc_hd__inv_2 _0714_ (.A(\frequency_counter_0.clk_counter[9] ),
    .Y(_0159_));
 sky130_fd_sc_hd__inv_2 _0715_ (.A(\frequency_counter_0.clk_counter[8] ),
    .Y(_0160_));
 sky130_fd_sc_hd__o22a_1 _0716_ (.A1(_0159_),
    .A2(\frequency_counter_0.update_period[9] ),
    .B1(\frequency_counter_0.update_period[8] ),
    .B2(_0160_),
    .X(_0161_));
 sky130_fd_sc_hd__nand2_1 _0717_ (.A(_0159_),
    .B(\frequency_counter_0.update_period[9] ),
    .Y(_0162_));
 sky130_fd_sc_hd__o2111a_1 _0718_ (.A1(\frequency_counter_0.clk_counter[8] ),
    .A2(_0156_),
    .B1(_0158_),
    .C1(_0161_),
    .D1(_0162_),
    .X(_0163_));
 sky130_fd_sc_hd__and3b_1 _0719_ (.A_N(_0161_),
    .B(_0162_),
    .C(_0158_),
    .X(_0164_));
 sky130_fd_sc_hd__a21oi_1 _0720_ (.A1(_0155_),
    .A2(_0163_),
    .B1(_0164_),
    .Y(_0165_));
 sky130_fd_sc_hd__nand2_1 _0721_ (.A(_0132_),
    .B(_0165_),
    .Y(_0166_));
 sky130_fd_sc_hd__clkbuf_4 _0722_ (.A(_0166_),
    .X(_0167_));
 sky130_fd_sc_hd__buf_2 _0723_ (.A(\frequency_counter_0.edge_counter[1] ),
    .X(_0168_));
 sky130_fd_sc_hd__o21a_1 _0724_ (.A1(\frequency_counter_0.edge_counter[2] ),
    .A2(_0168_),
    .B1(\frequency_counter_0.edge_counter[3] ),
    .X(_0169_));
 sky130_fd_sc_hd__or3_1 _0725_ (.A(\frequency_counter_0.dbg_edge_count[1] ),
    .B(\frequency_counter_0.dbg_edge_count[0] ),
    .C(_0169_),
    .X(_0170_));
 sky130_fd_sc_hd__clkinv_2 _0726_ (.A(\frequency_counter_0.dbg_state[0] ),
    .Y(_0171_));
 sky130_fd_sc_hd__or2_1 _0727_ (.A(\frequency_counter_0.dbg_state[1] ),
    .B(_0171_),
    .X(_0172_));
 sky130_fd_sc_hd__buf_2 _0728_ (.A(_0172_),
    .X(_0173_));
 sky130_fd_sc_hd__or3_1 _0729_ (.A(\frequency_counter_0.dbg_edge_count[2] ),
    .B(_0170_),
    .C(_0173_),
    .X(_0174_));
 sky130_fd_sc_hd__and2b_1 _0730_ (.A_N(\frequency_counter_0.dbg_state[1] ),
    .B(_0174_),
    .X(_0175_));
 sky130_fd_sc_hd__nand2_1 _0731_ (.A(_0167_),
    .B(_0175_),
    .Y(_0176_));
 sky130_fd_sc_hd__nor2_1 _0732_ (.A(_0081_),
    .B(_0176_),
    .Y(_0021_));
 sky130_fd_sc_hd__nor2_1 _0733_ (.A(_0081_),
    .B(_0174_),
    .Y(_0022_));
 sky130_fd_sc_hd__o211a_1 _0734_ (.A1(\frequency_counter_0.seven_segment0.load ),
    .A2(_0171_),
    .B1(_0083_),
    .C1(_0131_),
    .X(_0023_));
 sky130_fd_sc_hd__and2_1 _0735_ (.A(\frequency_counter_0.dbg_state[1] ),
    .B(_0171_),
    .X(_0177_));
 sky130_fd_sc_hd__clkbuf_2 _0736_ (.A(_0177_),
    .X(_0178_));
 sky130_fd_sc_hd__nand2_1 _0737_ (.A(\frequency_counter_0.edge_counter[0] ),
    .B(_0178_),
    .Y(_0179_));
 sky130_fd_sc_hd__a21bo_1 _0738_ (.A1(_0171_),
    .A2(_0167_),
    .B1_N(\frequency_counter_0.seven_segment0.unit_count[0] ),
    .X(_0180_));
 sky130_fd_sc_hd__a21oi_1 _0739_ (.A1(_0179_),
    .A2(_0180_),
    .B1(_0101_),
    .Y(_0024_));
 sky130_fd_sc_hd__nand2_1 _0740_ (.A(_0168_),
    .B(_0178_),
    .Y(_0181_));
 sky130_fd_sc_hd__a21bo_1 _0741_ (.A1(_0171_),
    .A2(_0167_),
    .B1_N(\frequency_counter_0.seven_segment0.unit_count[1] ),
    .X(_0182_));
 sky130_fd_sc_hd__a21oi_1 _0742_ (.A1(_0181_),
    .A2(_0182_),
    .B1(_0101_),
    .Y(_0025_));
 sky130_fd_sc_hd__nand2_1 _0743_ (.A(\frequency_counter_0.edge_counter[2] ),
    .B(_0178_),
    .Y(_0183_));
 sky130_fd_sc_hd__a21bo_1 _0744_ (.A1(_0171_),
    .A2(_0167_),
    .B1_N(\frequency_counter_0.seven_segment0.unit_count[2] ),
    .X(_0184_));
 sky130_fd_sc_hd__a21oi_1 _0745_ (.A1(_0183_),
    .A2(_0184_),
    .B1(_0101_),
    .Y(_0026_));
 sky130_fd_sc_hd__nand2_1 _0746_ (.A(\frequency_counter_0.edge_counter[3] ),
    .B(_0178_),
    .Y(_0185_));
 sky130_fd_sc_hd__a21bo_1 _0747_ (.A1(_0171_),
    .A2(_0167_),
    .B1_N(\frequency_counter_0.seven_segment0.unit_count[3] ),
    .X(_0186_));
 sky130_fd_sc_hd__a21oi_1 _0748_ (.A1(_0185_),
    .A2(_0186_),
    .B1(_0101_),
    .Y(_0027_));
 sky130_fd_sc_hd__inv_2 _0749_ (.A(\frequency_counter_0.seven_segment0.ten_count[0] ),
    .Y(_0187_));
 sky130_fd_sc_hd__a31o_1 _0750_ (.A1(\frequency_counter_0.dbg_state[0] ),
    .A2(_0167_),
    .A3(_0175_),
    .B1(\frequency_counter_0.seven_segment0.ten_count[0] ),
    .X(_0188_));
 sky130_fd_sc_hd__o211a_1 _0751_ (.A1(_0187_),
    .A2(_0176_),
    .B1(_0188_),
    .C1(_0083_),
    .X(_0028_));
 sky130_fd_sc_hd__a21oi_1 _0752_ (.A1(\frequency_counter_0.seven_segment0.ten_count[1] ),
    .A2(\frequency_counter_0.seven_segment0.ten_count[0] ),
    .B1(_0173_),
    .Y(_0189_));
 sky130_fd_sc_hd__a31o_1 _0753_ (.A1(\frequency_counter_0.seven_segment0.ten_count[0] ),
    .A2(_0167_),
    .A3(_0175_),
    .B1(\frequency_counter_0.seven_segment0.ten_count[1] ),
    .X(_0190_));
 sky130_fd_sc_hd__o211a_1 _0754_ (.A1(_0176_),
    .A2(_0189_),
    .B1(_0190_),
    .C1(_0083_),
    .X(_0029_));
 sky130_fd_sc_hd__and3_1 _0755_ (.A(\frequency_counter_0.seven_segment0.ten_count[2] ),
    .B(\frequency_counter_0.seven_segment0.ten_count[1] ),
    .C(\frequency_counter_0.seven_segment0.ten_count[0] ),
    .X(_0191_));
 sky130_fd_sc_hd__nor2_1 _0756_ (.A(_0173_),
    .B(_0191_),
    .Y(_0192_));
 sky130_fd_sc_hd__a41o_1 _0757_ (.A1(\frequency_counter_0.seven_segment0.ten_count[1] ),
    .A2(\frequency_counter_0.seven_segment0.ten_count[0] ),
    .A3(_0167_),
    .A4(_0175_),
    .B1(\frequency_counter_0.seven_segment0.ten_count[2] ),
    .X(_0193_));
 sky130_fd_sc_hd__o211a_1 _0758_ (.A1(_0176_),
    .A2(_0192_),
    .B1(_0193_),
    .C1(_0083_),
    .X(_0030_));
 sky130_fd_sc_hd__a41o_1 _0759_ (.A1(\frequency_counter_0.seven_segment0.ten_count[3] ),
    .A2(\frequency_counter_0.seven_segment0.ten_count[2] ),
    .A3(\frequency_counter_0.seven_segment0.ten_count[1] ),
    .A4(\frequency_counter_0.seven_segment0.ten_count[0] ),
    .B1(_0173_),
    .X(_0194_));
 sky130_fd_sc_hd__inv_2 _0760_ (.A(_0194_),
    .Y(_0195_));
 sky130_fd_sc_hd__a31o_1 _0761_ (.A1(_0167_),
    .A2(_0175_),
    .A3(_0191_),
    .B1(\frequency_counter_0.seven_segment0.ten_count[3] ),
    .X(_0196_));
 sky130_fd_sc_hd__o211a_1 _0762_ (.A1(_0176_),
    .A2(_0195_),
    .B1(_0196_),
    .C1(_0083_),
    .X(_0031_));
 sky130_fd_sc_hd__nor2_1 _0763_ (.A(\frequency_counter_0.dbg_state[1] ),
    .B(\frequency_counter_0.dbg_state[0] ),
    .Y(_0197_));
 sky130_fd_sc_hd__a21o_1 _0764_ (.A1(\frequency_counter_0.clk_counter[0] ),
    .A2(_0197_),
    .B1(_0080_),
    .X(_0198_));
 sky130_fd_sc_hd__a21oi_1 _0765_ (.A1(_0137_),
    .A2(_0167_),
    .B1(_0198_),
    .Y(_0032_));
 sky130_fd_sc_hd__clkbuf_4 _0766_ (.A(_0166_),
    .X(_0199_));
 sky130_fd_sc_hd__nor2_1 _0767_ (.A(\frequency_counter_0.clk_counter[1] ),
    .B(\frequency_counter_0.clk_counter[0] ),
    .Y(_0200_));
 sky130_fd_sc_hd__nor2_1 _0768_ (.A(_0136_),
    .B(_0137_),
    .Y(_0201_));
 sky130_fd_sc_hd__clkbuf_4 _0769_ (.A(_0197_),
    .X(_0202_));
 sky130_fd_sc_hd__o32a_1 _0770_ (.A1(_0199_),
    .A2(_0200_),
    .A3(_0201_),
    .B1(_0202_),
    .B2(_0136_),
    .X(_0203_));
 sky130_fd_sc_hd__nor2_1 _0771_ (.A(_0081_),
    .B(_0203_),
    .Y(_0033_));
 sky130_fd_sc_hd__nor2_1 _0772_ (.A(\frequency_counter_0.clk_counter[2] ),
    .B(_0201_),
    .Y(_0204_));
 sky130_fd_sc_hd__and3_1 _0773_ (.A(\frequency_counter_0.clk_counter[2] ),
    .B(\frequency_counter_0.clk_counter[1] ),
    .C(\frequency_counter_0.clk_counter[0] ),
    .X(_0205_));
 sky130_fd_sc_hd__o32a_1 _0774_ (.A1(_0199_),
    .A2(_0204_),
    .A3(_0205_),
    .B1(_0202_),
    .B2(_0139_),
    .X(_0206_));
 sky130_fd_sc_hd__nor2_1 _0775_ (.A(_0081_),
    .B(_0206_),
    .Y(_0034_));
 sky130_fd_sc_hd__nor2_1 _0776_ (.A(\frequency_counter_0.clk_counter[3] ),
    .B(_0205_),
    .Y(_0207_));
 sky130_fd_sc_hd__and2_1 _0777_ (.A(\frequency_counter_0.clk_counter[3] ),
    .B(_0205_),
    .X(_0208_));
 sky130_fd_sc_hd__o32a_1 _0778_ (.A1(_0199_),
    .A2(_0207_),
    .A3(_0208_),
    .B1(_0202_),
    .B2(_0141_),
    .X(_0209_));
 sky130_fd_sc_hd__nor2_1 _0779_ (.A(_0081_),
    .B(_0209_),
    .Y(_0035_));
 sky130_fd_sc_hd__nor2_1 _0780_ (.A(\frequency_counter_0.clk_counter[4] ),
    .B(_0208_),
    .Y(_0210_));
 sky130_fd_sc_hd__and3_1 _0781_ (.A(\frequency_counter_0.clk_counter[4] ),
    .B(\frequency_counter_0.clk_counter[3] ),
    .C(_0205_),
    .X(_0211_));
 sky130_fd_sc_hd__o32a_1 _0782_ (.A1(_0199_),
    .A2(_0210_),
    .A3(_0211_),
    .B1(_0202_),
    .B2(_0146_),
    .X(_0212_));
 sky130_fd_sc_hd__nor2_1 _0783_ (.A(_0081_),
    .B(_0212_),
    .Y(_0036_));
 sky130_fd_sc_hd__a21oi_1 _0784_ (.A1(\frequency_counter_0.clk_counter[4] ),
    .A2(_0208_),
    .B1(\frequency_counter_0.clk_counter[5] ),
    .Y(_0213_));
 sky130_fd_sc_hd__and3_1 _0785_ (.A(\frequency_counter_0.clk_counter[5] ),
    .B(\frequency_counter_0.clk_counter[4] ),
    .C(_0208_),
    .X(_0214_));
 sky130_fd_sc_hd__o32a_1 _0786_ (.A1(_0199_),
    .A2(_0213_),
    .A3(_0214_),
    .B1(_0202_),
    .B2(_0134_),
    .X(_0215_));
 sky130_fd_sc_hd__nor2_1 _0787_ (.A(_0081_),
    .B(_0215_),
    .Y(_0037_));
 sky130_fd_sc_hd__nor2_1 _0788_ (.A(\frequency_counter_0.clk_counter[6] ),
    .B(_0214_),
    .Y(_0216_));
 sky130_fd_sc_hd__and2_1 _0789_ (.A(\frequency_counter_0.clk_counter[6] ),
    .B(_0214_),
    .X(_0217_));
 sky130_fd_sc_hd__o32a_1 _0790_ (.A1(_0199_),
    .A2(_0216_),
    .A3(_0217_),
    .B1(_0202_),
    .B2(_0133_),
    .X(_0218_));
 sky130_fd_sc_hd__nor2_1 _0791_ (.A(_0081_),
    .B(_0218_),
    .Y(_0038_));
 sky130_fd_sc_hd__nor2_1 _0792_ (.A(\frequency_counter_0.clk_counter[7] ),
    .B(_0217_),
    .Y(_0219_));
 sky130_fd_sc_hd__and3_1 _0793_ (.A(\frequency_counter_0.clk_counter[7] ),
    .B(\frequency_counter_0.clk_counter[6] ),
    .C(_0214_),
    .X(_0220_));
 sky130_fd_sc_hd__o32a_1 _0794_ (.A1(_0199_),
    .A2(_0219_),
    .A3(_0220_),
    .B1(_0202_),
    .B2(_0144_),
    .X(_0221_));
 sky130_fd_sc_hd__nor2_1 _0795_ (.A(_0081_),
    .B(_0221_),
    .Y(_0039_));
 sky130_fd_sc_hd__nor2_1 _0796_ (.A(\frequency_counter_0.clk_counter[8] ),
    .B(_0220_),
    .Y(_0222_));
 sky130_fd_sc_hd__and2_1 _0797_ (.A(\frequency_counter_0.clk_counter[8] ),
    .B(_0220_),
    .X(_0223_));
 sky130_fd_sc_hd__o32a_1 _0798_ (.A1(_0199_),
    .A2(_0222_),
    .A3(_0223_),
    .B1(_0202_),
    .B2(_0160_),
    .X(_0224_));
 sky130_fd_sc_hd__nor2_1 _0799_ (.A(_0101_),
    .B(_0224_),
    .Y(_0040_));
 sky130_fd_sc_hd__nor2_1 _0800_ (.A(\frequency_counter_0.clk_counter[9] ),
    .B(_0223_),
    .Y(_0225_));
 sky130_fd_sc_hd__and3_1 _0801_ (.A(\frequency_counter_0.clk_counter[9] ),
    .B(\frequency_counter_0.clk_counter[8] ),
    .C(_0220_),
    .X(_0226_));
 sky130_fd_sc_hd__o32a_1 _0802_ (.A1(_0199_),
    .A2(_0225_),
    .A3(_0226_),
    .B1(_0202_),
    .B2(_0159_),
    .X(_0227_));
 sky130_fd_sc_hd__nor2_1 _0803_ (.A(_0101_),
    .B(_0227_),
    .Y(_0041_));
 sky130_fd_sc_hd__and2_1 _0804_ (.A(\frequency_counter_0.clk_counter[10] ),
    .B(_0226_),
    .X(_0228_));
 sky130_fd_sc_hd__nor2_1 _0805_ (.A(\frequency_counter_0.clk_counter[10] ),
    .B(_0226_),
    .Y(_0229_));
 sky130_fd_sc_hd__o32a_1 _0806_ (.A1(_0199_),
    .A2(_0228_),
    .A3(_0229_),
    .B1(_0202_),
    .B2(_0127_),
    .X(_0230_));
 sky130_fd_sc_hd__nor2_1 _0807_ (.A(_0101_),
    .B(_0230_),
    .Y(_0042_));
 sky130_fd_sc_hd__o211ai_1 _0808_ (.A1(_0166_),
    .A2(_0228_),
    .B1(\frequency_counter_0.clk_counter[11] ),
    .C1(_0197_),
    .Y(_0231_));
 sky130_fd_sc_hd__a31o_1 _0809_ (.A1(_0132_),
    .A2(_0165_),
    .A3(_0228_),
    .B1(\frequency_counter_0.clk_counter[11] ),
    .X(_0232_));
 sky130_fd_sc_hd__and3_1 _0810_ (.A(_0082_),
    .B(_0231_),
    .C(_0232_),
    .X(_0233_));
 sky130_fd_sc_hd__clkbuf_1 _0811_ (.A(_0233_),
    .X(_0043_));
 sky130_fd_sc_hd__nor2_1 _0812_ (.A(\frequency_counter_0.dbg_state[1] ),
    .B(_0171_),
    .Y(_0234_));
 sky130_fd_sc_hd__or2_1 _0813_ (.A(_0234_),
    .B(_0178_),
    .X(_0235_));
 sky130_fd_sc_hd__clkbuf_2 _0814_ (.A(_0235_),
    .X(_0236_));
 sky130_fd_sc_hd__clkinv_2 _0815_ (.A(\frequency_counter_0.edge_detect0.q2 ),
    .Y(_0237_));
 sky130_fd_sc_hd__and3_1 _0816_ (.A(_0171_),
    .B(\frequency_counter_0.edge_detect0.q1 ),
    .C(_0237_),
    .X(_0238_));
 sky130_fd_sc_hd__or2_1 _0817_ (.A(_0236_),
    .B(_0238_),
    .X(_0239_));
 sky130_fd_sc_hd__and2_1 _0818_ (.A(_0174_),
    .B(_0239_),
    .X(_0240_));
 sky130_fd_sc_hd__buf_2 _0819_ (.A(_0240_),
    .X(_0241_));
 sky130_fd_sc_hd__xnor2_1 _0820_ (.A(\frequency_counter_0.edge_counter[0] ),
    .B(_0168_),
    .Y(_0242_));
 sky130_fd_sc_hd__o221ai_1 _0821_ (.A1(_0168_),
    .A2(_0173_),
    .B1(_0236_),
    .B2(_0242_),
    .C1(_0241_),
    .Y(_0243_));
 sky130_fd_sc_hd__o211a_1 _0822_ (.A1(_0168_),
    .A2(_0241_),
    .B1(_0243_),
    .C1(_0083_),
    .X(_0044_));
 sky130_fd_sc_hd__a21oi_1 _0823_ (.A1(\frequency_counter_0.edge_counter[0] ),
    .A2(_0168_),
    .B1(\frequency_counter_0.edge_counter[2] ),
    .Y(_0244_));
 sky130_fd_sc_hd__and3_1 _0824_ (.A(\frequency_counter_0.edge_counter[0] ),
    .B(\frequency_counter_0.edge_counter[2] ),
    .C(_0168_),
    .X(_0245_));
 sky130_fd_sc_hd__xor2_1 _0825_ (.A(\frequency_counter_0.edge_counter[2] ),
    .B(_0168_),
    .X(_0246_));
 sky130_fd_sc_hd__o32a_1 _0826_ (.A1(_0236_),
    .A2(_0244_),
    .A3(_0245_),
    .B1(_0246_),
    .B2(_0173_),
    .X(_0247_));
 sky130_fd_sc_hd__nand2_1 _0827_ (.A(_0241_),
    .B(_0247_),
    .Y(_0248_));
 sky130_fd_sc_hd__o211a_1 _0828_ (.A1(\frequency_counter_0.edge_counter[2] ),
    .A2(_0241_),
    .B1(_0248_),
    .C1(_0083_),
    .X(_0045_));
 sky130_fd_sc_hd__nor2_1 _0829_ (.A(_0169_),
    .B(_0173_),
    .Y(_0249_));
 sky130_fd_sc_hd__o31a_1 _0830_ (.A1(\frequency_counter_0.edge_counter[3] ),
    .A2(\frequency_counter_0.edge_counter[2] ),
    .A3(_0168_),
    .B1(_0249_),
    .X(_0250_));
 sky130_fd_sc_hd__and2_1 _0831_ (.A(\frequency_counter_0.edge_counter[3] ),
    .B(_0245_),
    .X(_0251_));
 sky130_fd_sc_hd__nor2_1 _0832_ (.A(_0236_),
    .B(_0251_),
    .Y(_0252_));
 sky130_fd_sc_hd__o21ai_1 _0833_ (.A1(\frequency_counter_0.edge_counter[3] ),
    .A2(_0245_),
    .B1(_0252_),
    .Y(_0253_));
 sky130_fd_sc_hd__nand2_1 _0834_ (.A(_0241_),
    .B(_0253_),
    .Y(_0254_));
 sky130_fd_sc_hd__o221a_1 _0835_ (.A1(\frequency_counter_0.edge_counter[3] ),
    .A2(_0241_),
    .B1(_0250_),
    .B2(_0254_),
    .C1(_0083_),
    .X(_0046_));
 sky130_fd_sc_hd__and2b_1 _0836_ (.A_N(_0236_),
    .B(_0251_),
    .X(_0255_));
 sky130_fd_sc_hd__o21a_1 _0837_ (.A1(_0249_),
    .A2(_0255_),
    .B1(_0241_),
    .X(_0256_));
 sky130_fd_sc_hd__a21bo_1 _0838_ (.A1(_0169_),
    .A2(_0234_),
    .B1_N(\frequency_counter_0.dbg_edge_count[0] ),
    .X(_0257_));
 sky130_fd_sc_hd__or3b_1 _0839_ (.A(_0252_),
    .B(_0257_),
    .C_N(_0240_),
    .X(_0258_));
 sky130_fd_sc_hd__o211a_1 _0840_ (.A1(\frequency_counter_0.dbg_edge_count[0] ),
    .A2(_0256_),
    .B1(_0258_),
    .C1(_0083_),
    .X(_0047_));
 sky130_fd_sc_hd__a21oi_1 _0841_ (.A1(\frequency_counter_0.dbg_edge_count[0] ),
    .A2(_0251_),
    .B1(\frequency_counter_0.dbg_edge_count[1] ),
    .Y(_0259_));
 sky130_fd_sc_hd__and3_1 _0842_ (.A(\frequency_counter_0.dbg_edge_count[1] ),
    .B(\frequency_counter_0.dbg_edge_count[0] ),
    .C(_0251_),
    .X(_0260_));
 sky130_fd_sc_hd__or3_1 _0843_ (.A(_0236_),
    .B(_0259_),
    .C(_0260_),
    .X(_0261_));
 sky130_fd_sc_hd__o21ai_1 _0844_ (.A1(\frequency_counter_0.dbg_edge_count[0] ),
    .A2(_0169_),
    .B1(\frequency_counter_0.dbg_edge_count[1] ),
    .Y(_0262_));
 sky130_fd_sc_hd__a21o_1 _0845_ (.A1(_0170_),
    .A2(_0262_),
    .B1(_0173_),
    .X(_0263_));
 sky130_fd_sc_hd__a31o_1 _0846_ (.A1(_0241_),
    .A2(_0261_),
    .A3(_0263_),
    .B1(_0080_),
    .X(_0264_));
 sky130_fd_sc_hd__o21ba_1 _0847_ (.A1(\frequency_counter_0.dbg_edge_count[1] ),
    .A2(_0241_),
    .B1_N(_0264_),
    .X(_0048_));
 sky130_fd_sc_hd__a2bb2o_1 _0848_ (.A1_N(_0236_),
    .A2_N(_0260_),
    .B1(_0170_),
    .B2(_0234_),
    .X(_0265_));
 sky130_fd_sc_hd__nor2_1 _0849_ (.A(\frequency_counter_0.dbg_edge_count[2] ),
    .B(_0236_),
    .Y(_0266_));
 sky130_fd_sc_hd__a22o_1 _0850_ (.A1(\frequency_counter_0.dbg_edge_count[2] ),
    .A2(_0265_),
    .B1(_0266_),
    .B2(_0260_),
    .X(_0267_));
 sky130_fd_sc_hd__clkinv_2 _0851_ (.A(\frequency_counter_0.dbg_edge_count[2] ),
    .Y(_0268_));
 sky130_fd_sc_hd__o2bb2a_1 _0852_ (.A1_N(_0241_),
    .A2_N(_0267_),
    .B1(_0268_),
    .B2(_0239_),
    .X(_0269_));
 sky130_fd_sc_hd__nor2_1 _0853_ (.A(_0101_),
    .B(_0269_),
    .Y(_0049_));
 sky130_fd_sc_hd__a211o_1 _0854_ (.A1(\frequency_counter_0.edge_counter[0] ),
    .A2(_0238_),
    .B1(_0178_),
    .C1(_0080_),
    .X(_0270_));
 sky130_fd_sc_hd__o21ba_1 _0855_ (.A1(\frequency_counter_0.edge_counter[0] ),
    .A2(_0238_),
    .B1_N(_0270_),
    .X(_0050_));
 sky130_fd_sc_hd__dfxtp_2 _0856_ (.CLK(clknet_2_3__leaf_wb_clk_i),
    .D(_0000_),
    .Q(\frequency_counter_0.digit ));
 sky130_fd_sc_hd__dfxtp_1 _0857_ (.CLK(clknet_2_1__leaf_wb_clk_i),
    .D(_0001_),
    .Q(\frequency_counter_0.seven_segment0.ten_count_reg[0] ));
 sky130_fd_sc_hd__dfxtp_1 _0858_ (.CLK(clknet_2_0__leaf_wb_clk_i),
    .D(_0002_),
    .Q(\frequency_counter_0.seven_segment0.ten_count_reg[1] ));
 sky130_fd_sc_hd__dfxtp_1 _0859_ (.CLK(clknet_2_0__leaf_wb_clk_i),
    .D(_0003_),
    .Q(\frequency_counter_0.seven_segment0.ten_count_reg[2] ));
 sky130_fd_sc_hd__dfxtp_1 _0860_ (.CLK(clknet_2_0__leaf_wb_clk_i),
    .D(_0004_),
    .Q(\frequency_counter_0.seven_segment0.ten_count_reg[3] ));
 sky130_fd_sc_hd__dfxtp_1 _0861_ (.CLK(clknet_2_0__leaf_wb_clk_i),
    .D(_0005_),
    .Q(\frequency_counter_0.seven_segment0.unit_count_reg[0] ));
 sky130_fd_sc_hd__dfxtp_1 _0862_ (.CLK(clknet_2_0__leaf_wb_clk_i),
    .D(_0006_),
    .Q(\frequency_counter_0.seven_segment0.unit_count_reg[1] ));
 sky130_fd_sc_hd__dfxtp_1 _0863_ (.CLK(clknet_2_0__leaf_wb_clk_i),
    .D(_0007_),
    .Q(\frequency_counter_0.seven_segment0.unit_count_reg[2] ));
 sky130_fd_sc_hd__dfxtp_1 _0864_ (.CLK(clknet_2_2__leaf_wb_clk_i),
    .D(_0008_),
    .Q(\frequency_counter_0.seven_segment0.unit_count_reg[3] ));
 sky130_fd_sc_hd__dfxtp_1 _0865_ (.CLK(clknet_2_3__leaf_wb_clk_i),
    .D(net2),
    .Q(\frequency_counter_0.edge_detect0.q0 ));
 sky130_fd_sc_hd__dfxtp_1 _0866_ (.CLK(clknet_2_3__leaf_wb_clk_i),
    .D(net108),
    .Q(\frequency_counter_0.edge_detect0.q1 ));
 sky130_fd_sc_hd__dfxtp_1 _0867_ (.CLK(clknet_2_3__leaf_wb_clk_i),
    .D(net109),
    .Q(\frequency_counter_0.edge_detect0.q2 ));
 sky130_fd_sc_hd__dfxtp_1 _0868_ (.CLK(clknet_2_2__leaf_wb_clk_i),
    .D(_0009_),
    .Q(\frequency_counter_0.update_period[0] ));
 sky130_fd_sc_hd__dfxtp_1 _0869_ (.CLK(clknet_2_2__leaf_wb_clk_i),
    .D(_0010_),
    .Q(\frequency_counter_0.update_period[1] ));
 sky130_fd_sc_hd__dfxtp_1 _0870_ (.CLK(clknet_2_3__leaf_wb_clk_i),
    .D(_0011_),
    .Q(\frequency_counter_0.update_period[2] ));
 sky130_fd_sc_hd__dfxtp_1 _0871_ (.CLK(clknet_2_3__leaf_wb_clk_i),
    .D(_0012_),
    .Q(\frequency_counter_0.update_period[3] ));
 sky130_fd_sc_hd__dfxtp_1 _0872_ (.CLK(clknet_2_2__leaf_wb_clk_i),
    .D(_0013_),
    .Q(\frequency_counter_0.update_period[4] ));
 sky130_fd_sc_hd__dfxtp_1 _0873_ (.CLK(clknet_2_0__leaf_wb_clk_i),
    .D(_0014_),
    .Q(\frequency_counter_0.update_period[5] ));
 sky130_fd_sc_hd__dfxtp_1 _0874_ (.CLK(clknet_2_2__leaf_wb_clk_i),
    .D(_0015_),
    .Q(\frequency_counter_0.update_period[6] ));
 sky130_fd_sc_hd__dfxtp_1 _0875_ (.CLK(clknet_2_2__leaf_wb_clk_i),
    .D(_0016_),
    .Q(\frequency_counter_0.update_period[7] ));
 sky130_fd_sc_hd__dfxtp_1 _0876_ (.CLK(clknet_2_0__leaf_wb_clk_i),
    .D(_0017_),
    .Q(\frequency_counter_0.update_period[8] ));
 sky130_fd_sc_hd__dfxtp_1 _0877_ (.CLK(clknet_2_1__leaf_wb_clk_i),
    .D(_0018_),
    .Q(\frequency_counter_0.update_period[9] ));
 sky130_fd_sc_hd__dfxtp_1 _0878_ (.CLK(clknet_2_0__leaf_wb_clk_i),
    .D(_0019_),
    .Q(\frequency_counter_0.update_period[10] ));
 sky130_fd_sc_hd__dfxtp_1 _0879_ (.CLK(clknet_2_1__leaf_wb_clk_i),
    .D(_0020_),
    .Q(\frequency_counter_0.update_period[11] ));
 sky130_fd_sc_hd__dfxtp_2 _0880_ (.CLK(clknet_2_1__leaf_wb_clk_i),
    .D(_0021_),
    .Q(\frequency_counter_0.dbg_state[0] ));
 sky130_fd_sc_hd__dfxtp_2 _0881_ (.CLK(clknet_2_3__leaf_wb_clk_i),
    .D(_0022_),
    .Q(\frequency_counter_0.dbg_state[1] ));
 sky130_fd_sc_hd__dfxtp_2 _0882_ (.CLK(clknet_2_1__leaf_wb_clk_i),
    .D(_0023_),
    .Q(\frequency_counter_0.seven_segment0.load ));
 sky130_fd_sc_hd__dfxtp_1 _0883_ (.CLK(clknet_2_3__leaf_wb_clk_i),
    .D(_0024_),
    .Q(\frequency_counter_0.seven_segment0.unit_count[0] ));
 sky130_fd_sc_hd__dfxtp_1 _0884_ (.CLK(clknet_2_2__leaf_wb_clk_i),
    .D(_0025_),
    .Q(\frequency_counter_0.seven_segment0.unit_count[1] ));
 sky130_fd_sc_hd__dfxtp_1 _0885_ (.CLK(clknet_2_1__leaf_wb_clk_i),
    .D(_0026_),
    .Q(\frequency_counter_0.seven_segment0.unit_count[2] ));
 sky130_fd_sc_hd__dfxtp_1 _0886_ (.CLK(clknet_2_1__leaf_wb_clk_i),
    .D(_0027_),
    .Q(\frequency_counter_0.seven_segment0.unit_count[3] ));
 sky130_fd_sc_hd__dfxtp_2 _0887_ (.CLK(clknet_2_1__leaf_wb_clk_i),
    .D(_0028_),
    .Q(\frequency_counter_0.seven_segment0.ten_count[0] ));
 sky130_fd_sc_hd__dfxtp_1 _0888_ (.CLK(clknet_2_1__leaf_wb_clk_i),
    .D(_0029_),
    .Q(\frequency_counter_0.seven_segment0.ten_count[1] ));
 sky130_fd_sc_hd__dfxtp_1 _0889_ (.CLK(clknet_2_1__leaf_wb_clk_i),
    .D(_0030_),
    .Q(\frequency_counter_0.seven_segment0.ten_count[2] ));
 sky130_fd_sc_hd__dfxtp_1 _0890_ (.CLK(clknet_2_0__leaf_wb_clk_i),
    .D(_0031_),
    .Q(\frequency_counter_0.seven_segment0.ten_count[3] ));
 sky130_fd_sc_hd__dfxtp_1 _0891_ (.CLK(clknet_2_2__leaf_wb_clk_i),
    .D(_0032_),
    .Q(\frequency_counter_0.clk_counter[0] ));
 sky130_fd_sc_hd__dfxtp_1 _0892_ (.CLK(clknet_2_2__leaf_wb_clk_i),
    .D(_0033_),
    .Q(\frequency_counter_0.clk_counter[1] ));
 sky130_fd_sc_hd__dfxtp_1 _0893_ (.CLK(clknet_2_3__leaf_wb_clk_i),
    .D(_0034_),
    .Q(\frequency_counter_0.clk_counter[2] ));
 sky130_fd_sc_hd__dfxtp_1 _0894_ (.CLK(clknet_2_2__leaf_wb_clk_i),
    .D(_0035_),
    .Q(\frequency_counter_0.clk_counter[3] ));
 sky130_fd_sc_hd__dfxtp_1 _0895_ (.CLK(clknet_2_2__leaf_wb_clk_i),
    .D(_0036_),
    .Q(\frequency_counter_0.clk_counter[4] ));
 sky130_fd_sc_hd__dfxtp_1 _0896_ (.CLK(clknet_2_2__leaf_wb_clk_i),
    .D(_0037_),
    .Q(\frequency_counter_0.clk_counter[5] ));
 sky130_fd_sc_hd__dfxtp_1 _0897_ (.CLK(clknet_2_2__leaf_wb_clk_i),
    .D(_0038_),
    .Q(\frequency_counter_0.clk_counter[6] ));
 sky130_fd_sc_hd__dfxtp_1 _0898_ (.CLK(clknet_2_2__leaf_wb_clk_i),
    .D(_0039_),
    .Q(\frequency_counter_0.clk_counter[7] ));
 sky130_fd_sc_hd__dfxtp_1 _0899_ (.CLK(clknet_2_0__leaf_wb_clk_i),
    .D(_0040_),
    .Q(\frequency_counter_0.clk_counter[8] ));
 sky130_fd_sc_hd__dfxtp_2 _0900_ (.CLK(clknet_2_2__leaf_wb_clk_i),
    .D(_0041_),
    .Q(\frequency_counter_0.clk_counter[9] ));
 sky130_fd_sc_hd__dfxtp_1 _0901_ (.CLK(clknet_2_2__leaf_wb_clk_i),
    .D(_0042_),
    .Q(\frequency_counter_0.clk_counter[10] ));
 sky130_fd_sc_hd__dfxtp_1 _0902_ (.CLK(clknet_2_0__leaf_wb_clk_i),
    .D(_0043_),
    .Q(\frequency_counter_0.clk_counter[11] ));
 sky130_fd_sc_hd__dfxtp_1 _0903_ (.CLK(clknet_2_1__leaf_wb_clk_i),
    .D(_0044_),
    .Q(\frequency_counter_0.edge_counter[1] ));
 sky130_fd_sc_hd__dfxtp_2 _0904_ (.CLK(clknet_2_1__leaf_wb_clk_i),
    .D(_0045_),
    .Q(\frequency_counter_0.edge_counter[2] ));
 sky130_fd_sc_hd__dfxtp_1 _0905_ (.CLK(clknet_2_3__leaf_wb_clk_i),
    .D(_0046_),
    .Q(\frequency_counter_0.edge_counter[3] ));
 sky130_fd_sc_hd__dfxtp_1 _0906_ (.CLK(clknet_2_3__leaf_wb_clk_i),
    .D(_0047_),
    .Q(\frequency_counter_0.dbg_edge_count[0] ));
 sky130_fd_sc_hd__dfxtp_2 _0907_ (.CLK(clknet_2_1__leaf_wb_clk_i),
    .D(_0048_),
    .Q(\frequency_counter_0.dbg_edge_count[1] ));
 sky130_fd_sc_hd__dfxtp_1 _0908_ (.CLK(clknet_2_3__leaf_wb_clk_i),
    .D(_0049_),
    .Q(\frequency_counter_0.dbg_edge_count[2] ));
 sky130_fd_sc_hd__dfxtp_1 _0909_ (.CLK(clknet_2_3__leaf_wb_clk_i),
    .D(_0050_),
    .Q(\frequency_counter_0.edge_counter[0] ));
 sky130_fd_sc_hd__conb_1 _1002__18 (.LO(net18));
 sky130_fd_sc_hd__conb_1 _1003__19 (.LO(net19));
 sky130_fd_sc_hd__conb_1 _1004__20 (.LO(net20));
 sky130_fd_sc_hd__conb_1 _1005__21 (.LO(net21));
 sky130_fd_sc_hd__conb_1 _1006__22 (.LO(net22));
 sky130_fd_sc_hd__conb_1 _1007__23 (.LO(net23));
 sky130_fd_sc_hd__conb_1 _1008__24 (.LO(net24));
 sky130_fd_sc_hd__conb_1 _1009__25 (.LO(net25));
 sky130_fd_sc_hd__conb_1 _1010__26 (.LO(net26));
 sky130_fd_sc_hd__conb_1 _1011__27 (.LO(net27));
 sky130_fd_sc_hd__conb_1 _1012__28 (.LO(net28));
 sky130_fd_sc_hd__conb_1 _1013__29 (.LO(net29));
 sky130_fd_sc_hd__conb_1 _1014__30 (.LO(net30));
 sky130_fd_sc_hd__conb_1 _1015__31 (.LO(net31));
 sky130_fd_sc_hd__conb_1 _1016__32 (.LO(net32));
 sky130_fd_sc_hd__conb_1 _1017__33 (.LO(net33));
 sky130_fd_sc_hd__conb_1 _1018__34 (.LO(net34));
 sky130_fd_sc_hd__conb_1 _1019__35 (.LO(net35));
 sky130_fd_sc_hd__conb_1 _1020__36 (.LO(net36));
 sky130_fd_sc_hd__conb_1 _1021__37 (.LO(net37));
 sky130_fd_sc_hd__conb_1 _1022__38 (.LO(net38));
 sky130_fd_sc_hd__conb_1 _1023__39 (.LO(net39));
 sky130_fd_sc_hd__conb_1 _1024__40 (.LO(net40));
 sky130_fd_sc_hd__conb_1 _1025__41 (.LO(net41));
 sky130_fd_sc_hd__conb_1 _1026__42 (.LO(net42));
 sky130_fd_sc_hd__conb_1 _1027__43 (.LO(net43));
 sky130_fd_sc_hd__conb_1 _1028__44 (.LO(net44));
 sky130_fd_sc_hd__conb_1 _1029__45 (.LO(net45));
 sky130_fd_sc_hd__conb_1 _1030__46 (.LO(net46));
 sky130_fd_sc_hd__conb_1 _1031__47 (.LO(net47));
 sky130_fd_sc_hd__conb_1 _1032__48 (.LO(net48));
 sky130_fd_sc_hd__conb_1 _1033__49 (.LO(net49));
 sky130_fd_sc_hd__conb_1 _1034__50 (.LO(net50));
 sky130_fd_sc_hd__conb_1 _1035__51 (.LO(net51));
 sky130_fd_sc_hd__conb_1 _1036__52 (.LO(net52));
 sky130_fd_sc_hd__conb_1 _1037__53 (.LO(net53));
 sky130_fd_sc_hd__conb_1 _1038__54 (.LO(net54));
 sky130_fd_sc_hd__conb_1 _1039__55 (.LO(net55));
 sky130_fd_sc_hd__conb_1 _1040__56 (.LO(net56));
 sky130_fd_sc_hd__conb_1 _1041__57 (.LO(net57));
 sky130_fd_sc_hd__conb_1 _1059__58 (.LO(net58));
 sky130_fd_sc_hd__conb_1 _1060__59 (.LO(net59));
 sky130_fd_sc_hd__conb_1 _1061__60 (.LO(net60));
 sky130_fd_sc_hd__conb_1 _1062__61 (.LO(net61));
 sky130_fd_sc_hd__conb_1 _1063__62 (.LO(net62));
 sky130_fd_sc_hd__conb_1 _1064__63 (.LO(net63));
 sky130_fd_sc_hd__conb_1 _1065__64 (.LO(net64));
 sky130_fd_sc_hd__conb_1 _1066__65 (.LO(net65));
 sky130_fd_sc_hd__conb_1 _1067__66 (.LO(net66));
 sky130_fd_sc_hd__conb_1 _1068__67 (.LO(net67));
 sky130_fd_sc_hd__conb_1 _1069__68 (.LO(net68));
 sky130_fd_sc_hd__conb_1 _1070__69 (.LO(net69));
 sky130_fd_sc_hd__conb_1 _1071__70 (.LO(net70));
 sky130_fd_sc_hd__conb_1 _1072__71 (.LO(net71));
 sky130_fd_sc_hd__conb_1 _1073__72 (.LO(net72));
 sky130_fd_sc_hd__conb_1 _1074__73 (.LO(net73));
 sky130_fd_sc_hd__conb_1 _1075__74 (.LO(net74));
 sky130_fd_sc_hd__conb_1 _1076__75 (.LO(net75));
 sky130_fd_sc_hd__conb_1 _1077__76 (.LO(net76));
 sky130_fd_sc_hd__conb_1 _1078__77 (.LO(net77));
 sky130_fd_sc_hd__conb_1 _1079__78 (.LO(net78));
 sky130_fd_sc_hd__conb_1 _1080__79 (.LO(net79));
 sky130_fd_sc_hd__conb_1 _1081__80 (.LO(net80));
 sky130_fd_sc_hd__conb_1 _1082__81 (.LO(net81));
 sky130_fd_sc_hd__conb_1 _1083__82 (.LO(net82));
 sky130_fd_sc_hd__conb_1 _1084__83 (.LO(net83));
 sky130_fd_sc_hd__conb_1 _1085__84 (.LO(net84));
 sky130_fd_sc_hd__conb_1 _1086__85 (.LO(net85));
 sky130_fd_sc_hd__conb_1 _1087__86 (.LO(net86));
 sky130_fd_sc_hd__conb_1 _1088__87 (.LO(net87));
 sky130_fd_sc_hd__conb_1 _1089__88 (.LO(net88));
 sky130_fd_sc_hd__conb_1 _1090__89 (.LO(net89));
 sky130_fd_sc_hd__conb_1 _1091__90 (.LO(net90));
 sky130_fd_sc_hd__conb_1 _1092__91 (.LO(net91));
 sky130_fd_sc_hd__conb_1 _1093__92 (.LO(net92));
 sky130_fd_sc_hd__conb_1 _1094__93 (.LO(net93));
 sky130_fd_sc_hd__conb_1 _1095__94 (.LO(net94));
 sky130_fd_sc_hd__conb_1 _1096__95 (.LO(net95));
 sky130_fd_sc_hd__conb_1 _1097__96 (.LO(net96));
 sky130_fd_sc_hd__conb_1 _1098__97 (.LO(net97));
 sky130_fd_sc_hd__conb_1 _1099__98 (.LO(net98));
 sky130_fd_sc_hd__conb_1 _1100__99 (.LO(net99));
 sky130_fd_sc_hd__conb_1 _1101__100 (.LO(net100));
 sky130_fd_sc_hd__conb_1 _1102__101 (.LO(net101));
 sky130_fd_sc_hd__conb_1 _1103__102 (.LO(net102));
 sky130_fd_sc_hd__conb_1 _1104__103 (.LO(net103));
 sky130_fd_sc_hd__conb_1 _1105__104 (.LO(net104));
 sky130_fd_sc_hd__conb_1 _1106__105 (.LO(net105));
 sky130_fd_sc_hd__conb_1 _1107__106 (.LO(net106));
 sky130_fd_sc_hd__conb_1 _1108__107 (.LO(net107));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_wb_clk_i (.A(wb_clk_i),
    .X(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__ebufn_8 _1001_ (.A(net17),
    .TE_B(_0271_),
    .Z(la1_data_out[0]));
 sky130_fd_sc_hd__ebufn_8 _1002_ (.A(net18),
    .TE_B(_0272_),
    .Z(la1_data_out[1]));
 sky130_fd_sc_hd__ebufn_8 _1003_ (.A(net19),
    .TE_B(_0273_),
    .Z(la1_data_out[2]));
 sky130_fd_sc_hd__ebufn_8 _1004_ (.A(net20),
    .TE_B(_0274_),
    .Z(la1_data_out[3]));
 sky130_fd_sc_hd__ebufn_8 _1005_ (.A(net21),
    .TE_B(_0275_),
    .Z(la1_data_out[4]));
 sky130_fd_sc_hd__ebufn_8 _1006_ (.A(net22),
    .TE_B(_0276_),
    .Z(la1_data_out[5]));
 sky130_fd_sc_hd__ebufn_8 _1007_ (.A(net23),
    .TE_B(_0277_),
    .Z(la1_data_out[6]));
 sky130_fd_sc_hd__ebufn_8 _1008_ (.A(net24),
    .TE_B(_0278_),
    .Z(la1_data_out[7]));
 sky130_fd_sc_hd__ebufn_8 _1009_ (.A(net25),
    .TE_B(_0279_),
    .Z(la1_data_out[8]));
 sky130_fd_sc_hd__ebufn_8 _1010_ (.A(net26),
    .TE_B(_0280_),
    .Z(la1_data_out[9]));
 sky130_fd_sc_hd__ebufn_8 _1011_ (.A(net27),
    .TE_B(_0281_),
    .Z(la1_data_out[10]));
 sky130_fd_sc_hd__ebufn_8 _1012_ (.A(net28),
    .TE_B(_0282_),
    .Z(la1_data_out[11]));
 sky130_fd_sc_hd__ebufn_8 _1013_ (.A(net29),
    .TE_B(_0283_),
    .Z(la1_data_out[12]));
 sky130_fd_sc_hd__ebufn_8 _1014_ (.A(net30),
    .TE_B(_0284_),
    .Z(la1_data_out[13]));
 sky130_fd_sc_hd__ebufn_8 _1015_ (.A(net31),
    .TE_B(_0285_),
    .Z(la1_data_out[14]));
 sky130_fd_sc_hd__ebufn_8 _1016_ (.A(net32),
    .TE_B(_0286_),
    .Z(la1_data_out[15]));
 sky130_fd_sc_hd__ebufn_8 _1017_ (.A(net33),
    .TE_B(_0287_),
    .Z(la1_data_out[16]));
 sky130_fd_sc_hd__ebufn_8 _1018_ (.A(net34),
    .TE_B(_0288_),
    .Z(la1_data_out[17]));
 sky130_fd_sc_hd__ebufn_8 _1019_ (.A(net35),
    .TE_B(_0289_),
    .Z(la1_data_out[18]));
 sky130_fd_sc_hd__ebufn_8 _1020_ (.A(net36),
    .TE_B(_0290_),
    .Z(la1_data_out[19]));
 sky130_fd_sc_hd__ebufn_8 _1021_ (.A(net37),
    .TE_B(_0291_),
    .Z(la1_data_out[20]));
 sky130_fd_sc_hd__ebufn_8 _1022_ (.A(net38),
    .TE_B(_0292_),
    .Z(la1_data_out[21]));
 sky130_fd_sc_hd__ebufn_8 _1023_ (.A(net39),
    .TE_B(_0293_),
    .Z(la1_data_out[22]));
 sky130_fd_sc_hd__ebufn_8 _1024_ (.A(net40),
    .TE_B(_0294_),
    .Z(la1_data_out[23]));
 sky130_fd_sc_hd__ebufn_8 _1025_ (.A(net41),
    .TE_B(_0295_),
    .Z(la1_data_out[24]));
 sky130_fd_sc_hd__ebufn_8 _1026_ (.A(net42),
    .TE_B(_0296_),
    .Z(la1_data_out[25]));
 sky130_fd_sc_hd__ebufn_8 _1027_ (.A(net43),
    .TE_B(_0297_),
    .Z(la1_data_out[26]));
 sky130_fd_sc_hd__ebufn_8 _1028_ (.A(net44),
    .TE_B(_0298_),
    .Z(la1_data_out[27]));
 sky130_fd_sc_hd__ebufn_8 _1029_ (.A(net45),
    .TE_B(_0299_),
    .Z(la1_data_out[28]));
 sky130_fd_sc_hd__ebufn_8 _1030_ (.A(net46),
    .TE_B(_0300_),
    .Z(la1_data_out[29]));
 sky130_fd_sc_hd__ebufn_8 _1031_ (.A(net47),
    .TE_B(_0301_),
    .Z(la1_data_out[30]));
 sky130_fd_sc_hd__ebufn_8 _1032_ (.A(net48),
    .TE_B(_0302_),
    .Z(la1_data_out[31]));
 sky130_fd_sc_hd__ebufn_8 _1033_ (.A(net49),
    .TE_B(_0303_),
    .Z(io_out[0]));
 sky130_fd_sc_hd__ebufn_8 _1034_ (.A(net50),
    .TE_B(_0304_),
    .Z(io_out[1]));
 sky130_fd_sc_hd__ebufn_8 _1035_ (.A(net51),
    .TE_B(_0305_),
    .Z(io_out[2]));
 sky130_fd_sc_hd__ebufn_8 _1036_ (.A(net52),
    .TE_B(_0306_),
    .Z(io_out[3]));
 sky130_fd_sc_hd__ebufn_8 _1037_ (.A(net53),
    .TE_B(_0307_),
    .Z(io_out[4]));
 sky130_fd_sc_hd__ebufn_8 _1038_ (.A(net54),
    .TE_B(_0308_),
    .Z(io_out[5]));
 sky130_fd_sc_hd__ebufn_8 _1039_ (.A(net55),
    .TE_B(_0309_),
    .Z(io_out[6]));
 sky130_fd_sc_hd__ebufn_8 _1040_ (.A(net56),
    .TE_B(_0310_),
    .Z(io_out[7]));
 sky130_fd_sc_hd__ebufn_8 _1041_ (.A(net57),
    .TE_B(_0311_),
    .Z(io_out[8]));
 sky130_fd_sc_hd__ebufn_8 _1042_ (.A(\frequency_counter_0.segments[0] ),
    .TE_B(_0312_),
    .Z(io_out[9]));
 sky130_fd_sc_hd__ebufn_8 _1043_ (.A(\frequency_counter_0.segments[1] ),
    .TE_B(_0313_),
    .Z(io_out[10]));
 sky130_fd_sc_hd__ebufn_8 _1044_ (.A(\frequency_counter_0.segments[2] ),
    .TE_B(_0314_),
    .Z(io_out[11]));
 sky130_fd_sc_hd__ebufn_8 _1045_ (.A(\frequency_counter_0.segments[3] ),
    .TE_B(_0315_),
    .Z(io_out[12]));
 sky130_fd_sc_hd__ebufn_8 _1046_ (.A(\frequency_counter_0.segments[4] ),
    .TE_B(_0316_),
    .Z(io_out[13]));
 sky130_fd_sc_hd__ebufn_8 _1047_ (.A(\frequency_counter_0.segments[5] ),
    .TE_B(_0317_),
    .Z(io_out[14]));
 sky130_fd_sc_hd__ebufn_8 _1048_ (.A(\frequency_counter_0.segments[6] ),
    .TE_B(_0318_),
    .Z(io_out[15]));
 sky130_fd_sc_hd__ebufn_8 _1049_ (.A(\frequency_counter_0.digit ),
    .TE_B(_0319_),
    .Z(io_out[16]));
 sky130_fd_sc_hd__ebufn_8 _1050_ (.A(net1),
    .TE_B(_0320_),
    .Z(io_out[17]));
 sky130_fd_sc_hd__ebufn_8 _1051_ (.A(\frequency_counter_0.dbg_state[0] ),
    .TE_B(_0321_),
    .Z(io_out[18]));
 sky130_fd_sc_hd__ebufn_8 _1052_ (.A(\frequency_counter_0.dbg_state[1] ),
    .TE_B(_0322_),
    .Z(io_out[19]));
 sky130_fd_sc_hd__ebufn_8 _1053_ (.A(\frequency_counter_0.clk_counter[9] ),
    .TE_B(_0323_),
    .Z(io_out[20]));
 sky130_fd_sc_hd__ebufn_8 _1054_ (.A(\frequency_counter_0.clk_counter[10] ),
    .TE_B(_0324_),
    .Z(io_out[21]));
 sky130_fd_sc_hd__ebufn_8 _1055_ (.A(\frequency_counter_0.clk_counter[11] ),
    .TE_B(_0325_),
    .Z(io_out[22]));
 sky130_fd_sc_hd__ebufn_8 _1056_ (.A(\frequency_counter_0.dbg_edge_count[0] ),
    .TE_B(_0326_),
    .Z(io_out[23]));
 sky130_fd_sc_hd__ebufn_8 _1057_ (.A(\frequency_counter_0.dbg_edge_count[1] ),
    .TE_B(_0327_),
    .Z(io_out[24]));
 sky130_fd_sc_hd__ebufn_8 _1058_ (.A(\frequency_counter_0.dbg_edge_count[2] ),
    .TE_B(_0328_),
    .Z(io_out[25]));
 sky130_fd_sc_hd__ebufn_8 _1059_ (.A(net58),
    .TE_B(_0329_),
    .Z(io_out[26]));
 sky130_fd_sc_hd__ebufn_8 _1060_ (.A(net59),
    .TE_B(_0330_),
    .Z(io_out[27]));
 sky130_fd_sc_hd__ebufn_8 _1061_ (.A(net60),
    .TE_B(_0331_),
    .Z(io_out[28]));
 sky130_fd_sc_hd__ebufn_8 _1062_ (.A(net61),
    .TE_B(_0332_),
    .Z(io_out[29]));
 sky130_fd_sc_hd__ebufn_8 _1063_ (.A(net62),
    .TE_B(_0333_),
    .Z(io_out[30]));
 sky130_fd_sc_hd__ebufn_8 _1064_ (.A(net63),
    .TE_B(_0334_),
    .Z(io_out[31]));
 sky130_fd_sc_hd__ebufn_8 _1065_ (.A(net64),
    .TE_B(_0335_),
    .Z(io_out[32]));
 sky130_fd_sc_hd__ebufn_8 _1066_ (.A(net65),
    .TE_B(_0336_),
    .Z(io_out[33]));
 sky130_fd_sc_hd__ebufn_8 _1067_ (.A(net66),
    .TE_B(_0337_),
    .Z(io_out[34]));
 sky130_fd_sc_hd__ebufn_8 _1068_ (.A(net67),
    .TE_B(_0338_),
    .Z(io_out[35]));
 sky130_fd_sc_hd__ebufn_8 _1069_ (.A(net68),
    .TE_B(_0339_),
    .Z(io_out[36]));
 sky130_fd_sc_hd__ebufn_8 _1070_ (.A(net69),
    .TE_B(_0340_),
    .Z(io_out[37]));
 sky130_fd_sc_hd__ebufn_8 _1071_ (.A(net70),
    .TE_B(_0341_),
    .Z(io_oeb[0]));
 sky130_fd_sc_hd__ebufn_8 _1072_ (.A(net71),
    .TE_B(_0342_),
    .Z(io_oeb[1]));
 sky130_fd_sc_hd__ebufn_8 _1073_ (.A(net72),
    .TE_B(_0343_),
    .Z(io_oeb[2]));
 sky130_fd_sc_hd__ebufn_8 _1074_ (.A(net73),
    .TE_B(_0344_),
    .Z(io_oeb[3]));
 sky130_fd_sc_hd__ebufn_8 _1075_ (.A(net74),
    .TE_B(_0345_),
    .Z(io_oeb[4]));
 sky130_fd_sc_hd__ebufn_8 _1076_ (.A(net75),
    .TE_B(_0346_),
    .Z(io_oeb[5]));
 sky130_fd_sc_hd__ebufn_8 _1077_ (.A(net76),
    .TE_B(_0347_),
    .Z(io_oeb[6]));
 sky130_fd_sc_hd__ebufn_8 _1078_ (.A(net77),
    .TE_B(_0348_),
    .Z(io_oeb[7]));
 sky130_fd_sc_hd__ebufn_8 _1079_ (.A(net78),
    .TE_B(_0349_),
    .Z(io_oeb[8]));
 sky130_fd_sc_hd__ebufn_8 _1080_ (.A(net79),
    .TE_B(_0350_),
    .Z(io_oeb[9]));
 sky130_fd_sc_hd__ebufn_8 _1081_ (.A(net80),
    .TE_B(_0351_),
    .Z(io_oeb[10]));
 sky130_fd_sc_hd__ebufn_8 _1082_ (.A(net81),
    .TE_B(_0352_),
    .Z(io_oeb[11]));
 sky130_fd_sc_hd__ebufn_8 _1083_ (.A(net82),
    .TE_B(_0353_),
    .Z(io_oeb[12]));
 sky130_fd_sc_hd__ebufn_8 _1084_ (.A(net83),
    .TE_B(_0354_),
    .Z(io_oeb[13]));
 sky130_fd_sc_hd__ebufn_8 _1085_ (.A(net84),
    .TE_B(_0355_),
    .Z(io_oeb[14]));
 sky130_fd_sc_hd__ebufn_8 _1086_ (.A(net85),
    .TE_B(_0356_),
    .Z(io_oeb[15]));
 sky130_fd_sc_hd__ebufn_8 _1087_ (.A(net86),
    .TE_B(_0357_),
    .Z(io_oeb[16]));
 sky130_fd_sc_hd__ebufn_8 _1088_ (.A(net87),
    .TE_B(_0358_),
    .Z(io_oeb[17]));
 sky130_fd_sc_hd__ebufn_8 _1089_ (.A(net88),
    .TE_B(_0359_),
    .Z(io_oeb[18]));
 sky130_fd_sc_hd__ebufn_8 _1090_ (.A(net89),
    .TE_B(_0360_),
    .Z(io_oeb[19]));
 sky130_fd_sc_hd__ebufn_8 _1091_ (.A(net90),
    .TE_B(_0361_),
    .Z(io_oeb[20]));
 sky130_fd_sc_hd__ebufn_8 _1092_ (.A(net91),
    .TE_B(_0362_),
    .Z(io_oeb[21]));
 sky130_fd_sc_hd__ebufn_8 _1093_ (.A(net92),
    .TE_B(_0363_),
    .Z(io_oeb[22]));
 sky130_fd_sc_hd__ebufn_8 _1094_ (.A(net93),
    .TE_B(_0364_),
    .Z(io_oeb[23]));
 sky130_fd_sc_hd__ebufn_8 _1095_ (.A(net94),
    .TE_B(_0365_),
    .Z(io_oeb[24]));
 sky130_fd_sc_hd__ebufn_8 _1096_ (.A(net95),
    .TE_B(_0366_),
    .Z(io_oeb[25]));
 sky130_fd_sc_hd__ebufn_8 _1097_ (.A(net96),
    .TE_B(_0367_),
    .Z(io_oeb[26]));
 sky130_fd_sc_hd__ebufn_8 _1098_ (.A(net97),
    .TE_B(_0368_),
    .Z(io_oeb[27]));
 sky130_fd_sc_hd__ebufn_8 _1099_ (.A(net98),
    .TE_B(_0369_),
    .Z(io_oeb[28]));
 sky130_fd_sc_hd__ebufn_8 _1100_ (.A(net99),
    .TE_B(_0370_),
    .Z(io_oeb[29]));
 sky130_fd_sc_hd__ebufn_8 _1101_ (.A(net100),
    .TE_B(_0371_),
    .Z(io_oeb[30]));
 sky130_fd_sc_hd__ebufn_8 _1102_ (.A(net101),
    .TE_B(_0372_),
    .Z(io_oeb[31]));
 sky130_fd_sc_hd__ebufn_8 _1103_ (.A(net102),
    .TE_B(_0373_),
    .Z(io_oeb[32]));
 sky130_fd_sc_hd__ebufn_8 _1104_ (.A(net103),
    .TE_B(_0374_),
    .Z(io_oeb[33]));
 sky130_fd_sc_hd__ebufn_8 _1105_ (.A(net104),
    .TE_B(_0375_),
    .Z(io_oeb[34]));
 sky130_fd_sc_hd__ebufn_8 _1106_ (.A(net105),
    .TE_B(_0376_),
    .Z(io_oeb[35]));
 sky130_fd_sc_hd__ebufn_8 _1107_ (.A(net106),
    .TE_B(_0377_),
    .Z(io_oeb[36]));
 sky130_fd_sc_hd__ebufn_8 _1108_ (.A(net107),
    .TE_B(_0378_),
    .Z(io_oeb[37]));
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__decap_3 PHY_162 ();
 sky130_fd_sc_hd__decap_3 PHY_163 ();
 sky130_fd_sc_hd__decap_3 PHY_164 ();
 sky130_fd_sc_hd__decap_3 PHY_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__clkbuf_1 input1 (.A(active),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(io_in[8]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(la1_data_in[0]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(la1_data_in[10]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(la1_data_in[11]),
    .X(net5));
 sky130_fd_sc_hd__dlymetal6s2s_1 input6 (.A(la1_data_in[12]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_1 input7 (.A(la1_data_in[13]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_2 input8 (.A(la1_data_in[1]),
    .X(net8));
 sky130_fd_sc_hd__dlymetal6s2s_1 input9 (.A(la1_data_in[2]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_1 input10 (.A(la1_data_in[3]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_1 input11 (.A(la1_data_in[4]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_1 input12 (.A(la1_data_in[5]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_1 input13 (.A(la1_data_in[6]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_1 input14 (.A(la1_data_in[7]),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_1 input15 (.A(la1_data_in[8]),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_1 input16 (.A(la1_data_in[9]),
    .X(net16));
 sky130_fd_sc_hd__conb_1 _1001__17 (.LO(net17));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_0__f_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_2_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_1__f_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_2_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_2__f_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_2_2__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_3__f_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_2_3__leaf_wb_clk_i));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1 (.A(\frequency_counter_0.edge_detect0.q0 ),
    .X(net108));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(\frequency_counter_0.edge_detect0.q1 ),
    .X(net109));
 sky130_fd_sc_hd__decap_4 FILLER_0_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_28 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_84 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_192 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_71 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_10 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_24 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_87 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_99 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_268 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_227 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_45 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_291 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_13 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_36 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_291 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_58 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_267 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_10 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_260 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_297 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_12 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_36 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_28 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_77 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_124 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_155 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_272 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_240 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_236 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_296 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_286 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_170 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_235 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_180 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_238 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_10 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_155 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_187 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_229 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_244 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_286 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_244 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_183 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_210 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_188 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_286 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_174 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_259 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_298 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_228 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_235 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_170 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_163 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_234 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_206 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_267 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_260 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_230 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_267 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_272 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_168 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_224 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_243 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_295 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_43 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_213 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_155 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_291 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_43 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_296 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_174 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_182 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_239 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_286 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_210 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_217 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_40 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_248 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_268 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_171 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_236 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_258 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_183 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_286 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_17 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_157 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_182 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_297 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_12 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_185 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_10 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_182 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_297 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_13 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_16 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_298 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_13 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_286 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_20 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_100 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_52 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_72 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_107 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_146 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_186 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_190 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_126 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_207 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_286 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_13 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_62 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_298 ();
endmodule

