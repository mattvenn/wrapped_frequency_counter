// This is the unpowered netlist.
module wrapped_frequency_counter (active,
    wb_clk_i,
    io_in,
    io_oeb,
    io_out,
    la1_data_in,
    la1_data_out,
    la1_oenb);
 input active;
 input wb_clk_i;
 input [37:0] io_in;
 output [37:0] io_oeb;
 output [37:0] io_out;
 input [31:0] la1_data_in;
 output [31:0] la1_data_out;
 input [31:0] la1_oenb;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire clknet_0_wb_clk_i;
 wire \frequency_counter_0.clk_counter[0] ;
 wire \frequency_counter_0.clk_counter[10] ;
 wire \frequency_counter_0.clk_counter[11] ;
 wire \frequency_counter_0.clk_counter[1] ;
 wire \frequency_counter_0.clk_counter[2] ;
 wire \frequency_counter_0.clk_counter[3] ;
 wire \frequency_counter_0.clk_counter[4] ;
 wire \frequency_counter_0.clk_counter[5] ;
 wire \frequency_counter_0.clk_counter[6] ;
 wire \frequency_counter_0.clk_counter[7] ;
 wire \frequency_counter_0.clk_counter[8] ;
 wire \frequency_counter_0.clk_counter[9] ;
 wire \frequency_counter_0.digit ;
 wire \frequency_counter_0.edge_counter[0] ;
 wire \frequency_counter_0.edge_counter[1] ;
 wire \frequency_counter_0.edge_counter[2] ;
 wire \frequency_counter_0.edge_counter[3] ;
 wire \frequency_counter_0.edge_counter[4] ;
 wire \frequency_counter_0.edge_counter[5] ;
 wire \frequency_counter_0.edge_counter[6] ;
 wire \frequency_counter_0.edge_detect0.q0 ;
 wire \frequency_counter_0.edge_detect0.q1 ;
 wire \frequency_counter_0.edge_detect0.q2 ;
 wire \frequency_counter_0.segments[0] ;
 wire \frequency_counter_0.segments[1] ;
 wire \frequency_counter_0.segments[2] ;
 wire \frequency_counter_0.segments[3] ;
 wire \frequency_counter_0.segments[4] ;
 wire \frequency_counter_0.segments[5] ;
 wire \frequency_counter_0.segments[6] ;
 wire \frequency_counter_0.seven_segment0.load ;
 wire \frequency_counter_0.seven_segment0.ten_count[0] ;
 wire \frequency_counter_0.seven_segment0.ten_count[1] ;
 wire \frequency_counter_0.seven_segment0.ten_count[2] ;
 wire \frequency_counter_0.seven_segment0.ten_count[3] ;
 wire \frequency_counter_0.seven_segment0.ten_count_reg[0] ;
 wire \frequency_counter_0.seven_segment0.ten_count_reg[1] ;
 wire \frequency_counter_0.seven_segment0.ten_count_reg[2] ;
 wire \frequency_counter_0.seven_segment0.ten_count_reg[3] ;
 wire \frequency_counter_0.seven_segment0.unit_count[0] ;
 wire \frequency_counter_0.seven_segment0.unit_count[1] ;
 wire \frequency_counter_0.seven_segment0.unit_count[2] ;
 wire \frequency_counter_0.seven_segment0.unit_count[3] ;
 wire \frequency_counter_0.seven_segment0.unit_count_reg[0] ;
 wire \frequency_counter_0.seven_segment0.unit_count_reg[1] ;
 wire \frequency_counter_0.seven_segment0.unit_count_reg[2] ;
 wire \frequency_counter_0.seven_segment0.unit_count_reg[3] ;
 wire \frequency_counter_0.state[0] ;
 wire \frequency_counter_0.state[1] ;
 wire \frequency_counter_0.state[2] ;
 wire \frequency_counter_0.update_period[0] ;
 wire \frequency_counter_0.update_period[10] ;
 wire \frequency_counter_0.update_period[11] ;
 wire \frequency_counter_0.update_period[1] ;
 wire \frequency_counter_0.update_period[2] ;
 wire \frequency_counter_0.update_period[3] ;
 wire \frequency_counter_0.update_period[4] ;
 wire \frequency_counter_0.update_period[5] ;
 wire \frequency_counter_0.update_period[6] ;
 wire \frequency_counter_0.update_period[7] ;
 wire \frequency_counter_0.update_period[8] ;
 wire \frequency_counter_0.update_period[9] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire clknet_2_0__leaf_wb_clk_i;
 wire clknet_2_1__leaf_wb_clk_i;
 wire clknet_2_2__leaf_wb_clk_i;
 wire clknet_2_3__leaf_wb_clk_i;
 wire net117;
 wire net118;

 sky130_fd_sc_hd__clkbuf_8 _0475_ (.A(net1),
    .X(_0052_));
 sky130_fd_sc_hd__buf_8 _0476_ (.A(_0052_),
    .X(_0053_));
 sky130_fd_sc_hd__buf_8 _0477_ (.A(_0053_),
    .X(_0054_));
 sky130_fd_sc_hd__inv_2 _0478_ (.A(_0054_),
    .Y(_0373_));
 sky130_fd_sc_hd__inv_2 _0479_ (.A(_0054_),
    .Y(_0372_));
 sky130_fd_sc_hd__inv_2 _0480_ (.A(_0054_),
    .Y(_0371_));
 sky130_fd_sc_hd__inv_2 _0481_ (.A(_0054_),
    .Y(_0370_));
 sky130_fd_sc_hd__inv_2 _0482_ (.A(_0054_),
    .Y(_0369_));
 sky130_fd_sc_hd__inv_2 _0483_ (.A(_0054_),
    .Y(_0368_));
 sky130_fd_sc_hd__inv_2 _0484_ (.A(_0054_),
    .Y(_0367_));
 sky130_fd_sc_hd__inv_2 _0485_ (.A(_0054_),
    .Y(_0366_));
 sky130_fd_sc_hd__inv_2 _0486_ (.A(_0054_),
    .Y(_0365_));
 sky130_fd_sc_hd__inv_2 _0487_ (.A(_0054_),
    .Y(_0364_));
 sky130_fd_sc_hd__buf_8 _0488_ (.A(_0053_),
    .X(_0055_));
 sky130_fd_sc_hd__inv_2 _0489_ (.A(_0055_),
    .Y(_0363_));
 sky130_fd_sc_hd__inv_2 _0490_ (.A(_0055_),
    .Y(_0362_));
 sky130_fd_sc_hd__inv_2 _0491_ (.A(_0055_),
    .Y(_0361_));
 sky130_fd_sc_hd__inv_2 _0492_ (.A(_0055_),
    .Y(_0360_));
 sky130_fd_sc_hd__inv_2 _0493_ (.A(_0055_),
    .Y(_0359_));
 sky130_fd_sc_hd__inv_2 _0494_ (.A(_0055_),
    .Y(_0358_));
 sky130_fd_sc_hd__inv_2 _0495_ (.A(_0055_),
    .Y(_0357_));
 sky130_fd_sc_hd__inv_2 _0496_ (.A(_0055_),
    .Y(_0356_));
 sky130_fd_sc_hd__inv_2 _0497_ (.A(_0055_),
    .Y(_0355_));
 sky130_fd_sc_hd__inv_2 _0498_ (.A(_0055_),
    .Y(_0354_));
 sky130_fd_sc_hd__buf_8 _0499_ (.A(_0052_),
    .X(_0056_));
 sky130_fd_sc_hd__inv_2 _0500_ (.A(_0056_),
    .Y(_0353_));
 sky130_fd_sc_hd__inv_2 _0501_ (.A(_0056_),
    .Y(_0352_));
 sky130_fd_sc_hd__inv_2 _0502_ (.A(_0056_),
    .Y(_0351_));
 sky130_fd_sc_hd__inv_2 _0503_ (.A(_0056_),
    .Y(_0350_));
 sky130_fd_sc_hd__inv_2 _0504_ (.A(_0056_),
    .Y(_0349_));
 sky130_fd_sc_hd__inv_2 _0505_ (.A(_0056_),
    .Y(_0348_));
 sky130_fd_sc_hd__inv_2 _0506_ (.A(_0056_),
    .Y(_0347_));
 sky130_fd_sc_hd__inv_2 _0507_ (.A(_0056_),
    .Y(_0346_));
 sky130_fd_sc_hd__inv_2 _0508_ (.A(_0056_),
    .Y(_0345_));
 sky130_fd_sc_hd__inv_2 _0509_ (.A(_0056_),
    .Y(_0344_));
 sky130_fd_sc_hd__buf_8 _0510_ (.A(_0052_),
    .X(_0057_));
 sky130_fd_sc_hd__inv_2 _0511_ (.A(_0057_),
    .Y(_0343_));
 sky130_fd_sc_hd__inv_2 _0512_ (.A(_0057_),
    .Y(_0342_));
 sky130_fd_sc_hd__inv_2 _0513_ (.A(_0057_),
    .Y(_0341_));
 sky130_fd_sc_hd__inv_2 _0514_ (.A(_0057_),
    .Y(_0340_));
 sky130_fd_sc_hd__inv_2 _0515_ (.A(_0057_),
    .Y(_0339_));
 sky130_fd_sc_hd__inv_2 _0516_ (.A(_0057_),
    .Y(_0338_));
 sky130_fd_sc_hd__inv_2 _0517_ (.A(_0057_),
    .Y(_0336_));
 sky130_fd_sc_hd__inv_2 _0518_ (.A(_0057_),
    .Y(_0335_));
 sky130_fd_sc_hd__inv_2 _0519_ (.A(_0057_),
    .Y(_0334_));
 sky130_fd_sc_hd__inv_2 _0520_ (.A(_0057_),
    .Y(_0333_));
 sky130_fd_sc_hd__buf_8 _0521_ (.A(_0052_),
    .X(_0058_));
 sky130_fd_sc_hd__inv_2 _0522_ (.A(_0058_),
    .Y(_0325_));
 sky130_fd_sc_hd__inv_2 _0523_ (.A(_0058_),
    .Y(_0326_));
 sky130_fd_sc_hd__inv_2 _0524_ (.A(_0058_),
    .Y(_0327_));
 sky130_fd_sc_hd__inv_2 _0525_ (.A(_0058_),
    .Y(_0328_));
 sky130_fd_sc_hd__inv_2 _0526_ (.A(_0058_),
    .Y(_0329_));
 sky130_fd_sc_hd__inv_2 _0527_ (.A(_0058_),
    .Y(_0330_));
 sky130_fd_sc_hd__inv_2 _0528_ (.A(_0058_),
    .Y(_0331_));
 sky130_fd_sc_hd__inv_2 _0529_ (.A(_0058_),
    .Y(_0276_));
 sky130_fd_sc_hd__inv_2 _0530_ (.A(_0058_),
    .Y(_0283_));
 sky130_fd_sc_hd__inv_2 _0531_ (.A(_0058_),
    .Y(_0287_));
 sky130_fd_sc_hd__buf_6 _0532_ (.A(_0052_),
    .X(_0059_));
 sky130_fd_sc_hd__inv_2 _0533_ (.A(_0059_),
    .Y(_0311_));
 sky130_fd_sc_hd__inv_2 _0534_ (.A(_0059_),
    .Y(_0312_));
 sky130_fd_sc_hd__inv_2 _0535_ (.A(_0059_),
    .Y(_0313_));
 sky130_fd_sc_hd__inv_2 _0536_ (.A(_0059_),
    .Y(_0267_));
 sky130_fd_sc_hd__inv_2 _0537_ (.A(_0059_),
    .Y(_0268_));
 sky130_fd_sc_hd__inv_2 _0538_ (.A(_0059_),
    .Y(_0269_));
 sky130_fd_sc_hd__inv_2 _0539_ (.A(_0059_),
    .Y(_0270_));
 sky130_fd_sc_hd__inv_2 _0540_ (.A(_0059_),
    .Y(_0271_));
 sky130_fd_sc_hd__inv_2 _0541_ (.A(_0059_),
    .Y(_0272_));
 sky130_fd_sc_hd__inv_2 _0542_ (.A(_0059_),
    .Y(_0273_));
 sky130_fd_sc_hd__buf_8 _0543_ (.A(_0052_),
    .X(_0060_));
 sky130_fd_sc_hd__inv_2 _0544_ (.A(_0060_),
    .Y(_0274_));
 sky130_fd_sc_hd__inv_2 _0545_ (.A(_0060_),
    .Y(_0275_));
 sky130_fd_sc_hd__inv_2 _0546_ (.A(_0060_),
    .Y(_0314_));
 sky130_fd_sc_hd__inv_2 _0547_ (.A(_0060_),
    .Y(_0288_));
 sky130_fd_sc_hd__inv_2 _0548_ (.A(_0060_),
    .Y(_0289_));
 sky130_fd_sc_hd__inv_2 _0549_ (.A(_0060_),
    .Y(_0315_));
 sky130_fd_sc_hd__inv_2 _0550_ (.A(_0060_),
    .Y(_0290_));
 sky130_fd_sc_hd__inv_2 _0551_ (.A(_0060_),
    .Y(_0291_));
 sky130_fd_sc_hd__inv_2 _0552_ (.A(_0060_),
    .Y(_0316_));
 sky130_fd_sc_hd__inv_2 _0553_ (.A(_0060_),
    .Y(_0292_));
 sky130_fd_sc_hd__buf_8 _0554_ (.A(_0052_),
    .X(_0061_));
 sky130_fd_sc_hd__inv_2 _0555_ (.A(_0061_),
    .Y(_0293_));
 sky130_fd_sc_hd__inv_2 _0556_ (.A(_0061_),
    .Y(_0317_));
 sky130_fd_sc_hd__inv_2 _0557_ (.A(_0061_),
    .Y(_0294_));
 sky130_fd_sc_hd__inv_2 _0558_ (.A(_0061_),
    .Y(_0295_));
 sky130_fd_sc_hd__inv_2 _0559_ (.A(_0061_),
    .Y(_0318_));
 sky130_fd_sc_hd__inv_2 _0560_ (.A(_0061_),
    .Y(_0296_));
 sky130_fd_sc_hd__inv_2 _0561_ (.A(_0061_),
    .Y(_0297_));
 sky130_fd_sc_hd__inv_2 _0562_ (.A(_0061_),
    .Y(_0319_));
 sky130_fd_sc_hd__inv_2 _0563_ (.A(_0061_),
    .Y(_0320_));
 sky130_fd_sc_hd__inv_2 _0564_ (.A(_0061_),
    .Y(_0324_));
 sky130_fd_sc_hd__buf_8 _0565_ (.A(_0052_),
    .X(_0062_));
 sky130_fd_sc_hd__inv_2 _0566_ (.A(_0062_),
    .Y(_0298_));
 sky130_fd_sc_hd__inv_2 _0567_ (.A(_0062_),
    .Y(_0300_));
 sky130_fd_sc_hd__inv_2 _0568_ (.A(_0062_),
    .Y(_0301_));
 sky130_fd_sc_hd__inv_2 _0569_ (.A(_0062_),
    .Y(_0302_));
 sky130_fd_sc_hd__inv_2 _0570_ (.A(_0062_),
    .Y(_0321_));
 sky130_fd_sc_hd__inv_2 _0571_ (.A(_0062_),
    .Y(_0303_));
 sky130_fd_sc_hd__inv_2 _0572_ (.A(_0062_),
    .Y(_0322_));
 sky130_fd_sc_hd__inv_2 _0573_ (.A(_0062_),
    .Y(_0304_));
 sky130_fd_sc_hd__inv_2 _0574_ (.A(_0062_),
    .Y(_0305_));
 sky130_fd_sc_hd__inv_2 _0575_ (.A(_0062_),
    .Y(_0306_));
 sky130_fd_sc_hd__buf_8 _0576_ (.A(_0052_),
    .X(_0063_));
 sky130_fd_sc_hd__inv_2 _0577_ (.A(_0063_),
    .Y(_0307_));
 sky130_fd_sc_hd__inv_2 _0578_ (.A(_0063_),
    .Y(_0308_));
 sky130_fd_sc_hd__inv_2 _0579_ (.A(_0063_),
    .Y(_0309_));
 sky130_fd_sc_hd__inv_2 _0580_ (.A(_0063_),
    .Y(_0310_));
 sky130_fd_sc_hd__inv_2 _0581_ (.A(_0063_),
    .Y(_0323_));
 sky130_fd_sc_hd__inv_2 _0582_ (.A(_0063_),
    .Y(_0277_));
 sky130_fd_sc_hd__inv_2 _0583_ (.A(_0063_),
    .Y(_0278_));
 sky130_fd_sc_hd__inv_2 _0584_ (.A(_0063_),
    .Y(_0279_));
 sky130_fd_sc_hd__inv_2 _0585_ (.A(_0063_),
    .Y(_0280_));
 sky130_fd_sc_hd__inv_2 _0586_ (.A(_0063_),
    .Y(_0281_));
 sky130_fd_sc_hd__inv_2 _0587_ (.A(_0053_),
    .Y(_0282_));
 sky130_fd_sc_hd__inv_2 _0588_ (.A(_0053_),
    .Y(_0285_));
 sky130_fd_sc_hd__inv_2 _0589_ (.A(_0053_),
    .Y(_0286_));
 sky130_fd_sc_hd__inv_2 _0590_ (.A(_0053_),
    .Y(_0284_));
 sky130_fd_sc_hd__inv_2 _0591_ (.A(_0053_),
    .Y(_0332_));
 sky130_fd_sc_hd__inv_2 _0592_ (.A(_0053_),
    .Y(_0337_));
 sky130_fd_sc_hd__inv_2 _0593_ (.A(_0053_),
    .Y(_0299_));
 sky130_fd_sc_hd__clkbuf_4 _0594_ (.A(net3),
    .X(_0064_));
 sky130_fd_sc_hd__clkbuf_4 _0595_ (.A(_0064_),
    .X(_0065_));
 sky130_fd_sc_hd__clkbuf_4 _0596_ (.A(\frequency_counter_0.state[0] ),
    .X(_0066_));
 sky130_fd_sc_hd__inv_2 _0597_ (.A(\frequency_counter_0.clk_counter[6] ),
    .Y(_0067_));
 sky130_fd_sc_hd__inv_2 _0598_ (.A(\frequency_counter_0.clk_counter[5] ),
    .Y(_0068_));
 sky130_fd_sc_hd__a22oi_1 _0599_ (.A1(_0067_),
    .A2(\frequency_counter_0.update_period[6] ),
    .B1(\frequency_counter_0.update_period[5] ),
    .B2(_0068_),
    .Y(_0069_));
 sky130_fd_sc_hd__inv_2 _0600_ (.A(\frequency_counter_0.update_period[1] ),
    .Y(_0070_));
 sky130_fd_sc_hd__inv_2 _0601_ (.A(\frequency_counter_0.update_period[0] ),
    .Y(_0071_));
 sky130_fd_sc_hd__a211o_1 _0602_ (.A1(\frequency_counter_0.clk_counter[1] ),
    .A2(_0070_),
    .B1(_0071_),
    .C1(\frequency_counter_0.clk_counter[0] ),
    .X(_0072_));
 sky130_fd_sc_hd__inv_2 _0603_ (.A(\frequency_counter_0.update_period[2] ),
    .Y(_0073_));
 sky130_fd_sc_hd__o22a_1 _0604_ (.A1(\frequency_counter_0.clk_counter[2] ),
    .A2(_0073_),
    .B1(_0070_),
    .B2(\frequency_counter_0.clk_counter[1] ),
    .X(_0074_));
 sky130_fd_sc_hd__inv_2 _0605_ (.A(\frequency_counter_0.update_period[3] ),
    .Y(_0075_));
 sky130_fd_sc_hd__a22o_1 _0606_ (.A1(\frequency_counter_0.clk_counter[3] ),
    .A2(_0075_),
    .B1(_0073_),
    .B2(\frequency_counter_0.clk_counter[2] ),
    .X(_0076_));
 sky130_fd_sc_hd__a21o_1 _0607_ (.A1(_0072_),
    .A2(_0074_),
    .B1(_0076_),
    .X(_0077_));
 sky130_fd_sc_hd__inv_2 _0608_ (.A(\frequency_counter_0.clk_counter[7] ),
    .Y(_0078_));
 sky130_fd_sc_hd__o22a_1 _0609_ (.A1(_0078_),
    .A2(\frequency_counter_0.update_period[7] ),
    .B1(\frequency_counter_0.update_period[6] ),
    .B2(_0067_),
    .X(_0079_));
 sky130_fd_sc_hd__inv_2 _0610_ (.A(\frequency_counter_0.clk_counter[4] ),
    .Y(_0080_));
 sky130_fd_sc_hd__o22a_1 _0611_ (.A1(_0068_),
    .A2(\frequency_counter_0.update_period[5] ),
    .B1(\frequency_counter_0.update_period[4] ),
    .B2(_0080_),
    .X(_0081_));
 sky130_fd_sc_hd__inv_2 _0612_ (.A(\frequency_counter_0.update_period[4] ),
    .Y(_0082_));
 sky130_fd_sc_hd__or2b_1 _0613_ (.A(\frequency_counter_0.clk_counter[7] ),
    .B_N(\frequency_counter_0.update_period[7] ),
    .X(_0083_));
 sky130_fd_sc_hd__o221a_1 _0614_ (.A1(\frequency_counter_0.clk_counter[4] ),
    .A2(_0082_),
    .B1(_0075_),
    .B2(\frequency_counter_0.clk_counter[3] ),
    .C1(_0083_),
    .X(_0084_));
 sky130_fd_sc_hd__and3_1 _0615_ (.A(_0079_),
    .B(_0081_),
    .C(_0084_),
    .X(_0085_));
 sky130_fd_sc_hd__a22o_1 _0616_ (.A1(_0067_),
    .A2(\frequency_counter_0.update_period[6] ),
    .B1(\frequency_counter_0.update_period[5] ),
    .B2(_0068_),
    .X(_0086_));
 sky130_fd_sc_hd__o21ai_1 _0617_ (.A1(_0086_),
    .A2(_0081_),
    .B1(_0079_),
    .Y(_0087_));
 sky130_fd_sc_hd__a32o_1 _0618_ (.A1(_0069_),
    .A2(_0077_),
    .A3(_0085_),
    .B1(_0087_),
    .B2(_0083_),
    .X(_0088_));
 sky130_fd_sc_hd__inv_2 _0619_ (.A(\frequency_counter_0.clk_counter[10] ),
    .Y(_0089_));
 sky130_fd_sc_hd__inv_2 _0620_ (.A(\frequency_counter_0.clk_counter[9] ),
    .Y(_0090_));
 sky130_fd_sc_hd__and2_1 _0621_ (.A(_0090_),
    .B(\frequency_counter_0.update_period[9] ),
    .X(_0091_));
 sky130_fd_sc_hd__inv_2 _0622_ (.A(\frequency_counter_0.clk_counter[8] ),
    .Y(_0092_));
 sky130_fd_sc_hd__or2b_1 _0623_ (.A(\frequency_counter_0.clk_counter[11] ),
    .B_N(\frequency_counter_0.update_period[11] ),
    .X(_0093_));
 sky130_fd_sc_hd__a21bo_1 _0624_ (.A1(_0092_),
    .A2(\frequency_counter_0.update_period[8] ),
    .B1_N(_0093_),
    .X(_0094_));
 sky130_fd_sc_hd__a211oi_1 _0625_ (.A1(_0089_),
    .A2(\frequency_counter_0.update_period[10] ),
    .B1(_0091_),
    .C1(_0094_),
    .Y(_0095_));
 sky130_fd_sc_hd__inv_2 _0626_ (.A(\frequency_counter_0.clk_counter[11] ),
    .Y(_0096_));
 sky130_fd_sc_hd__o22a_1 _0627_ (.A1(_0096_),
    .A2(\frequency_counter_0.update_period[11] ),
    .B1(\frequency_counter_0.update_period[10] ),
    .B2(_0089_),
    .X(_0097_));
 sky130_fd_sc_hd__o22a_1 _0628_ (.A1(_0090_),
    .A2(\frequency_counter_0.update_period[9] ),
    .B1(\frequency_counter_0.update_period[8] ),
    .B2(_0092_),
    .X(_0098_));
 sky130_fd_sc_hd__and3_1 _0629_ (.A(_0095_),
    .B(_0097_),
    .C(_0098_),
    .X(_0099_));
 sky130_fd_sc_hd__a211o_1 _0630_ (.A1(_0089_),
    .A2(\frequency_counter_0.update_period[10] ),
    .B1(_0091_),
    .C1(_0098_),
    .X(_0100_));
 sky130_fd_sc_hd__a21boi_2 _0631_ (.A1(_0097_),
    .A2(_0100_),
    .B1_N(_0093_),
    .Y(_0101_));
 sky130_fd_sc_hd__a21o_1 _0632_ (.A1(_0088_),
    .A2(_0099_),
    .B1(_0101_),
    .X(_0102_));
 sky130_fd_sc_hd__buf_2 _0633_ (.A(\frequency_counter_0.edge_counter[1] ),
    .X(_0103_));
 sky130_fd_sc_hd__o21a_1 _0634_ (.A1(\frequency_counter_0.edge_counter[2] ),
    .A2(_0103_),
    .B1(\frequency_counter_0.edge_counter[3] ),
    .X(_0104_));
 sky130_fd_sc_hd__or3_1 _0635_ (.A(\frequency_counter_0.edge_counter[5] ),
    .B(\frequency_counter_0.edge_counter[4] ),
    .C(_0104_),
    .X(_0105_));
 sky130_fd_sc_hd__o21a_1 _0636_ (.A1(\frequency_counter_0.edge_counter[6] ),
    .A2(_0105_),
    .B1(\frequency_counter_0.state[2] ),
    .X(_0106_));
 sky130_fd_sc_hd__a21oi_1 _0637_ (.A1(_0066_),
    .A2(_0102_),
    .B1(_0106_),
    .Y(_0107_));
 sky130_fd_sc_hd__nor2_1 _0638_ (.A(_0065_),
    .B(_0107_),
    .Y(_0002_));
 sky130_fd_sc_hd__inv_2 _0639_ (.A(\frequency_counter_0.state[0] ),
    .Y(_0108_));
 sky130_fd_sc_hd__a211o_2 _0640_ (.A1(_0088_),
    .A2(_0099_),
    .B1(_0101_),
    .C1(_0108_),
    .X(_0109_));
 sky130_fd_sc_hd__buf_2 _0641_ (.A(_0109_),
    .X(_0110_));
 sky130_fd_sc_hd__or3b_1 _0642_ (.A(\frequency_counter_0.state[1] ),
    .B(_0064_),
    .C_N(_0110_),
    .X(_0111_));
 sky130_fd_sc_hd__clkbuf_1 _0643_ (.A(_0111_),
    .X(_0001_));
 sky130_fd_sc_hd__mux2_2 _0644_ (.A0(\frequency_counter_0.seven_segment0.unit_count_reg[3] ),
    .A1(\frequency_counter_0.seven_segment0.ten_count_reg[3] ),
    .S(\frequency_counter_0.digit ),
    .X(_0112_));
 sky130_fd_sc_hd__inv_2 _0645_ (.A(_0112_),
    .Y(_0113_));
 sky130_fd_sc_hd__mux2_1 _0646_ (.A0(\frequency_counter_0.seven_segment0.unit_count_reg[2] ),
    .A1(\frequency_counter_0.seven_segment0.ten_count_reg[2] ),
    .S(\frequency_counter_0.digit ),
    .X(_0114_));
 sky130_fd_sc_hd__mux2_2 _0647_ (.A0(\frequency_counter_0.seven_segment0.unit_count_reg[0] ),
    .A1(\frequency_counter_0.seven_segment0.ten_count_reg[0] ),
    .S(\frequency_counter_0.digit ),
    .X(_0115_));
 sky130_fd_sc_hd__nor2_1 _0648_ (.A(_0114_),
    .B(_0115_),
    .Y(_0116_));
 sky130_fd_sc_hd__mux2_2 _0649_ (.A0(\frequency_counter_0.seven_segment0.unit_count_reg[1] ),
    .A1(\frequency_counter_0.seven_segment0.ten_count_reg[1] ),
    .S(\frequency_counter_0.digit ),
    .X(_0117_));
 sky130_fd_sc_hd__nor2_1 _0650_ (.A(_0114_),
    .B(_0117_),
    .Y(_0118_));
 sky130_fd_sc_hd__nor2_1 _0651_ (.A(_0118_),
    .B(_0112_),
    .Y(_0119_));
 sky130_fd_sc_hd__and2_1 _0652_ (.A(_0118_),
    .B(_0112_),
    .X(_0120_));
 sky130_fd_sc_hd__a221o_1 _0653_ (.A1(_0113_),
    .A2(_0116_),
    .B1(_0119_),
    .B2(_0115_),
    .C1(_0120_),
    .X(\frequency_counter_0.segments[0] ));
 sky130_fd_sc_hd__a21bo_1 _0654_ (.A1(_0117_),
    .A2(_0115_),
    .B1_N(_0114_),
    .X(_0121_));
 sky130_fd_sc_hd__or2_1 _0655_ (.A(_0117_),
    .B(_0115_),
    .X(_0122_));
 sky130_fd_sc_hd__or2b_1 _0656_ (.A(_0121_),
    .B_N(_0122_),
    .X(_0123_));
 sky130_fd_sc_hd__a21o_1 _0657_ (.A1(_0113_),
    .A2(_0123_),
    .B1(_0120_),
    .X(\frequency_counter_0.segments[1] ));
 sky130_fd_sc_hd__o21bai_2 _0658_ (.A1(_0112_),
    .A2(_0116_),
    .B1_N(_0118_),
    .Y(\frequency_counter_0.segments[2] ));
 sky130_fd_sc_hd__nand2_1 _0659_ (.A(_0114_),
    .B(_0117_),
    .Y(_0124_));
 sky130_fd_sc_hd__a21oi_1 _0660_ (.A1(_0117_),
    .A2(_0113_),
    .B1(_0118_),
    .Y(_0125_));
 sky130_fd_sc_hd__nor2_2 _0661_ (.A(_0115_),
    .B(_0125_),
    .Y(\frequency_counter_0.segments[4] ));
 sky130_fd_sc_hd__a31o_1 _0662_ (.A1(_0119_),
    .A2(_0122_),
    .A3(_0124_),
    .B1(\frequency_counter_0.segments[4] ),
    .X(\frequency_counter_0.segments[3] ));
 sky130_fd_sc_hd__a21oi_1 _0663_ (.A1(_0121_),
    .A2(_0122_),
    .B1(_0112_),
    .Y(_0126_));
 sky130_fd_sc_hd__or2_1 _0664_ (.A(_0120_),
    .B(_0126_),
    .X(_0127_));
 sky130_fd_sc_hd__clkbuf_1 _0665_ (.A(_0127_),
    .X(\frequency_counter_0.segments[5] ));
 sky130_fd_sc_hd__nand3_1 _0666_ (.A(_0114_),
    .B(_0117_),
    .C(_0115_),
    .Y(_0128_));
 sky130_fd_sc_hd__a21o_1 _0667_ (.A1(_0119_),
    .A2(_0128_),
    .B1(_0120_),
    .X(\frequency_counter_0.segments[6] ));
 sky130_fd_sc_hd__clkinv_2 _0668_ (.A(\frequency_counter_0.state[2] ),
    .Y(_0129_));
 sky130_fd_sc_hd__or3_1 _0669_ (.A(\frequency_counter_0.edge_counter[6] ),
    .B(_0129_),
    .C(_0105_),
    .X(_0130_));
 sky130_fd_sc_hd__nor2_1 _0670_ (.A(_0065_),
    .B(_0130_),
    .Y(_0000_));
 sky130_fd_sc_hd__inv_2 _0671_ (.A(_0053_),
    .Y(_0374_));
 sky130_fd_sc_hd__inv_2 _0672_ (.A(_0130_),
    .Y(_0131_));
 sky130_fd_sc_hd__nor2_1 _0673_ (.A(\frequency_counter_0.state[1] ),
    .B(\frequency_counter_0.state[2] ),
    .Y(_0132_));
 sky130_fd_sc_hd__nand2_1 _0674_ (.A(_0066_),
    .B(\frequency_counter_0.edge_detect0.q1 ),
    .Y(_0133_));
 sky130_fd_sc_hd__o22a_2 _0675_ (.A1(_0066_),
    .A2(_0132_),
    .B1(_0133_),
    .B2(\frequency_counter_0.edge_detect0.q2 ),
    .X(_0134_));
 sky130_fd_sc_hd__nor2_4 _0676_ (.A(_0131_),
    .B(_0134_),
    .Y(_0135_));
 sky130_fd_sc_hd__or2_2 _0677_ (.A(\frequency_counter_0.state[1] ),
    .B(\frequency_counter_0.state[2] ),
    .X(_0136_));
 sky130_fd_sc_hd__xnor2_1 _0678_ (.A(\frequency_counter_0.edge_counter[0] ),
    .B(_0103_),
    .Y(_0137_));
 sky130_fd_sc_hd__o221ai_1 _0679_ (.A1(_0103_),
    .A2(_0129_),
    .B1(_0136_),
    .B2(_0137_),
    .C1(_0135_),
    .Y(_0138_));
 sky130_fd_sc_hd__inv_2 _0680_ (.A(net3),
    .Y(_0139_));
 sky130_fd_sc_hd__clkbuf_4 _0681_ (.A(_0139_),
    .X(_0140_));
 sky130_fd_sc_hd__o211a_1 _0682_ (.A1(_0103_),
    .A2(_0135_),
    .B1(_0138_),
    .C1(_0140_),
    .X(_0003_));
 sky130_fd_sc_hd__a21oi_1 _0683_ (.A1(\frequency_counter_0.edge_counter[0] ),
    .A2(_0103_),
    .B1(\frequency_counter_0.edge_counter[2] ),
    .Y(_0141_));
 sky130_fd_sc_hd__and3_1 _0684_ (.A(\frequency_counter_0.edge_counter[0] ),
    .B(\frequency_counter_0.edge_counter[2] ),
    .C(_0103_),
    .X(_0142_));
 sky130_fd_sc_hd__xor2_1 _0685_ (.A(\frequency_counter_0.edge_counter[2] ),
    .B(_0103_),
    .X(_0143_));
 sky130_fd_sc_hd__o32a_1 _0686_ (.A1(_0136_),
    .A2(_0141_),
    .A3(_0142_),
    .B1(_0143_),
    .B2(_0129_),
    .X(_0144_));
 sky130_fd_sc_hd__nand2_1 _0687_ (.A(_0135_),
    .B(_0144_),
    .Y(_0145_));
 sky130_fd_sc_hd__o211a_1 _0688_ (.A1(\frequency_counter_0.edge_counter[2] ),
    .A2(_0135_),
    .B1(_0145_),
    .C1(_0140_),
    .X(_0004_));
 sky130_fd_sc_hd__o21ai_1 _0689_ (.A1(\frequency_counter_0.edge_counter[2] ),
    .A2(_0103_),
    .B1(\frequency_counter_0.edge_counter[3] ),
    .Y(_0146_));
 sky130_fd_sc_hd__or3_1 _0690_ (.A(\frequency_counter_0.edge_counter[3] ),
    .B(\frequency_counter_0.edge_counter[2] ),
    .C(_0103_),
    .X(_0147_));
 sky130_fd_sc_hd__or2_1 _0691_ (.A(\frequency_counter_0.edge_counter[3] ),
    .B(_0142_),
    .X(_0148_));
 sky130_fd_sc_hd__and2_1 _0692_ (.A(\frequency_counter_0.edge_counter[3] ),
    .B(_0142_),
    .X(_0149_));
 sky130_fd_sc_hd__nor2_1 _0693_ (.A(_0136_),
    .B(_0149_),
    .Y(_0150_));
 sky130_fd_sc_hd__a32o_1 _0694_ (.A1(\frequency_counter_0.state[2] ),
    .A2(_0146_),
    .A3(_0147_),
    .B1(_0148_),
    .B2(_0150_),
    .X(_0151_));
 sky130_fd_sc_hd__or3_1 _0695_ (.A(_0131_),
    .B(_0134_),
    .C(_0151_),
    .X(_0152_));
 sky130_fd_sc_hd__o211a_1 _0696_ (.A1(\frequency_counter_0.edge_counter[3] ),
    .A2(_0135_),
    .B1(_0152_),
    .C1(_0140_),
    .X(_0005_));
 sky130_fd_sc_hd__a22o_1 _0697_ (.A1(\frequency_counter_0.state[2] ),
    .A2(_0146_),
    .B1(_0132_),
    .B2(_0149_),
    .X(_0153_));
 sky130_fd_sc_hd__a21oi_1 _0698_ (.A1(_0135_),
    .A2(_0153_),
    .B1(\frequency_counter_0.edge_counter[4] ),
    .Y(_0154_));
 sky130_fd_sc_hd__a21oi_1 _0699_ (.A1(\frequency_counter_0.state[2] ),
    .A2(_0104_),
    .B1(_0150_),
    .Y(_0155_));
 sky130_fd_sc_hd__a31o_1 _0700_ (.A1(\frequency_counter_0.edge_counter[4] ),
    .A2(_0135_),
    .A3(_0155_),
    .B1(_0064_),
    .X(_0156_));
 sky130_fd_sc_hd__nor2_1 _0701_ (.A(_0154_),
    .B(_0156_),
    .Y(_0006_));
 sky130_fd_sc_hd__a21oi_1 _0702_ (.A1(\frequency_counter_0.edge_counter[4] ),
    .A2(_0149_),
    .B1(\frequency_counter_0.edge_counter[5] ),
    .Y(_0157_));
 sky130_fd_sc_hd__and3_1 _0703_ (.A(\frequency_counter_0.edge_counter[5] ),
    .B(\frequency_counter_0.edge_counter[4] ),
    .C(_0149_),
    .X(_0158_));
 sky130_fd_sc_hd__or2_1 _0704_ (.A(_0136_),
    .B(_0158_),
    .X(_0159_));
 sky130_fd_sc_hd__o21ai_1 _0705_ (.A1(\frequency_counter_0.edge_counter[4] ),
    .A2(_0104_),
    .B1(\frequency_counter_0.edge_counter[5] ),
    .Y(_0160_));
 sky130_fd_sc_hd__a21o_1 _0706_ (.A1(_0105_),
    .A2(_0160_),
    .B1(_0129_),
    .X(_0161_));
 sky130_fd_sc_hd__o211ai_1 _0707_ (.A1(_0157_),
    .A2(_0159_),
    .B1(_0161_),
    .C1(_0135_),
    .Y(_0162_));
 sky130_fd_sc_hd__o211a_1 _0708_ (.A1(\frequency_counter_0.edge_counter[5] ),
    .A2(_0135_),
    .B1(_0162_),
    .C1(_0140_),
    .X(_0007_));
 sky130_fd_sc_hd__a21oi_1 _0709_ (.A1(\frequency_counter_0.state[2] ),
    .A2(_0105_),
    .B1(_0134_),
    .Y(_0163_));
 sky130_fd_sc_hd__o211a_1 _0710_ (.A1(\frequency_counter_0.edge_counter[6] ),
    .A2(_0136_),
    .B1(_0159_),
    .C1(_0163_),
    .X(_0164_));
 sky130_fd_sc_hd__nor2_1 _0711_ (.A(_0136_),
    .B(_0134_),
    .Y(_0165_));
 sky130_fd_sc_hd__a21oi_1 _0712_ (.A1(_0158_),
    .A2(_0165_),
    .B1(\frequency_counter_0.edge_counter[6] ),
    .Y(_0166_));
 sky130_fd_sc_hd__nor3_1 _0713_ (.A(_0065_),
    .B(_0164_),
    .C(_0166_),
    .Y(_0008_));
 sky130_fd_sc_hd__mux2_1 _0714_ (.A0(\frequency_counter_0.seven_segment0.ten_count_reg[0] ),
    .A1(\frequency_counter_0.seven_segment0.ten_count[0] ),
    .S(\frequency_counter_0.seven_segment0.load ),
    .X(_0167_));
 sky130_fd_sc_hd__and2_1 _0715_ (.A(_0140_),
    .B(_0167_),
    .X(_0168_));
 sky130_fd_sc_hd__clkbuf_1 _0716_ (.A(_0168_),
    .X(_0009_));
 sky130_fd_sc_hd__buf_2 _0717_ (.A(_0139_),
    .X(_0169_));
 sky130_fd_sc_hd__mux2_1 _0718_ (.A0(\frequency_counter_0.seven_segment0.ten_count_reg[1] ),
    .A1(\frequency_counter_0.seven_segment0.ten_count[1] ),
    .S(\frequency_counter_0.seven_segment0.load ),
    .X(_0170_));
 sky130_fd_sc_hd__and2_1 _0719_ (.A(_0169_),
    .B(_0170_),
    .X(_0171_));
 sky130_fd_sc_hd__clkbuf_1 _0720_ (.A(_0171_),
    .X(_0010_));
 sky130_fd_sc_hd__mux2_1 _0721_ (.A0(\frequency_counter_0.seven_segment0.ten_count_reg[2] ),
    .A1(\frequency_counter_0.seven_segment0.ten_count[2] ),
    .S(\frequency_counter_0.seven_segment0.load ),
    .X(_0172_));
 sky130_fd_sc_hd__and2_1 _0722_ (.A(_0169_),
    .B(_0172_),
    .X(_0173_));
 sky130_fd_sc_hd__clkbuf_1 _0723_ (.A(_0173_),
    .X(_0011_));
 sky130_fd_sc_hd__mux2_1 _0724_ (.A0(\frequency_counter_0.seven_segment0.ten_count_reg[3] ),
    .A1(\frequency_counter_0.seven_segment0.ten_count[3] ),
    .S(\frequency_counter_0.seven_segment0.load ),
    .X(_0174_));
 sky130_fd_sc_hd__and2_1 _0725_ (.A(_0169_),
    .B(_0174_),
    .X(_0175_));
 sky130_fd_sc_hd__clkbuf_1 _0726_ (.A(_0175_),
    .X(_0012_));
 sky130_fd_sc_hd__mux2_1 _0727_ (.A0(\frequency_counter_0.seven_segment0.unit_count_reg[0] ),
    .A1(\frequency_counter_0.seven_segment0.unit_count[0] ),
    .S(\frequency_counter_0.seven_segment0.load ),
    .X(_0176_));
 sky130_fd_sc_hd__and2_1 _0728_ (.A(_0169_),
    .B(_0176_),
    .X(_0177_));
 sky130_fd_sc_hd__clkbuf_1 _0729_ (.A(_0177_),
    .X(_0013_));
 sky130_fd_sc_hd__mux2_1 _0730_ (.A0(\frequency_counter_0.seven_segment0.unit_count_reg[1] ),
    .A1(\frequency_counter_0.seven_segment0.unit_count[1] ),
    .S(\frequency_counter_0.seven_segment0.load ),
    .X(_0178_));
 sky130_fd_sc_hd__and2_1 _0731_ (.A(_0169_),
    .B(_0178_),
    .X(_0179_));
 sky130_fd_sc_hd__clkbuf_1 _0732_ (.A(_0179_),
    .X(_0014_));
 sky130_fd_sc_hd__mux2_1 _0733_ (.A0(\frequency_counter_0.seven_segment0.unit_count_reg[2] ),
    .A1(\frequency_counter_0.seven_segment0.unit_count[2] ),
    .S(\frequency_counter_0.seven_segment0.load ),
    .X(_0180_));
 sky130_fd_sc_hd__and2_1 _0734_ (.A(_0169_),
    .B(_0180_),
    .X(_0181_));
 sky130_fd_sc_hd__clkbuf_1 _0735_ (.A(_0181_),
    .X(_0015_));
 sky130_fd_sc_hd__mux2_1 _0736_ (.A0(\frequency_counter_0.seven_segment0.unit_count_reg[3] ),
    .A1(\frequency_counter_0.seven_segment0.unit_count[3] ),
    .S(\frequency_counter_0.seven_segment0.load ),
    .X(_0182_));
 sky130_fd_sc_hd__and2_1 _0737_ (.A(_0169_),
    .B(_0182_),
    .X(_0183_));
 sky130_fd_sc_hd__clkbuf_1 _0738_ (.A(_0183_),
    .X(_0016_));
 sky130_fd_sc_hd__buf_4 _0739_ (.A(net8),
    .X(_0184_));
 sky130_fd_sc_hd__mux2_1 _0740_ (.A0(\frequency_counter_0.update_period[0] ),
    .A1(net9),
    .S(_0184_),
    .X(_0185_));
 sky130_fd_sc_hd__or2_1 _0741_ (.A(_0065_),
    .B(_0185_),
    .X(_0186_));
 sky130_fd_sc_hd__clkbuf_1 _0742_ (.A(_0186_),
    .X(_0017_));
 sky130_fd_sc_hd__mux2_1 _0743_ (.A0(\frequency_counter_0.update_period[1] ),
    .A1(net10),
    .S(_0184_),
    .X(_0187_));
 sky130_fd_sc_hd__or2_1 _0744_ (.A(_0065_),
    .B(_0187_),
    .X(_0188_));
 sky130_fd_sc_hd__clkbuf_1 _0745_ (.A(_0188_),
    .X(_0018_));
 sky130_fd_sc_hd__mux2_1 _0746_ (.A0(\frequency_counter_0.update_period[2] ),
    .A1(net11),
    .S(_0184_),
    .X(_0189_));
 sky130_fd_sc_hd__or2_1 _0747_ (.A(_0065_),
    .B(_0189_),
    .X(_0190_));
 sky130_fd_sc_hd__clkbuf_1 _0748_ (.A(_0190_),
    .X(_0019_));
 sky130_fd_sc_hd__mux2_1 _0749_ (.A0(\frequency_counter_0.update_period[3] ),
    .A1(net12),
    .S(_0184_),
    .X(_0191_));
 sky130_fd_sc_hd__or2_1 _0750_ (.A(_0064_),
    .B(_0191_),
    .X(_0192_));
 sky130_fd_sc_hd__clkbuf_1 _0751_ (.A(_0192_),
    .X(_0020_));
 sky130_fd_sc_hd__mux2_1 _0752_ (.A0(\frequency_counter_0.update_period[4] ),
    .A1(net13),
    .S(_0184_),
    .X(_0193_));
 sky130_fd_sc_hd__and2_1 _0753_ (.A(_0169_),
    .B(_0193_),
    .X(_0194_));
 sky130_fd_sc_hd__clkbuf_1 _0754_ (.A(_0194_),
    .X(_0021_));
 sky130_fd_sc_hd__mux2_1 _0755_ (.A0(\frequency_counter_0.update_period[5] ),
    .A1(net14),
    .S(_0184_),
    .X(_0195_));
 sky130_fd_sc_hd__or2_1 _0756_ (.A(_0064_),
    .B(_0195_),
    .X(_0196_));
 sky130_fd_sc_hd__clkbuf_1 _0757_ (.A(_0196_),
    .X(_0022_));
 sky130_fd_sc_hd__mux2_1 _0758_ (.A0(\frequency_counter_0.update_period[6] ),
    .A1(net15),
    .S(_0184_),
    .X(_0197_));
 sky130_fd_sc_hd__and2_1 _0759_ (.A(_0169_),
    .B(_0197_),
    .X(_0198_));
 sky130_fd_sc_hd__clkbuf_1 _0760_ (.A(_0198_),
    .X(_0023_));
 sky130_fd_sc_hd__mux2_1 _0761_ (.A0(\frequency_counter_0.update_period[7] ),
    .A1(net16),
    .S(net8),
    .X(_0199_));
 sky130_fd_sc_hd__or2_1 _0762_ (.A(_0064_),
    .B(_0199_),
    .X(_0200_));
 sky130_fd_sc_hd__clkbuf_1 _0763_ (.A(_0200_),
    .X(_0024_));
 sky130_fd_sc_hd__mux2_1 _0764_ (.A0(\frequency_counter_0.update_period[8] ),
    .A1(net4),
    .S(_0184_),
    .X(_0201_));
 sky130_fd_sc_hd__and2_1 _0765_ (.A(_0169_),
    .B(_0201_),
    .X(_0202_));
 sky130_fd_sc_hd__clkbuf_1 _0766_ (.A(_0202_),
    .X(_0025_));
 sky130_fd_sc_hd__mux2_1 _0767_ (.A0(\frequency_counter_0.update_period[9] ),
    .A1(net5),
    .S(_0184_),
    .X(_0203_));
 sky130_fd_sc_hd__and2_1 _0768_ (.A(_0139_),
    .B(_0203_),
    .X(_0204_));
 sky130_fd_sc_hd__clkbuf_1 _0769_ (.A(_0204_),
    .X(_0026_));
 sky130_fd_sc_hd__mux2_1 _0770_ (.A0(\frequency_counter_0.update_period[10] ),
    .A1(net6),
    .S(net8),
    .X(_0205_));
 sky130_fd_sc_hd__or2_1 _0771_ (.A(_0064_),
    .B(_0205_),
    .X(_0206_));
 sky130_fd_sc_hd__clkbuf_1 _0772_ (.A(_0206_),
    .X(_0027_));
 sky130_fd_sc_hd__mux2_1 _0773_ (.A0(\frequency_counter_0.update_period[11] ),
    .A1(net7),
    .S(_0184_),
    .X(_0207_));
 sky130_fd_sc_hd__and2_1 _0774_ (.A(_0139_),
    .B(_0207_),
    .X(_0208_));
 sky130_fd_sc_hd__clkbuf_1 _0775_ (.A(_0208_),
    .X(_0028_));
 sky130_fd_sc_hd__a21oi_1 _0776_ (.A1(_0108_),
    .A2(\frequency_counter_0.seven_segment0.load ),
    .B1(\frequency_counter_0.state[1] ),
    .Y(_0209_));
 sky130_fd_sc_hd__nor2_1 _0777_ (.A(_0065_),
    .B(_0209_),
    .Y(_0029_));
 sky130_fd_sc_hd__or2_1 _0778_ (.A(_0066_),
    .B(\frequency_counter_0.state[1] ),
    .X(_0210_));
 sky130_fd_sc_hd__a21boi_1 _0779_ (.A1(_0110_),
    .A2(_0210_),
    .B1_N(\frequency_counter_0.seven_segment0.unit_count[0] ),
    .Y(_0211_));
 sky130_fd_sc_hd__and3_1 _0780_ (.A(\frequency_counter_0.edge_counter[0] ),
    .B(\frequency_counter_0.state[1] ),
    .C(_0110_),
    .X(_0212_));
 sky130_fd_sc_hd__o21a_1 _0781_ (.A1(_0211_),
    .A2(_0212_),
    .B1(_0140_),
    .X(_0030_));
 sky130_fd_sc_hd__a21boi_1 _0782_ (.A1(_0110_),
    .A2(_0210_),
    .B1_N(\frequency_counter_0.seven_segment0.unit_count[1] ),
    .Y(_0213_));
 sky130_fd_sc_hd__and3_1 _0783_ (.A(\frequency_counter_0.state[1] ),
    .B(_0103_),
    .C(_0110_),
    .X(_0214_));
 sky130_fd_sc_hd__o21a_1 _0784_ (.A1(_0213_),
    .A2(_0214_),
    .B1(_0140_),
    .X(_0031_));
 sky130_fd_sc_hd__a21boi_1 _0785_ (.A1(_0110_),
    .A2(_0210_),
    .B1_N(\frequency_counter_0.seven_segment0.unit_count[2] ),
    .Y(_0215_));
 sky130_fd_sc_hd__and3_1 _0786_ (.A(\frequency_counter_0.state[1] ),
    .B(\frequency_counter_0.edge_counter[2] ),
    .C(_0110_),
    .X(_0216_));
 sky130_fd_sc_hd__o21a_1 _0787_ (.A1(_0215_),
    .A2(_0216_),
    .B1(_0140_),
    .X(_0032_));
 sky130_fd_sc_hd__a21boi_1 _0788_ (.A1(_0110_),
    .A2(_0210_),
    .B1_N(\frequency_counter_0.seven_segment0.unit_count[3] ),
    .Y(_0217_));
 sky130_fd_sc_hd__and3_1 _0789_ (.A(\frequency_counter_0.state[1] ),
    .B(\frequency_counter_0.edge_counter[3] ),
    .C(_0109_),
    .X(_0218_));
 sky130_fd_sc_hd__o21a_1 _0790_ (.A1(_0217_),
    .A2(_0218_),
    .B1(_0140_),
    .X(_0033_));
 sky130_fd_sc_hd__a21oi_1 _0791_ (.A1(_0106_),
    .A2(_0110_),
    .B1(\frequency_counter_0.seven_segment0.ten_count[0] ),
    .Y(_0219_));
 sky130_fd_sc_hd__o21a_1 _0792_ (.A1(_0066_),
    .A2(\frequency_counter_0.state[2] ),
    .B1(_0130_),
    .X(_0220_));
 sky130_fd_sc_hd__and3_1 _0793_ (.A(\frequency_counter_0.seven_segment0.ten_count[0] ),
    .B(_0109_),
    .C(_0220_),
    .X(_0221_));
 sky130_fd_sc_hd__nor3_1 _0794_ (.A(_0065_),
    .B(_0219_),
    .C(_0221_),
    .Y(_0034_));
 sky130_fd_sc_hd__a21o_1 _0795_ (.A1(\frequency_counter_0.seven_segment0.ten_count[1] ),
    .A2(\frequency_counter_0.seven_segment0.ten_count[0] ),
    .B1(_0129_),
    .X(_0222_));
 sky130_fd_sc_hd__a31o_1 _0796_ (.A1(_0110_),
    .A2(_0220_),
    .A3(_0222_),
    .B1(_0064_),
    .X(_0223_));
 sky130_fd_sc_hd__o21ba_1 _0797_ (.A1(\frequency_counter_0.seven_segment0.ten_count[1] ),
    .A2(_0221_),
    .B1_N(_0223_),
    .X(_0035_));
 sky130_fd_sc_hd__and3_1 _0798_ (.A(\frequency_counter_0.seven_segment0.ten_count[2] ),
    .B(\frequency_counter_0.seven_segment0.ten_count[1] ),
    .C(\frequency_counter_0.seven_segment0.ten_count[0] ),
    .X(_0224_));
 sky130_fd_sc_hd__or2_1 _0799_ (.A(_0129_),
    .B(_0224_),
    .X(_0225_));
 sky130_fd_sc_hd__a31o_1 _0800_ (.A1(_0109_),
    .A2(_0220_),
    .A3(_0225_),
    .B1(_0064_),
    .X(_0226_));
 sky130_fd_sc_hd__a41o_1 _0801_ (.A1(\frequency_counter_0.seven_segment0.ten_count[1] ),
    .A2(\frequency_counter_0.seven_segment0.ten_count[0] ),
    .A3(_0109_),
    .A4(_0220_),
    .B1(\frequency_counter_0.seven_segment0.ten_count[2] ),
    .X(_0227_));
 sky130_fd_sc_hd__and2b_1 _0802_ (.A_N(_0226_),
    .B(_0227_),
    .X(_0228_));
 sky130_fd_sc_hd__clkbuf_1 _0803_ (.A(_0228_),
    .X(_0036_));
 sky130_fd_sc_hd__nand4_1 _0804_ (.A(\frequency_counter_0.seven_segment0.ten_count[3] ),
    .B(_0109_),
    .C(_0220_),
    .D(_0225_),
    .Y(_0229_));
 sky130_fd_sc_hd__a31o_1 _0805_ (.A1(_0106_),
    .A2(_0109_),
    .A3(_0224_),
    .B1(\frequency_counter_0.seven_segment0.ten_count[3] ),
    .X(_0230_));
 sky130_fd_sc_hd__and3_1 _0806_ (.A(_0139_),
    .B(_0229_),
    .C(_0230_),
    .X(_0231_));
 sky130_fd_sc_hd__clkbuf_1 _0807_ (.A(_0231_),
    .X(_0037_));
 sky130_fd_sc_hd__mux2_1 _0808_ (.A0(_0109_),
    .A1(_0066_),
    .S(\frequency_counter_0.clk_counter[0] ),
    .X(_0232_));
 sky130_fd_sc_hd__nor2_1 _0809_ (.A(_0065_),
    .B(_0232_),
    .Y(_0038_));
 sky130_fd_sc_hd__and3_1 _0810_ (.A(_0066_),
    .B(\frequency_counter_0.clk_counter[1] ),
    .C(\frequency_counter_0.clk_counter[0] ),
    .X(_0233_));
 sky130_fd_sc_hd__a21oi_1 _0811_ (.A1(_0066_),
    .A2(_0102_),
    .B1(_0064_),
    .Y(_0234_));
 sky130_fd_sc_hd__buf_2 _0812_ (.A(_0234_),
    .X(_0235_));
 sky130_fd_sc_hd__a21o_1 _0813_ (.A1(_0066_),
    .A2(\frequency_counter_0.clk_counter[0] ),
    .B1(\frequency_counter_0.clk_counter[1] ),
    .X(_0236_));
 sky130_fd_sc_hd__and3b_1 _0814_ (.A_N(_0233_),
    .B(_0235_),
    .C(_0236_),
    .X(_0237_));
 sky130_fd_sc_hd__clkbuf_1 _0815_ (.A(_0237_),
    .X(_0039_));
 sky130_fd_sc_hd__or2_1 _0816_ (.A(\frequency_counter_0.clk_counter[2] ),
    .B(_0233_),
    .X(_0238_));
 sky130_fd_sc_hd__nand2_1 _0817_ (.A(\frequency_counter_0.clk_counter[2] ),
    .B(_0233_),
    .Y(_0239_));
 sky130_fd_sc_hd__and3_1 _0818_ (.A(_0235_),
    .B(_0238_),
    .C(_0239_),
    .X(_0240_));
 sky130_fd_sc_hd__clkbuf_1 _0819_ (.A(_0240_),
    .X(_0040_));
 sky130_fd_sc_hd__and4_1 _0820_ (.A(\frequency_counter_0.clk_counter[3] ),
    .B(\frequency_counter_0.clk_counter[2] ),
    .C(\frequency_counter_0.clk_counter[1] ),
    .D(\frequency_counter_0.clk_counter[0] ),
    .X(_0241_));
 sky130_fd_sc_hd__nand2_1 _0821_ (.A(_0066_),
    .B(_0241_),
    .Y(_0242_));
 sky130_fd_sc_hd__a21o_1 _0822_ (.A1(\frequency_counter_0.clk_counter[2] ),
    .A2(_0233_),
    .B1(\frequency_counter_0.clk_counter[3] ),
    .X(_0243_));
 sky130_fd_sc_hd__and3_1 _0823_ (.A(_0235_),
    .B(_0242_),
    .C(_0243_),
    .X(_0244_));
 sky130_fd_sc_hd__clkbuf_1 _0824_ (.A(_0244_),
    .X(_0041_));
 sky130_fd_sc_hd__nand2_1 _0825_ (.A(_0080_),
    .B(_0242_),
    .Y(_0245_));
 sky130_fd_sc_hd__or3b_1 _0826_ (.A(_0108_),
    .B(_0080_),
    .C_N(_0241_),
    .X(_0246_));
 sky130_fd_sc_hd__and3_1 _0827_ (.A(_0235_),
    .B(_0245_),
    .C(_0246_),
    .X(_0247_));
 sky130_fd_sc_hd__clkbuf_1 _0828_ (.A(_0247_),
    .X(_0042_));
 sky130_fd_sc_hd__or2_1 _0829_ (.A(_0068_),
    .B(_0246_),
    .X(_0248_));
 sky130_fd_sc_hd__nand2_1 _0830_ (.A(_0068_),
    .B(_0246_),
    .Y(_0249_));
 sky130_fd_sc_hd__and3_1 _0831_ (.A(_0235_),
    .B(_0248_),
    .C(_0249_),
    .X(_0250_));
 sky130_fd_sc_hd__clkbuf_1 _0832_ (.A(_0250_),
    .X(_0043_));
 sky130_fd_sc_hd__or3_1 _0833_ (.A(_0067_),
    .B(_0068_),
    .C(_0246_),
    .X(_0251_));
 sky130_fd_sc_hd__nand2_1 _0834_ (.A(_0067_),
    .B(_0248_),
    .Y(_0252_));
 sky130_fd_sc_hd__and3_1 _0835_ (.A(_0235_),
    .B(_0251_),
    .C(_0252_),
    .X(_0253_));
 sky130_fd_sc_hd__clkbuf_1 _0836_ (.A(_0253_),
    .X(_0044_));
 sky130_fd_sc_hd__nor2_1 _0837_ (.A(_0078_),
    .B(_0251_),
    .Y(_0254_));
 sky130_fd_sc_hd__nand2_1 _0838_ (.A(_0078_),
    .B(_0251_),
    .Y(_0255_));
 sky130_fd_sc_hd__and3b_1 _0839_ (.A_N(_0254_),
    .B(_0235_),
    .C(_0255_),
    .X(_0256_));
 sky130_fd_sc_hd__clkbuf_1 _0840_ (.A(_0256_),
    .X(_0045_));
 sky130_fd_sc_hd__and2_1 _0841_ (.A(\frequency_counter_0.clk_counter[8] ),
    .B(_0254_),
    .X(_0257_));
 sky130_fd_sc_hd__or2_1 _0842_ (.A(\frequency_counter_0.clk_counter[8] ),
    .B(_0254_),
    .X(_0258_));
 sky130_fd_sc_hd__and3b_1 _0843_ (.A_N(_0257_),
    .B(_0235_),
    .C(_0258_),
    .X(_0259_));
 sky130_fd_sc_hd__clkbuf_1 _0844_ (.A(_0259_),
    .X(_0046_));
 sky130_fd_sc_hd__and3_1 _0845_ (.A(\frequency_counter_0.clk_counter[9] ),
    .B(\frequency_counter_0.clk_counter[8] ),
    .C(_0254_),
    .X(_0260_));
 sky130_fd_sc_hd__or2_1 _0846_ (.A(\frequency_counter_0.clk_counter[9] ),
    .B(_0257_),
    .X(_0261_));
 sky130_fd_sc_hd__and3b_1 _0847_ (.A_N(_0260_),
    .B(_0234_),
    .C(_0261_),
    .X(_0262_));
 sky130_fd_sc_hd__clkbuf_1 _0848_ (.A(_0262_),
    .X(_0047_));
 sky130_fd_sc_hd__or2_1 _0849_ (.A(\frequency_counter_0.clk_counter[10] ),
    .B(_0260_),
    .X(_0263_));
 sky130_fd_sc_hd__nand2_1 _0850_ (.A(\frequency_counter_0.clk_counter[10] ),
    .B(_0260_),
    .Y(_0264_));
 sky130_fd_sc_hd__and3_1 _0851_ (.A(_0235_),
    .B(_0263_),
    .C(_0264_),
    .X(_0265_));
 sky130_fd_sc_hd__clkbuf_1 _0852_ (.A(_0265_),
    .X(_0048_));
 sky130_fd_sc_hd__a21boi_1 _0853_ (.A1(_0096_),
    .A2(_0264_),
    .B1_N(_0235_),
    .Y(_0049_));
 sky130_fd_sc_hd__or3b_1 _0854_ (.A(\frequency_counter_0.state[2] ),
    .B(_0134_),
    .C_N(\frequency_counter_0.edge_counter[0] ),
    .X(_0266_));
 sky130_fd_sc_hd__o211a_1 _0855_ (.A1(\frequency_counter_0.edge_counter[0] ),
    .A2(_0165_),
    .B1(_0266_),
    .C1(_0140_),
    .X(_0050_));
 sky130_fd_sc_hd__nor2_1 _0856_ (.A(_0065_),
    .B(\frequency_counter_0.digit ),
    .Y(_0051_));
 sky130_fd_sc_hd__dfxtp_1 _0857_ (.CLK(clknet_2_3__leaf_wb_clk_i),
    .D(_0001_),
    .Q(\frequency_counter_0.state[0] ));
 sky130_fd_sc_hd__dfxtp_2 _0858_ (.CLK(clknet_2_3__leaf_wb_clk_i),
    .D(_0000_),
    .Q(\frequency_counter_0.state[1] ));
 sky130_fd_sc_hd__dfxtp_2 _0859_ (.CLK(clknet_2_3__leaf_wb_clk_i),
    .D(_0002_),
    .Q(\frequency_counter_0.state[2] ));
 sky130_fd_sc_hd__dfxtp_1 _0860_ (.CLK(clknet_2_1__leaf_wb_clk_i),
    .D(_0003_),
    .Q(\frequency_counter_0.edge_counter[1] ));
 sky130_fd_sc_hd__dfxtp_2 _0861_ (.CLK(clknet_2_1__leaf_wb_clk_i),
    .D(_0004_),
    .Q(\frequency_counter_0.edge_counter[2] ));
 sky130_fd_sc_hd__dfxtp_1 _0862_ (.CLK(clknet_2_1__leaf_wb_clk_i),
    .D(_0005_),
    .Q(\frequency_counter_0.edge_counter[3] ));
 sky130_fd_sc_hd__dfxtp_1 _0863_ (.CLK(clknet_2_3__leaf_wb_clk_i),
    .D(_0006_),
    .Q(\frequency_counter_0.edge_counter[4] ));
 sky130_fd_sc_hd__dfxtp_1 _0864_ (.CLK(clknet_2_3__leaf_wb_clk_i),
    .D(_0007_),
    .Q(\frequency_counter_0.edge_counter[5] ));
 sky130_fd_sc_hd__dfxtp_1 _0865_ (.CLK(clknet_2_3__leaf_wb_clk_i),
    .D(_0008_),
    .Q(\frequency_counter_0.edge_counter[6] ));
 sky130_fd_sc_hd__dfxtp_1 _0866_ (.CLK(clknet_2_0__leaf_wb_clk_i),
    .D(_0009_),
    .Q(\frequency_counter_0.seven_segment0.ten_count_reg[0] ));
 sky130_fd_sc_hd__dfxtp_1 _0867_ (.CLK(clknet_2_0__leaf_wb_clk_i),
    .D(_0010_),
    .Q(\frequency_counter_0.seven_segment0.ten_count_reg[1] ));
 sky130_fd_sc_hd__dfxtp_1 _0868_ (.CLK(clknet_2_0__leaf_wb_clk_i),
    .D(_0011_),
    .Q(\frequency_counter_0.seven_segment0.ten_count_reg[2] ));
 sky130_fd_sc_hd__dfxtp_1 _0869_ (.CLK(clknet_2_0__leaf_wb_clk_i),
    .D(_0012_),
    .Q(\frequency_counter_0.seven_segment0.ten_count_reg[3] ));
 sky130_fd_sc_hd__dfxtp_1 _0870_ (.CLK(clknet_2_0__leaf_wb_clk_i),
    .D(_0013_),
    .Q(\frequency_counter_0.seven_segment0.unit_count_reg[0] ));
 sky130_fd_sc_hd__dfxtp_1 _0871_ (.CLK(clknet_2_2__leaf_wb_clk_i),
    .D(_0014_),
    .Q(\frequency_counter_0.seven_segment0.unit_count_reg[1] ));
 sky130_fd_sc_hd__dfxtp_1 _0872_ (.CLK(clknet_2_0__leaf_wb_clk_i),
    .D(_0015_),
    .Q(\frequency_counter_0.seven_segment0.unit_count_reg[2] ));
 sky130_fd_sc_hd__dfxtp_1 _0873_ (.CLK(clknet_2_0__leaf_wb_clk_i),
    .D(_0016_),
    .Q(\frequency_counter_0.seven_segment0.unit_count_reg[3] ));
 sky130_fd_sc_hd__dfxtp_1 _0874_ (.CLK(clknet_2_3__leaf_wb_clk_i),
    .D(net2),
    .Q(\frequency_counter_0.edge_detect0.q0 ));
 sky130_fd_sc_hd__dfxtp_1 _0875_ (.CLK(clknet_2_3__leaf_wb_clk_i),
    .D(net117),
    .Q(\frequency_counter_0.edge_detect0.q1 ));
 sky130_fd_sc_hd__dfxtp_1 _0876_ (.CLK(clknet_2_3__leaf_wb_clk_i),
    .D(net118),
    .Q(\frequency_counter_0.edge_detect0.q2 ));
 sky130_fd_sc_hd__dfxtp_1 _0877_ (.CLK(clknet_2_0__leaf_wb_clk_i),
    .D(_0017_),
    .Q(\frequency_counter_0.update_period[0] ));
 sky130_fd_sc_hd__dfxtp_1 _0878_ (.CLK(clknet_2_2__leaf_wb_clk_i),
    .D(_0018_),
    .Q(\frequency_counter_0.update_period[1] ));
 sky130_fd_sc_hd__dfxtp_1 _0879_ (.CLK(clknet_2_3__leaf_wb_clk_i),
    .D(_0019_),
    .Q(\frequency_counter_0.update_period[2] ));
 sky130_fd_sc_hd__dfxtp_1 _0880_ (.CLK(clknet_2_3__leaf_wb_clk_i),
    .D(_0020_),
    .Q(\frequency_counter_0.update_period[3] ));
 sky130_fd_sc_hd__dfxtp_1 _0881_ (.CLK(clknet_2_2__leaf_wb_clk_i),
    .D(_0021_),
    .Q(\frequency_counter_0.update_period[4] ));
 sky130_fd_sc_hd__dfxtp_1 _0882_ (.CLK(clknet_2_0__leaf_wb_clk_i),
    .D(_0022_),
    .Q(\frequency_counter_0.update_period[5] ));
 sky130_fd_sc_hd__dfxtp_1 _0883_ (.CLK(clknet_2_2__leaf_wb_clk_i),
    .D(_0023_),
    .Q(\frequency_counter_0.update_period[6] ));
 sky130_fd_sc_hd__dfxtp_1 _0884_ (.CLK(clknet_2_2__leaf_wb_clk_i),
    .D(_0024_),
    .Q(\frequency_counter_0.update_period[7] ));
 sky130_fd_sc_hd__dfxtp_1 _0885_ (.CLK(clknet_2_0__leaf_wb_clk_i),
    .D(_0025_),
    .Q(\frequency_counter_0.update_period[8] ));
 sky130_fd_sc_hd__dfxtp_1 _0886_ (.CLK(clknet_2_1__leaf_wb_clk_i),
    .D(_0026_),
    .Q(\frequency_counter_0.update_period[9] ));
 sky130_fd_sc_hd__dfxtp_1 _0887_ (.CLK(clknet_2_0__leaf_wb_clk_i),
    .D(_0027_),
    .Q(\frequency_counter_0.update_period[10] ));
 sky130_fd_sc_hd__dfxtp_1 _0888_ (.CLK(clknet_2_1__leaf_wb_clk_i),
    .D(_0028_),
    .Q(\frequency_counter_0.update_period[11] ));
 sky130_fd_sc_hd__dfxtp_4 _0889_ (.CLK(clknet_2_2__leaf_wb_clk_i),
    .D(_0029_),
    .Q(\frequency_counter_0.seven_segment0.load ));
 sky130_fd_sc_hd__dfxtp_1 _0890_ (.CLK(clknet_2_1__leaf_wb_clk_i),
    .D(_0030_),
    .Q(\frequency_counter_0.seven_segment0.unit_count[0] ));
 sky130_fd_sc_hd__dfxtp_1 _0891_ (.CLK(clknet_2_2__leaf_wb_clk_i),
    .D(_0031_),
    .Q(\frequency_counter_0.seven_segment0.unit_count[1] ));
 sky130_fd_sc_hd__dfxtp_1 _0892_ (.CLK(clknet_2_1__leaf_wb_clk_i),
    .D(_0032_),
    .Q(\frequency_counter_0.seven_segment0.unit_count[2] ));
 sky130_fd_sc_hd__dfxtp_1 _0893_ (.CLK(clknet_2_0__leaf_wb_clk_i),
    .D(_0033_),
    .Q(\frequency_counter_0.seven_segment0.unit_count[3] ));
 sky130_fd_sc_hd__dfxtp_1 _0894_ (.CLK(clknet_2_1__leaf_wb_clk_i),
    .D(_0034_),
    .Q(\frequency_counter_0.seven_segment0.ten_count[0] ));
 sky130_fd_sc_hd__dfxtp_1 _0895_ (.CLK(clknet_2_1__leaf_wb_clk_i),
    .D(_0035_),
    .Q(\frequency_counter_0.seven_segment0.ten_count[1] ));
 sky130_fd_sc_hd__dfxtp_1 _0896_ (.CLK(clknet_2_1__leaf_wb_clk_i),
    .D(_0036_),
    .Q(\frequency_counter_0.seven_segment0.ten_count[2] ));
 sky130_fd_sc_hd__dfxtp_1 _0897_ (.CLK(clknet_2_1__leaf_wb_clk_i),
    .D(_0037_),
    .Q(\frequency_counter_0.seven_segment0.ten_count[3] ));
 sky130_fd_sc_hd__dfxtp_1 _0898_ (.CLK(clknet_2_2__leaf_wb_clk_i),
    .D(_0038_),
    .Q(\frequency_counter_0.clk_counter[0] ));
 sky130_fd_sc_hd__dfxtp_1 _0899_ (.CLK(clknet_2_2__leaf_wb_clk_i),
    .D(_0039_),
    .Q(\frequency_counter_0.clk_counter[1] ));
 sky130_fd_sc_hd__dfxtp_1 _0900_ (.CLK(clknet_2_3__leaf_wb_clk_i),
    .D(_0040_),
    .Q(\frequency_counter_0.clk_counter[2] ));
 sky130_fd_sc_hd__dfxtp_1 _0901_ (.CLK(clknet_2_2__leaf_wb_clk_i),
    .D(_0041_),
    .Q(\frequency_counter_0.clk_counter[3] ));
 sky130_fd_sc_hd__dfxtp_1 _0902_ (.CLK(clknet_2_2__leaf_wb_clk_i),
    .D(_0042_),
    .Q(\frequency_counter_0.clk_counter[4] ));
 sky130_fd_sc_hd__dfxtp_1 _0903_ (.CLK(clknet_2_2__leaf_wb_clk_i),
    .D(_0043_),
    .Q(\frequency_counter_0.clk_counter[5] ));
 sky130_fd_sc_hd__dfxtp_1 _0904_ (.CLK(clknet_2_2__leaf_wb_clk_i),
    .D(_0044_),
    .Q(\frequency_counter_0.clk_counter[6] ));
 sky130_fd_sc_hd__dfxtp_1 _0905_ (.CLK(clknet_2_2__leaf_wb_clk_i),
    .D(_0045_),
    .Q(\frequency_counter_0.clk_counter[7] ));
 sky130_fd_sc_hd__dfxtp_1 _0906_ (.CLK(clknet_2_0__leaf_wb_clk_i),
    .D(_0046_),
    .Q(\frequency_counter_0.clk_counter[8] ));
 sky130_fd_sc_hd__dfxtp_1 _0907_ (.CLK(clknet_2_0__leaf_wb_clk_i),
    .D(_0047_),
    .Q(\frequency_counter_0.clk_counter[9] ));
 sky130_fd_sc_hd__dfxtp_1 _0908_ (.CLK(clknet_2_0__leaf_wb_clk_i),
    .D(_0048_),
    .Q(\frequency_counter_0.clk_counter[10] ));
 sky130_fd_sc_hd__dfxtp_1 _0909_ (.CLK(clknet_2_0__leaf_wb_clk_i),
    .D(_0049_),
    .Q(\frequency_counter_0.clk_counter[11] ));
 sky130_fd_sc_hd__dfxtp_1 _0910_ (.CLK(clknet_2_1__leaf_wb_clk_i),
    .D(_0050_),
    .Q(\frequency_counter_0.edge_counter[0] ));
 sky130_fd_sc_hd__dfxtp_2 _0911_ (.CLK(clknet_2_3__leaf_wb_clk_i),
    .D(_0051_),
    .Q(\frequency_counter_0.digit ));
 sky130_fd_sc_hd__conb_1 _1013__18 (.LO(net18));
 sky130_fd_sc_hd__conb_1 _1014__19 (.LO(net19));
 sky130_fd_sc_hd__conb_1 _1015__20 (.LO(net20));
 sky130_fd_sc_hd__conb_1 _1016__21 (.LO(net21));
 sky130_fd_sc_hd__conb_1 _1017__22 (.LO(net22));
 sky130_fd_sc_hd__conb_1 _1018__23 (.LO(net23));
 sky130_fd_sc_hd__conb_1 _1019__24 (.LO(net24));
 sky130_fd_sc_hd__conb_1 _1020__25 (.LO(net25));
 sky130_fd_sc_hd__conb_1 _1021__26 (.LO(net26));
 sky130_fd_sc_hd__conb_1 _1022__27 (.LO(net27));
 sky130_fd_sc_hd__conb_1 _1023__28 (.LO(net28));
 sky130_fd_sc_hd__conb_1 _1024__29 (.LO(net29));
 sky130_fd_sc_hd__conb_1 _1025__30 (.LO(net30));
 sky130_fd_sc_hd__conb_1 _1026__31 (.LO(net31));
 sky130_fd_sc_hd__conb_1 _1027__32 (.LO(net32));
 sky130_fd_sc_hd__conb_1 _1028__33 (.LO(net33));
 sky130_fd_sc_hd__conb_1 _1029__34 (.LO(net34));
 sky130_fd_sc_hd__conb_1 _1030__35 (.LO(net35));
 sky130_fd_sc_hd__conb_1 _1031__36 (.LO(net36));
 sky130_fd_sc_hd__conb_1 _1032__37 (.LO(net37));
 sky130_fd_sc_hd__conb_1 _1033__38 (.LO(net38));
 sky130_fd_sc_hd__conb_1 _1034__39 (.LO(net39));
 sky130_fd_sc_hd__conb_1 _1035__40 (.LO(net40));
 sky130_fd_sc_hd__conb_1 _1036__41 (.LO(net41));
 sky130_fd_sc_hd__conb_1 _1037__42 (.LO(net42));
 sky130_fd_sc_hd__conb_1 _1038__43 (.LO(net43));
 sky130_fd_sc_hd__conb_1 _1039__44 (.LO(net44));
 sky130_fd_sc_hd__conb_1 _1040__45 (.LO(net45));
 sky130_fd_sc_hd__conb_1 _1041__46 (.LO(net46));
 sky130_fd_sc_hd__conb_1 _1042__47 (.LO(net47));
 sky130_fd_sc_hd__conb_1 _1043__48 (.LO(net48));
 sky130_fd_sc_hd__conb_1 _1044__49 (.LO(net49));
 sky130_fd_sc_hd__conb_1 _1045__50 (.LO(net50));
 sky130_fd_sc_hd__conb_1 _1046__51 (.LO(net51));
 sky130_fd_sc_hd__conb_1 _1047__52 (.LO(net52));
 sky130_fd_sc_hd__conb_1 _1048__53 (.LO(net53));
 sky130_fd_sc_hd__conb_1 _1049__54 (.LO(net54));
 sky130_fd_sc_hd__conb_1 _1050__55 (.LO(net55));
 sky130_fd_sc_hd__conb_1 _1051__56 (.LO(net56));
 sky130_fd_sc_hd__conb_1 _1052__57 (.LO(net57));
 sky130_fd_sc_hd__conb_1 _1061__58 (.LO(net58));
 sky130_fd_sc_hd__conb_1 _1062__59 (.LO(net59));
 sky130_fd_sc_hd__conb_1 _1063__60 (.LO(net60));
 sky130_fd_sc_hd__conb_1 _1064__61 (.LO(net61));
 sky130_fd_sc_hd__conb_1 _1065__62 (.LO(net62));
 sky130_fd_sc_hd__conb_1 _1066__63 (.LO(net63));
 sky130_fd_sc_hd__conb_1 _1067__64 (.LO(net64));
 sky130_fd_sc_hd__conb_1 _1068__65 (.LO(net65));
 sky130_fd_sc_hd__conb_1 _1069__66 (.LO(net66));
 sky130_fd_sc_hd__conb_1 _1070__67 (.LO(net67));
 sky130_fd_sc_hd__conb_1 _1071__68 (.LO(net68));
 sky130_fd_sc_hd__conb_1 _1072__69 (.LO(net69));
 sky130_fd_sc_hd__conb_1 _1073__70 (.LO(net70));
 sky130_fd_sc_hd__conb_1 _1074__71 (.LO(net71));
 sky130_fd_sc_hd__conb_1 _1075__72 (.LO(net72));
 sky130_fd_sc_hd__conb_1 _1076__73 (.LO(net73));
 sky130_fd_sc_hd__conb_1 _1077__74 (.LO(net74));
 sky130_fd_sc_hd__conb_1 _1078__75 (.LO(net75));
 sky130_fd_sc_hd__conb_1 _1079__76 (.LO(net76));
 sky130_fd_sc_hd__conb_1 _1080__77 (.LO(net77));
 sky130_fd_sc_hd__conb_1 _1081__78 (.LO(net78));
 sky130_fd_sc_hd__conb_1 _1082__79 (.LO(net79));
 sky130_fd_sc_hd__conb_1 _1083__80 (.LO(net80));
 sky130_fd_sc_hd__conb_1 _1084__81 (.LO(net81));
 sky130_fd_sc_hd__conb_1 _1085__82 (.LO(net82));
 sky130_fd_sc_hd__conb_1 _1086__83 (.LO(net83));
 sky130_fd_sc_hd__conb_1 _1087__84 (.LO(net84));
 sky130_fd_sc_hd__conb_1 _1088__85 (.LO(net85));
 sky130_fd_sc_hd__conb_1 _1089__86 (.LO(net86));
 sky130_fd_sc_hd__conb_1 _1090__87 (.LO(net87));
 sky130_fd_sc_hd__conb_1 _1091__88 (.LO(net88));
 sky130_fd_sc_hd__conb_1 _1092__89 (.LO(net89));
 sky130_fd_sc_hd__conb_1 _1093__90 (.LO(net90));
 sky130_fd_sc_hd__conb_1 _1094__91 (.LO(net91));
 sky130_fd_sc_hd__conb_1 _1095__92 (.LO(net92));
 sky130_fd_sc_hd__conb_1 _1096__93 (.LO(net93));
 sky130_fd_sc_hd__conb_1 _1097__94 (.LO(net94));
 sky130_fd_sc_hd__conb_1 _1098__95 (.LO(net95));
 sky130_fd_sc_hd__conb_1 _1099__96 (.LO(net96));
 sky130_fd_sc_hd__conb_1 _1100__97 (.LO(net97));
 sky130_fd_sc_hd__conb_1 _1101__98 (.LO(net98));
 sky130_fd_sc_hd__conb_1 _1102__99 (.LO(net99));
 sky130_fd_sc_hd__conb_1 _1103__100 (.LO(net100));
 sky130_fd_sc_hd__conb_1 _1104__101 (.LO(net101));
 sky130_fd_sc_hd__conb_1 _1105__102 (.LO(net102));
 sky130_fd_sc_hd__conb_1 _1106__103 (.LO(net103));
 sky130_fd_sc_hd__conb_1 _1107__104 (.LO(net104));
 sky130_fd_sc_hd__conb_1 _1108__105 (.LO(net105));
 sky130_fd_sc_hd__conb_1 _1109__106 (.LO(net106));
 sky130_fd_sc_hd__conb_1 _1110__107 (.LO(net107));
 sky130_fd_sc_hd__conb_1 _1111__108 (.LO(net108));
 sky130_fd_sc_hd__conb_1 _1112__109 (.LO(net109));
 sky130_fd_sc_hd__conb_1 _1113__110 (.LO(net110));
 sky130_fd_sc_hd__conb_1 _1114__111 (.LO(net111));
 sky130_fd_sc_hd__conb_1 _1115__112 (.LO(net112));
 sky130_fd_sc_hd__conb_1 _1116__113 (.LO(net113));
 sky130_fd_sc_hd__conb_1 _1117__114 (.LO(net114));
 sky130_fd_sc_hd__conb_1 _1118__115 (.LO(net115));
 sky130_fd_sc_hd__conb_1 _1119__116 (.LO(net116));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_wb_clk_i (.A(wb_clk_i),
    .X(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__ebufn_8 _1012_ (.A(net17),
    .TE_B(_0267_),
    .Z(la1_data_out[0]));
 sky130_fd_sc_hd__ebufn_8 _1013_ (.A(net18),
    .TE_B(_0268_),
    .Z(la1_data_out[1]));
 sky130_fd_sc_hd__ebufn_8 _1014_ (.A(net19),
    .TE_B(_0269_),
    .Z(la1_data_out[2]));
 sky130_fd_sc_hd__ebufn_8 _1015_ (.A(net20),
    .TE_B(_0270_),
    .Z(la1_data_out[3]));
 sky130_fd_sc_hd__ebufn_8 _1016_ (.A(net21),
    .TE_B(_0271_),
    .Z(la1_data_out[4]));
 sky130_fd_sc_hd__ebufn_8 _1017_ (.A(net22),
    .TE_B(_0272_),
    .Z(la1_data_out[5]));
 sky130_fd_sc_hd__ebufn_8 _1018_ (.A(net23),
    .TE_B(_0273_),
    .Z(la1_data_out[6]));
 sky130_fd_sc_hd__ebufn_8 _1019_ (.A(net24),
    .TE_B(_0274_),
    .Z(la1_data_out[7]));
 sky130_fd_sc_hd__ebufn_8 _1020_ (.A(net25),
    .TE_B(_0275_),
    .Z(la1_data_out[8]));
 sky130_fd_sc_hd__ebufn_8 _1021_ (.A(net26),
    .TE_B(_0276_),
    .Z(la1_data_out[9]));
 sky130_fd_sc_hd__ebufn_8 _1022_ (.A(net27),
    .TE_B(_0277_),
    .Z(la1_data_out[10]));
 sky130_fd_sc_hd__ebufn_8 _1023_ (.A(net28),
    .TE_B(_0278_),
    .Z(la1_data_out[11]));
 sky130_fd_sc_hd__ebufn_8 _1024_ (.A(net29),
    .TE_B(_0279_),
    .Z(la1_data_out[12]));
 sky130_fd_sc_hd__ebufn_8 _1025_ (.A(net30),
    .TE_B(_0280_),
    .Z(la1_data_out[13]));
 sky130_fd_sc_hd__ebufn_8 _1026_ (.A(net31),
    .TE_B(_0281_),
    .Z(la1_data_out[14]));
 sky130_fd_sc_hd__ebufn_8 _1027_ (.A(net32),
    .TE_B(_0282_),
    .Z(la1_data_out[15]));
 sky130_fd_sc_hd__ebufn_8 _1028_ (.A(net33),
    .TE_B(_0283_),
    .Z(la1_data_out[16]));
 sky130_fd_sc_hd__ebufn_8 _1029_ (.A(net34),
    .TE_B(_0284_),
    .Z(la1_data_out[17]));
 sky130_fd_sc_hd__ebufn_8 _1030_ (.A(net35),
    .TE_B(_0285_),
    .Z(la1_data_out[18]));
 sky130_fd_sc_hd__ebufn_8 _1031_ (.A(net36),
    .TE_B(_0286_),
    .Z(la1_data_out[19]));
 sky130_fd_sc_hd__ebufn_8 _1032_ (.A(net37),
    .TE_B(_0287_),
    .Z(la1_data_out[20]));
 sky130_fd_sc_hd__ebufn_8 _1033_ (.A(net38),
    .TE_B(_0288_),
    .Z(la1_data_out[21]));
 sky130_fd_sc_hd__ebufn_8 _1034_ (.A(net39),
    .TE_B(_0289_),
    .Z(la1_data_out[22]));
 sky130_fd_sc_hd__ebufn_8 _1035_ (.A(net40),
    .TE_B(_0290_),
    .Z(la1_data_out[23]));
 sky130_fd_sc_hd__ebufn_8 _1036_ (.A(net41),
    .TE_B(_0291_),
    .Z(la1_data_out[24]));
 sky130_fd_sc_hd__ebufn_8 _1037_ (.A(net42),
    .TE_B(_0292_),
    .Z(la1_data_out[25]));
 sky130_fd_sc_hd__ebufn_8 _1038_ (.A(net43),
    .TE_B(_0293_),
    .Z(la1_data_out[26]));
 sky130_fd_sc_hd__ebufn_8 _1039_ (.A(net44),
    .TE_B(_0294_),
    .Z(la1_data_out[27]));
 sky130_fd_sc_hd__ebufn_8 _1040_ (.A(net45),
    .TE_B(_0295_),
    .Z(la1_data_out[28]));
 sky130_fd_sc_hd__ebufn_8 _1041_ (.A(net46),
    .TE_B(_0296_),
    .Z(la1_data_out[29]));
 sky130_fd_sc_hd__ebufn_8 _1042_ (.A(net47),
    .TE_B(_0297_),
    .Z(la1_data_out[30]));
 sky130_fd_sc_hd__ebufn_8 _1043_ (.A(net48),
    .TE_B(_0298_),
    .Z(la1_data_out[31]));
 sky130_fd_sc_hd__ebufn_8 _1044_ (.A(net49),
    .TE_B(_0299_),
    .Z(io_out[0]));
 sky130_fd_sc_hd__ebufn_8 _1045_ (.A(net50),
    .TE_B(_0300_),
    .Z(io_out[1]));
 sky130_fd_sc_hd__ebufn_8 _1046_ (.A(net51),
    .TE_B(_0301_),
    .Z(io_out[2]));
 sky130_fd_sc_hd__ebufn_8 _1047_ (.A(net52),
    .TE_B(_0302_),
    .Z(io_out[3]));
 sky130_fd_sc_hd__ebufn_8 _1048_ (.A(net53),
    .TE_B(_0303_),
    .Z(io_out[4]));
 sky130_fd_sc_hd__ebufn_8 _1049_ (.A(net54),
    .TE_B(_0304_),
    .Z(io_out[5]));
 sky130_fd_sc_hd__ebufn_8 _1050_ (.A(net55),
    .TE_B(_0305_),
    .Z(io_out[6]));
 sky130_fd_sc_hd__ebufn_8 _1051_ (.A(net56),
    .TE_B(_0306_),
    .Z(io_out[7]));
 sky130_fd_sc_hd__ebufn_8 _1052_ (.A(net57),
    .TE_B(_0307_),
    .Z(io_out[8]));
 sky130_fd_sc_hd__ebufn_8 _1053_ (.A(\frequency_counter_0.segments[0] ),
    .TE_B(_0308_),
    .Z(io_out[9]));
 sky130_fd_sc_hd__ebufn_8 _1054_ (.A(\frequency_counter_0.segments[1] ),
    .TE_B(_0309_),
    .Z(io_out[10]));
 sky130_fd_sc_hd__ebufn_8 _1055_ (.A(\frequency_counter_0.segments[2] ),
    .TE_B(_0310_),
    .Z(io_out[11]));
 sky130_fd_sc_hd__ebufn_8 _1056_ (.A(\frequency_counter_0.segments[3] ),
    .TE_B(_0311_),
    .Z(io_out[12]));
 sky130_fd_sc_hd__ebufn_8 _1057_ (.A(\frequency_counter_0.segments[4] ),
    .TE_B(_0312_),
    .Z(io_out[13]));
 sky130_fd_sc_hd__ebufn_8 _1058_ (.A(\frequency_counter_0.segments[5] ),
    .TE_B(_0313_),
    .Z(io_out[14]));
 sky130_fd_sc_hd__ebufn_8 _1059_ (.A(\frequency_counter_0.segments[6] ),
    .TE_B(_0314_),
    .Z(io_out[15]));
 sky130_fd_sc_hd__ebufn_8 _1060_ (.A(\frequency_counter_0.digit ),
    .TE_B(_0315_),
    .Z(io_out[16]));
 sky130_fd_sc_hd__ebufn_8 _1061_ (.A(net58),
    .TE_B(_0316_),
    .Z(io_out[17]));
 sky130_fd_sc_hd__ebufn_8 _1062_ (.A(net59),
    .TE_B(_0317_),
    .Z(io_out[18]));
 sky130_fd_sc_hd__ebufn_8 _1063_ (.A(net60),
    .TE_B(_0318_),
    .Z(io_out[19]));
 sky130_fd_sc_hd__ebufn_8 _1064_ (.A(net61),
    .TE_B(_0319_),
    .Z(io_out[20]));
 sky130_fd_sc_hd__ebufn_8 _1065_ (.A(net62),
    .TE_B(_0320_),
    .Z(io_out[21]));
 sky130_fd_sc_hd__ebufn_8 _1066_ (.A(net63),
    .TE_B(_0321_),
    .Z(io_out[22]));
 sky130_fd_sc_hd__ebufn_8 _1067_ (.A(net64),
    .TE_B(_0322_),
    .Z(io_out[23]));
 sky130_fd_sc_hd__ebufn_8 _1068_ (.A(net65),
    .TE_B(_0323_),
    .Z(io_out[24]));
 sky130_fd_sc_hd__ebufn_8 _1069_ (.A(net66),
    .TE_B(_0324_),
    .Z(io_out[25]));
 sky130_fd_sc_hd__ebufn_8 _1070_ (.A(net67),
    .TE_B(_0325_),
    .Z(io_out[26]));
 sky130_fd_sc_hd__ebufn_8 _1071_ (.A(net68),
    .TE_B(_0326_),
    .Z(io_out[27]));
 sky130_fd_sc_hd__ebufn_8 _1072_ (.A(net69),
    .TE_B(_0327_),
    .Z(io_out[28]));
 sky130_fd_sc_hd__ebufn_8 _1073_ (.A(net70),
    .TE_B(_0328_),
    .Z(io_out[29]));
 sky130_fd_sc_hd__ebufn_8 _1074_ (.A(net71),
    .TE_B(_0329_),
    .Z(io_out[30]));
 sky130_fd_sc_hd__ebufn_8 _1075_ (.A(net72),
    .TE_B(_0330_),
    .Z(io_out[31]));
 sky130_fd_sc_hd__ebufn_8 _1076_ (.A(net73),
    .TE_B(_0331_),
    .Z(io_out[32]));
 sky130_fd_sc_hd__ebufn_8 _1077_ (.A(net74),
    .TE_B(_0332_),
    .Z(io_out[33]));
 sky130_fd_sc_hd__ebufn_8 _1078_ (.A(net75),
    .TE_B(_0333_),
    .Z(io_out[34]));
 sky130_fd_sc_hd__ebufn_8 _1079_ (.A(net76),
    .TE_B(_0334_),
    .Z(io_out[35]));
 sky130_fd_sc_hd__ebufn_8 _1080_ (.A(net77),
    .TE_B(_0335_),
    .Z(io_out[36]));
 sky130_fd_sc_hd__ebufn_8 _1081_ (.A(net78),
    .TE_B(_0336_),
    .Z(io_out[37]));
 sky130_fd_sc_hd__ebufn_8 _1082_ (.A(net79),
    .TE_B(_0337_),
    .Z(io_oeb[0]));
 sky130_fd_sc_hd__ebufn_8 _1083_ (.A(net80),
    .TE_B(_0338_),
    .Z(io_oeb[1]));
 sky130_fd_sc_hd__ebufn_8 _1084_ (.A(net81),
    .TE_B(_0339_),
    .Z(io_oeb[2]));
 sky130_fd_sc_hd__ebufn_8 _1085_ (.A(net82),
    .TE_B(_0340_),
    .Z(io_oeb[3]));
 sky130_fd_sc_hd__ebufn_8 _1086_ (.A(net83),
    .TE_B(_0341_),
    .Z(io_oeb[4]));
 sky130_fd_sc_hd__ebufn_8 _1087_ (.A(net84),
    .TE_B(_0342_),
    .Z(io_oeb[5]));
 sky130_fd_sc_hd__ebufn_8 _1088_ (.A(net85),
    .TE_B(_0343_),
    .Z(io_oeb[6]));
 sky130_fd_sc_hd__ebufn_8 _1089_ (.A(net86),
    .TE_B(_0344_),
    .Z(io_oeb[7]));
 sky130_fd_sc_hd__ebufn_8 _1090_ (.A(net87),
    .TE_B(_0345_),
    .Z(io_oeb[8]));
 sky130_fd_sc_hd__ebufn_8 _1091_ (.A(net88),
    .TE_B(_0346_),
    .Z(io_oeb[9]));
 sky130_fd_sc_hd__ebufn_8 _1092_ (.A(net89),
    .TE_B(_0347_),
    .Z(io_oeb[10]));
 sky130_fd_sc_hd__ebufn_8 _1093_ (.A(net90),
    .TE_B(_0348_),
    .Z(io_oeb[11]));
 sky130_fd_sc_hd__ebufn_8 _1094_ (.A(net91),
    .TE_B(_0349_),
    .Z(io_oeb[12]));
 sky130_fd_sc_hd__ebufn_8 _1095_ (.A(net92),
    .TE_B(_0350_),
    .Z(io_oeb[13]));
 sky130_fd_sc_hd__ebufn_8 _1096_ (.A(net93),
    .TE_B(_0351_),
    .Z(io_oeb[14]));
 sky130_fd_sc_hd__ebufn_8 _1097_ (.A(net94),
    .TE_B(_0352_),
    .Z(io_oeb[15]));
 sky130_fd_sc_hd__ebufn_8 _1098_ (.A(net95),
    .TE_B(_0353_),
    .Z(io_oeb[16]));
 sky130_fd_sc_hd__ebufn_8 _1099_ (.A(net96),
    .TE_B(_0354_),
    .Z(io_oeb[17]));
 sky130_fd_sc_hd__ebufn_8 _1100_ (.A(net97),
    .TE_B(_0355_),
    .Z(io_oeb[18]));
 sky130_fd_sc_hd__ebufn_8 _1101_ (.A(net98),
    .TE_B(_0356_),
    .Z(io_oeb[19]));
 sky130_fd_sc_hd__ebufn_8 _1102_ (.A(net99),
    .TE_B(_0357_),
    .Z(io_oeb[20]));
 sky130_fd_sc_hd__ebufn_8 _1103_ (.A(net100),
    .TE_B(_0358_),
    .Z(io_oeb[21]));
 sky130_fd_sc_hd__ebufn_8 _1104_ (.A(net101),
    .TE_B(_0359_),
    .Z(io_oeb[22]));
 sky130_fd_sc_hd__ebufn_8 _1105_ (.A(net102),
    .TE_B(_0360_),
    .Z(io_oeb[23]));
 sky130_fd_sc_hd__ebufn_8 _1106_ (.A(net103),
    .TE_B(_0361_),
    .Z(io_oeb[24]));
 sky130_fd_sc_hd__ebufn_8 _1107_ (.A(net104),
    .TE_B(_0362_),
    .Z(io_oeb[25]));
 sky130_fd_sc_hd__ebufn_8 _1108_ (.A(net105),
    .TE_B(_0363_),
    .Z(io_oeb[26]));
 sky130_fd_sc_hd__ebufn_8 _1109_ (.A(net106),
    .TE_B(_0364_),
    .Z(io_oeb[27]));
 sky130_fd_sc_hd__ebufn_8 _1110_ (.A(net107),
    .TE_B(_0365_),
    .Z(io_oeb[28]));
 sky130_fd_sc_hd__ebufn_8 _1111_ (.A(net108),
    .TE_B(_0366_),
    .Z(io_oeb[29]));
 sky130_fd_sc_hd__ebufn_8 _1112_ (.A(net109),
    .TE_B(_0367_),
    .Z(io_oeb[30]));
 sky130_fd_sc_hd__ebufn_8 _1113_ (.A(net110),
    .TE_B(_0368_),
    .Z(io_oeb[31]));
 sky130_fd_sc_hd__ebufn_8 _1114_ (.A(net111),
    .TE_B(_0369_),
    .Z(io_oeb[32]));
 sky130_fd_sc_hd__ebufn_8 _1115_ (.A(net112),
    .TE_B(_0370_),
    .Z(io_oeb[33]));
 sky130_fd_sc_hd__ebufn_8 _1116_ (.A(net113),
    .TE_B(_0371_),
    .Z(io_oeb[34]));
 sky130_fd_sc_hd__ebufn_8 _1117_ (.A(net114),
    .TE_B(_0372_),
    .Z(io_oeb[35]));
 sky130_fd_sc_hd__ebufn_8 _1118_ (.A(net115),
    .TE_B(_0373_),
    .Z(io_oeb[36]));
 sky130_fd_sc_hd__ebufn_8 _1119_ (.A(net116),
    .TE_B(_0374_),
    .Z(io_oeb[37]));
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__decap_3 PHY_162 ();
 sky130_fd_sc_hd__decap_3 PHY_163 ();
 sky130_fd_sc_hd__decap_3 PHY_164 ();
 sky130_fd_sc_hd__decap_3 PHY_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__clkbuf_1 input1 (.A(active),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(io_in[8]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(la1_data_in[0]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(la1_data_in[10]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(la1_data_in[11]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(la1_data_in[12]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_1 input7 (.A(la1_data_in[13]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_2 input8 (.A(la1_data_in[1]),
    .X(net8));
 sky130_fd_sc_hd__dlymetal6s2s_1 input9 (.A(la1_data_in[2]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_1 input10 (.A(la1_data_in[3]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_1 input11 (.A(la1_data_in[4]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_1 input12 (.A(la1_data_in[5]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_1 input13 (.A(la1_data_in[6]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_1 input14 (.A(la1_data_in[7]),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_1 input15 (.A(la1_data_in[8]),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_1 input16 (.A(la1_data_in[9]),
    .X(net16));
 sky130_fd_sc_hd__conb_1 _1012__17 (.LO(net17));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_0__f_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_2_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_1__f_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_2_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_2__f_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_2_2__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_3__f_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_2_3__leaf_wb_clk_i));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1 (.A(\frequency_counter_0.edge_detect0.q0 ),
    .X(net117));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(\frequency_counter_0.edge_detect0.q1 ),
    .X(net118));
 sky130_fd_sc_hd__fill_2 FILLER_0_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_286 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_10 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_24 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_84 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_196 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_248 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_286 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_72 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_90 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_180 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_117 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_127 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_40 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_286 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_49 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_10 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_286 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_16 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_58 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_10 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_286 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_17 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_204 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_286 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_10 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_43 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_212 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_238 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_247 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_190 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_238 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_295 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_28 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_185 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_204 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_176 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_298 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_107 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_187 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_199 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_10 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_236 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_28 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_148 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_200 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_270 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_142 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_184 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_246 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_260 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_10 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_208 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_236 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_196 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_136 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_28 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_189 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_236 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_201 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_224 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_187 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_220 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_232 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_246 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_217 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_232 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_247 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_12 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_168 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_208 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_286 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_10 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_258 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_174 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_268 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_286 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_168 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_229 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_246 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_263 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_170 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_238 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_246 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_213 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_236 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_248 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_297 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_159 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_171 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_229 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_246 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_204 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_257 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_10 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_190 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_199 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_243 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_298 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_235 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_10 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_43 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_176 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_286 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_10 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_43 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_191 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_286 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_10 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_10 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_298 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_10 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_10 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_297 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_272 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_286 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_96 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_208 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_70 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_130 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_168 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_140 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_192 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_286 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_70 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_118 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_126 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_186 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_286 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_293 ();
endmodule

