VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO wrapped_frequency_counter
  CLASS BLOCK ;
  FOREIGN wrapped_frequency_counter ;
  ORIGIN 0.000 0.000 ;
  SIZE 150.000 BY 210.000 ;
  PIN active
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 194.520 4.000 195.120 ;
    END
  END active
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.090 0.000 46.370 4.000 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.810 206.000 84.090 210.000 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.010 206.000 1.290 210.000 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 176.840 150.000 177.440 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.930 0.000 71.210 4.000 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.210 206.000 56.490 210.000 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 185.000 150.000 185.600 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 17.720 150.000 18.320 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.370 206.000 31.650 210.000 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.890 206.000 37.170 210.000 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.890 0.000 129.170 4.000 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.040 4.000 68.640 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 121.080 4.000 121.680 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 80.280 4.000 80.880 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 66.680 150.000 67.280 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.610 206.000 28.890 210.000 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.330 206.000 20.610 210.000 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.330 0.000 112.610 4.000 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.570 0.000 109.850 4.000 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 46.280 150.000 46.880 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.530 0.000 98.810 4.000 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 149.130 206.000 149.410 210.000 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.850 0.000 49.130 4.000 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 83.000 150.000 83.600 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 186.360 4.000 186.960 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.010 0.000 93.290 4.000 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 108.840 4.000 109.440 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 114.170 206.000 114.450 210.000 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 130.730 206.000 131.010 210.000 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 131.960 150.000 132.560 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.490 206.000 133.770 210.000 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 86.570 206.000 86.850 210.000 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 127.880 150.000 128.480 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 201.320 150.000 201.920 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 129.240 4.000 129.840 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 88.440 4.000 89.040 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 140.120 150.000 140.720 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.850 206.000 26.130 210.000 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.210 0.000 79.490 4.000 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 72.120 4.000 72.720 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 119.720 150.000 120.320 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 62.600 150.000 63.200 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 58.520 150.000 59.120 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 19.080 4.000 19.680 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.410 206.000 42.690 210.000 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 9.560 150.000 10.160 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.570 0.000 40.850 4.000 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 108.650 206.000 108.930 210.000 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.170 206.000 45.450 210.000 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 117.850 0.000 118.130 4.000 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 91.160 150.000 91.760 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.530 206.000 6.810 210.000 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 15.730 0.000 16.010 4.000 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.530 206.000 75.810 210.000 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.290 206.000 78.570 210.000 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 142.690 0.000 142.970 4.000 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 164.600 150.000 165.200 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.330 206.000 89.610 210.000 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 126.130 0.000 126.410 4.000 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 136.040 150.000 136.640 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.210 206.000 125.490 210.000 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.290 206.000 9.570 210.000 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 123.370 0.000 123.650 4.000 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 104.760 4.000 105.360 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 145.450 0.000 145.730 4.000 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.130 206.000 34.410 210.000 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 92.520 4.000 93.120 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 47.640 4.000 48.240 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 76.200 4.000 76.800 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.450 0.000 76.730 4.000 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 1.400 150.000 2.000 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 137.400 4.000 138.000 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 74.840 150.000 75.440 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.650 206.000 39.930 210.000 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.970 0.000 13.250 4.000 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.290 0.000 32.570 4.000 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 197.240 150.000 197.840 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 115.640 150.000 116.240 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 10.920 4.000 11.520 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 31.320 4.000 31.920 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 120.610 0.000 120.890 4.000 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 168.680 150.000 169.280 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 174.120 4.000 174.720 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 111.560 150.000 112.160 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.010 206.000 139.290 210.000 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.930 0.000 140.210 4.000 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 100.680 4.000 101.280 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 100.370 206.000 100.650 210.000 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.450 206.000 122.730 210.000 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 170.040 4.000 170.640 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 95.770 0.000 96.050 4.000 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 95.240 150.000 95.840 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.970 0.000 82.250 4.000 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 111.410 206.000 111.690 210.000 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 23.160 4.000 23.760 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.930 206.000 117.210 210.000 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.610 0.000 51.890 4.000 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 5.480 150.000 6.080 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.250 0.000 21.530 4.000 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.240 4.000 27.840 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 59.880 4.000 60.480 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 198.600 4.000 199.200 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 29.960 150.000 30.560 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 172.760 150.000 173.360 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 160.520 150.000 161.120 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.930 206.000 48.210 210.000 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 189.080 150.000 189.680 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 182.280 4.000 182.880 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 123.800 150.000 124.400 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.010 206.000 70.290 210.000 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.530 206.000 144.810 210.000 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 84.360 4.000 84.960 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.130 0.000 57.410 4.000 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 63.960 4.000 64.560 ;
    END
  END io_out[9]
  PIN la1_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 34.040 150.000 34.640 ;
    END
  END la1_data_in[0]
  PIN la1_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.410 0.000 65.690 4.000 ;
    END
  END la1_data_in[10]
  PIN la1_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 25.880 150.000 26.480 ;
    END
  END la1_data_in[11]
  PIN la1_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 157.800 4.000 158.400 ;
    END
  END la1_data_in[12]
  PIN la1_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 101.290 0.000 101.570 4.000 ;
    END
  END la1_data_in[13]
  PIN la1_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 55.800 4.000 56.400 ;
    END
  END la1_data_in[14]
  PIN la1_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.690 206.000 50.970 210.000 ;
    END
  END la1_data_in[15]
  PIN la1_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.850 206.000 95.130 210.000 ;
    END
  END la1_data_in[16]
  PIN la1_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.770 206.000 73.050 210.000 ;
    END
  END la1_data_in[17]
  PIN la1_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 131.650 0.000 131.930 4.000 ;
    END
  END la1_data_in[18]
  PIN la1_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.450 206.000 53.730 210.000 ;
    END
  END la1_data_in[19]
  PIN la1_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.890 0.000 60.170 4.000 ;
    END
  END la1_data_in[1]
  PIN la1_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 153.720 4.000 154.320 ;
    END
  END la1_data_in[20]
  PIN la1_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 147.290 206.000 147.570 210.000 ;
    END
  END la1_data_in[21]
  PIN la1_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 38.120 150.000 38.720 ;
    END
  END la1_data_in[22]
  PIN la1_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2.760 4.000 3.360 ;
    END
  END la1_data_in[23]
  PIN la1_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.330 0.000 43.610 4.000 ;
    END
  END la1_data_in[24]
  PIN la1_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 161.880 4.000 162.480 ;
    END
  END la1_data_in[25]
  PIN la1_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 13.640 150.000 14.240 ;
    END
  END la1_data_in[26]
  PIN la1_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.490 0.000 87.770 4.000 ;
    END
  END la1_data_in[27]
  PIN la1_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 141.480 4.000 142.080 ;
    END
  END la1_data_in[28]
  PIN la1_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.770 206.000 4.050 210.000 ;
    END
  END la1_data_in[29]
  PIN la1_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.050 0.000 35.330 4.000 ;
    END
  END la1_data_in[2]
  PIN la1_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.690 0.000 4.970 4.000 ;
    END
  END la1_data_in[30]
  PIN la1_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 115.090 0.000 115.370 4.000 ;
    END
  END la1_data_in[31]
  PIN la1_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 133.320 4.000 133.920 ;
    END
  END la1_data_in[3]
  PIN la1_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.970 206.000 128.250 210.000 ;
    END
  END la1_data_in[4]
  PIN la1_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 103.400 150.000 104.000 ;
    END
  END la1_data_in[5]
  PIN la1_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.970 206.000 59.250 210.000 ;
    END
  END la1_data_in[6]
  PIN la1_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 96.600 4.000 97.200 ;
    END
  END la1_data_in[7]
  PIN la1_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.730 206.000 62.010 210.000 ;
    END
  END la1_data_in[8]
  PIN la1_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 145.560 4.000 146.160 ;
    END
  END la1_data_in[9]
  PIN la1_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.010 0.000 24.290 4.000 ;
    END
  END la1_data_out[0]
  PIN la1_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 50.360 150.000 50.960 ;
    END
  END la1_data_out[10]
  PIN la1_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.170 0.000 68.450 4.000 ;
    END
  END la1_data_out[11]
  PIN la1_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 193.160 150.000 193.760 ;
    END
  END la1_data_out[12]
  PIN la1_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.810 206.000 15.090 210.000 ;
    END
  END la1_data_out[13]
  PIN la1_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.050 206.000 81.330 210.000 ;
    END
  END la1_data_out[14]
  PIN la1_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 6.840 4.000 7.440 ;
    END
  END la1_data_out[15]
  PIN la1_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 70.760 150.000 71.360 ;
    END
  END la1_data_out[16]
  PIN la1_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 152.360 150.000 152.960 ;
    END
  END la1_data_out[17]
  PIN la1_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.570 206.000 17.850 210.000 ;
    END
  END la1_data_out[18]
  PIN la1_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 107.480 150.000 108.080 ;
    END
  END la1_data_out[19]
  PIN la1_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 190.440 4.000 191.040 ;
    END
  END la1_data_out[1]
  PIN la1_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 43.560 4.000 44.160 ;
    END
  END la1_data_out[20]
  PIN la1_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 180.920 150.000 181.520 ;
    END
  END la1_data_out[21]
  PIN la1_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 92.090 206.000 92.370 210.000 ;
    END
  END la1_data_out[22]
  PIN la1_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.810 0.000 38.090 4.000 ;
    END
  END la1_data_out[23]
  PIN la1_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 78.920 150.000 79.520 ;
    END
  END la1_data_out[24]
  PIN la1_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 15.000 4.000 15.600 ;
    END
  END la1_data_out[25]
  PIN la1_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 21.800 150.000 22.400 ;
    END
  END la1_data_out[26]
  PIN la1_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 202.680 4.000 203.280 ;
    END
  END la1_data_out[27]
  PIN la1_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 134.410 0.000 134.690 4.000 ;
    END
  END la1_data_out[28]
  PIN la1_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.490 0.000 18.770 4.000 ;
    END
  END la1_data_out[29]
  PIN la1_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.650 0.000 62.930 4.000 ;
    END
  END la1_data_out[2]
  PIN la1_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 54.440 150.000 55.040 ;
    END
  END la1_data_out[30]
  PIN la1_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 205.400 150.000 206.000 ;
    END
  END la1_data_out[31]
  PIN la1_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 39.480 4.000 40.080 ;
    END
  END la1_data_out[3]
  PIN la1_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 137.170 0.000 137.450 4.000 ;
    END
  END la1_data_out[4]
  PIN la1_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.210 0.000 10.490 4.000 ;
    END
  END la1_data_out[5]
  PIN la1_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 87.080 150.000 87.680 ;
    END
  END la1_data_out[6]
  PIN la1_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.930 0.000 2.210 4.000 ;
    END
  END la1_data_out[7]
  PIN la1_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 156.440 150.000 157.040 ;
    END
  END la1_data_out[8]
  PIN la1_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 141.770 206.000 142.050 210.000 ;
    END
  END la1_data_out[9]
  PIN la1_oenb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.210 0.000 148.490 4.000 ;
    END
  END la1_oenb[0]
  PIN la1_oenb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 136.250 206.000 136.530 210.000 ;
    END
  END la1_oenb[10]
  PIN la1_oenb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 117.000 4.000 117.600 ;
    END
  END la1_oenb[11]
  PIN la1_oenb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 125.160 4.000 125.760 ;
    END
  END la1_oenb[12]
  PIN la1_oenb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.250 0.000 90.530 4.000 ;
    END
  END la1_oenb[13]
  PIN la1_oenb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END la1_oenb[14]
  PIN la1_oenb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.810 0.000 107.090 4.000 ;
    END
  END la1_oenb[15]
  PIN la1_oenb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 149.640 4.000 150.240 ;
    END
  END la1_oenb[16]
  PIN la1_oenb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.050 206.000 12.330 210.000 ;
    END
  END la1_oenb[17]
  PIN la1_oenb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.250 206.000 67.530 210.000 ;
    END
  END la1_oenb[18]
  PIN la1_oenb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 112.920 4.000 113.520 ;
    END
  END la1_oenb[19]
  PIN la1_oenb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.770 0.000 27.050 4.000 ;
    END
  END la1_oenb[1]
  PIN la1_oenb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.450 0.000 7.730 4.000 ;
    END
  END la1_oenb[20]
  PIN la1_oenb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 97.610 206.000 97.890 210.000 ;
    END
  END la1_oenb[21]
  PIN la1_oenb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.490 206.000 64.770 210.000 ;
    END
  END la1_oenb[22]
  PIN la1_oenb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.690 0.000 73.970 4.000 ;
    END
  END la1_oenb[23]
  PIN la1_oenb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.690 206.000 119.970 210.000 ;
    END
  END la1_oenb[24]
  PIN la1_oenb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 42.200 150.000 42.800 ;
    END
  END la1_oenb[25]
  PIN la1_oenb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 165.960 4.000 166.560 ;
    END
  END la1_oenb[26]
  PIN la1_oenb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 148.280 150.000 148.880 ;
    END
  END la1_oenb[27]
  PIN la1_oenb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.530 0.000 29.810 4.000 ;
    END
  END la1_oenb[28]
  PIN la1_oenb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.370 0.000 54.650 4.000 ;
    END
  END la1_oenb[29]
  PIN la1_oenb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 35.400 4.000 36.000 ;
    END
  END la1_oenb[2]
  PIN la1_oenb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 144.200 150.000 144.800 ;
    END
  END la1_oenb[30]
  PIN la1_oenb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 84.730 0.000 85.010 4.000 ;
    END
  END la1_oenb[31]
  PIN la1_oenb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 105.890 206.000 106.170 210.000 ;
    END
  END la1_oenb[3]
  PIN la1_oenb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.130 206.000 103.410 210.000 ;
    END
  END la1_oenb[4]
  PIN la1_oenb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 206.760 4.000 207.360 ;
    END
  END la1_oenb[5]
  PIN la1_oenb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.090 206.000 23.370 210.000 ;
    END
  END la1_oenb[6]
  PIN la1_oenb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.050 0.000 104.330 4.000 ;
    END
  END la1_oenb[7]
  PIN la1_oenb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.720 4.000 52.320 ;
    END
  END la1_oenb[8]
  PIN la1_oenb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 178.200 4.000 178.800 ;
    END
  END la1_oenb[9]
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 27.875 10.640 29.475 198.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 74.195 10.640 75.795 198.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 120.515 10.640 122.115 198.800 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 51.035 10.640 52.635 198.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 97.355 10.640 98.955 198.800 ;
    END
  END vssd1
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 99.320 150.000 99.920 ;
    END
  END wb_clk_i
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 146.595 198.645 ;
      LAYER met1 ;
        RECT 1.910 10.640 146.655 198.800 ;
      LAYER met2 ;
        RECT 1.940 205.720 3.490 206.450 ;
        RECT 4.330 205.720 6.250 206.450 ;
        RECT 7.090 205.720 9.010 206.450 ;
        RECT 9.850 205.720 11.770 206.450 ;
        RECT 12.610 205.720 14.530 206.450 ;
        RECT 15.370 205.720 17.290 206.450 ;
        RECT 18.130 205.720 20.050 206.450 ;
        RECT 20.890 205.720 22.810 206.450 ;
        RECT 23.650 205.720 25.570 206.450 ;
        RECT 26.410 205.720 28.330 206.450 ;
        RECT 29.170 205.720 31.090 206.450 ;
        RECT 31.930 205.720 33.850 206.450 ;
        RECT 34.690 205.720 36.610 206.450 ;
        RECT 37.450 205.720 39.370 206.450 ;
        RECT 40.210 205.720 42.130 206.450 ;
        RECT 42.970 205.720 44.890 206.450 ;
        RECT 45.730 205.720 47.650 206.450 ;
        RECT 48.490 205.720 50.410 206.450 ;
        RECT 51.250 205.720 53.170 206.450 ;
        RECT 54.010 205.720 55.930 206.450 ;
        RECT 56.770 205.720 58.690 206.450 ;
        RECT 59.530 205.720 61.450 206.450 ;
        RECT 62.290 205.720 64.210 206.450 ;
        RECT 65.050 205.720 66.970 206.450 ;
        RECT 67.810 205.720 69.730 206.450 ;
        RECT 70.570 205.720 72.490 206.450 ;
        RECT 73.330 205.720 75.250 206.450 ;
        RECT 76.090 205.720 78.010 206.450 ;
        RECT 78.850 205.720 80.770 206.450 ;
        RECT 81.610 205.720 83.530 206.450 ;
        RECT 84.370 205.720 86.290 206.450 ;
        RECT 87.130 205.720 89.050 206.450 ;
        RECT 89.890 205.720 91.810 206.450 ;
        RECT 92.650 205.720 94.570 206.450 ;
        RECT 95.410 205.720 97.330 206.450 ;
        RECT 98.170 205.720 100.090 206.450 ;
        RECT 100.930 205.720 102.850 206.450 ;
        RECT 103.690 205.720 105.610 206.450 ;
        RECT 106.450 205.720 108.370 206.450 ;
        RECT 109.210 205.720 111.130 206.450 ;
        RECT 111.970 205.720 113.890 206.450 ;
        RECT 114.730 205.720 116.650 206.450 ;
        RECT 117.490 205.720 119.410 206.450 ;
        RECT 120.250 205.720 122.170 206.450 ;
        RECT 123.010 205.720 124.930 206.450 ;
        RECT 125.770 205.720 127.690 206.450 ;
        RECT 128.530 205.720 130.450 206.450 ;
        RECT 131.290 205.720 133.210 206.450 ;
        RECT 134.050 205.720 135.970 206.450 ;
        RECT 136.810 205.720 138.730 206.450 ;
        RECT 139.570 205.720 141.490 206.450 ;
        RECT 142.330 205.720 144.250 206.450 ;
        RECT 145.090 205.720 145.720 206.450 ;
        RECT 1.940 4.280 145.720 205.720 ;
        RECT 2.490 1.515 4.410 4.280 ;
        RECT 5.250 1.515 7.170 4.280 ;
        RECT 8.010 1.515 9.930 4.280 ;
        RECT 10.770 1.515 12.690 4.280 ;
        RECT 13.530 1.515 15.450 4.280 ;
        RECT 16.290 1.515 18.210 4.280 ;
        RECT 19.050 1.515 20.970 4.280 ;
        RECT 21.810 1.515 23.730 4.280 ;
        RECT 24.570 1.515 26.490 4.280 ;
        RECT 27.330 1.515 29.250 4.280 ;
        RECT 30.090 1.515 32.010 4.280 ;
        RECT 32.850 1.515 34.770 4.280 ;
        RECT 35.610 1.515 37.530 4.280 ;
        RECT 38.370 1.515 40.290 4.280 ;
        RECT 41.130 1.515 43.050 4.280 ;
        RECT 43.890 1.515 45.810 4.280 ;
        RECT 46.650 1.515 48.570 4.280 ;
        RECT 49.410 1.515 51.330 4.280 ;
        RECT 52.170 1.515 54.090 4.280 ;
        RECT 54.930 1.515 56.850 4.280 ;
        RECT 57.690 1.515 59.610 4.280 ;
        RECT 60.450 1.515 62.370 4.280 ;
        RECT 63.210 1.515 65.130 4.280 ;
        RECT 65.970 1.515 67.890 4.280 ;
        RECT 68.730 1.515 70.650 4.280 ;
        RECT 71.490 1.515 73.410 4.280 ;
        RECT 74.250 1.515 76.170 4.280 ;
        RECT 77.010 1.515 78.930 4.280 ;
        RECT 79.770 1.515 81.690 4.280 ;
        RECT 82.530 1.515 84.450 4.280 ;
        RECT 85.290 1.515 87.210 4.280 ;
        RECT 88.050 1.515 89.970 4.280 ;
        RECT 90.810 1.515 92.730 4.280 ;
        RECT 93.570 1.515 95.490 4.280 ;
        RECT 96.330 1.515 98.250 4.280 ;
        RECT 99.090 1.515 101.010 4.280 ;
        RECT 101.850 1.515 103.770 4.280 ;
        RECT 104.610 1.515 106.530 4.280 ;
        RECT 107.370 1.515 109.290 4.280 ;
        RECT 110.130 1.515 112.050 4.280 ;
        RECT 112.890 1.515 114.810 4.280 ;
        RECT 115.650 1.515 117.570 4.280 ;
        RECT 118.410 1.515 120.330 4.280 ;
        RECT 121.170 1.515 123.090 4.280 ;
        RECT 123.930 1.515 125.850 4.280 ;
        RECT 126.690 1.515 128.610 4.280 ;
        RECT 129.450 1.515 131.370 4.280 ;
        RECT 132.210 1.515 134.130 4.280 ;
        RECT 134.970 1.515 136.890 4.280 ;
        RECT 137.730 1.515 139.650 4.280 ;
        RECT 140.490 1.515 142.410 4.280 ;
        RECT 143.250 1.515 145.170 4.280 ;
      LAYER met3 ;
        RECT 4.000 205.000 145.600 205.865 ;
        RECT 4.000 203.680 146.000 205.000 ;
        RECT 4.400 202.320 146.000 203.680 ;
        RECT 4.400 202.280 145.600 202.320 ;
        RECT 4.000 200.920 145.600 202.280 ;
        RECT 4.000 199.600 146.000 200.920 ;
        RECT 4.400 198.240 146.000 199.600 ;
        RECT 4.400 198.200 145.600 198.240 ;
        RECT 4.000 196.840 145.600 198.200 ;
        RECT 4.000 195.520 146.000 196.840 ;
        RECT 4.400 194.160 146.000 195.520 ;
        RECT 4.400 194.120 145.600 194.160 ;
        RECT 4.000 192.760 145.600 194.120 ;
        RECT 4.000 191.440 146.000 192.760 ;
        RECT 4.400 190.080 146.000 191.440 ;
        RECT 4.400 190.040 145.600 190.080 ;
        RECT 4.000 188.680 145.600 190.040 ;
        RECT 4.000 187.360 146.000 188.680 ;
        RECT 4.400 186.000 146.000 187.360 ;
        RECT 4.400 185.960 145.600 186.000 ;
        RECT 4.000 184.600 145.600 185.960 ;
        RECT 4.000 183.280 146.000 184.600 ;
        RECT 4.400 181.920 146.000 183.280 ;
        RECT 4.400 181.880 145.600 181.920 ;
        RECT 4.000 180.520 145.600 181.880 ;
        RECT 4.000 179.200 146.000 180.520 ;
        RECT 4.400 177.840 146.000 179.200 ;
        RECT 4.400 177.800 145.600 177.840 ;
        RECT 4.000 176.440 145.600 177.800 ;
        RECT 4.000 175.120 146.000 176.440 ;
        RECT 4.400 173.760 146.000 175.120 ;
        RECT 4.400 173.720 145.600 173.760 ;
        RECT 4.000 172.360 145.600 173.720 ;
        RECT 4.000 171.040 146.000 172.360 ;
        RECT 4.400 169.680 146.000 171.040 ;
        RECT 4.400 169.640 145.600 169.680 ;
        RECT 4.000 168.280 145.600 169.640 ;
        RECT 4.000 166.960 146.000 168.280 ;
        RECT 4.400 165.600 146.000 166.960 ;
        RECT 4.400 165.560 145.600 165.600 ;
        RECT 4.000 164.200 145.600 165.560 ;
        RECT 4.000 162.880 146.000 164.200 ;
        RECT 4.400 161.520 146.000 162.880 ;
        RECT 4.400 161.480 145.600 161.520 ;
        RECT 4.000 160.120 145.600 161.480 ;
        RECT 4.000 158.800 146.000 160.120 ;
        RECT 4.400 157.440 146.000 158.800 ;
        RECT 4.400 157.400 145.600 157.440 ;
        RECT 4.000 156.040 145.600 157.400 ;
        RECT 4.000 154.720 146.000 156.040 ;
        RECT 4.400 153.360 146.000 154.720 ;
        RECT 4.400 153.320 145.600 153.360 ;
        RECT 4.000 151.960 145.600 153.320 ;
        RECT 4.000 150.640 146.000 151.960 ;
        RECT 4.400 149.280 146.000 150.640 ;
        RECT 4.400 149.240 145.600 149.280 ;
        RECT 4.000 147.880 145.600 149.240 ;
        RECT 4.000 146.560 146.000 147.880 ;
        RECT 4.400 145.200 146.000 146.560 ;
        RECT 4.400 145.160 145.600 145.200 ;
        RECT 4.000 143.800 145.600 145.160 ;
        RECT 4.000 142.480 146.000 143.800 ;
        RECT 4.400 141.120 146.000 142.480 ;
        RECT 4.400 141.080 145.600 141.120 ;
        RECT 4.000 139.720 145.600 141.080 ;
        RECT 4.000 138.400 146.000 139.720 ;
        RECT 4.400 137.040 146.000 138.400 ;
        RECT 4.400 137.000 145.600 137.040 ;
        RECT 4.000 135.640 145.600 137.000 ;
        RECT 4.000 134.320 146.000 135.640 ;
        RECT 4.400 132.960 146.000 134.320 ;
        RECT 4.400 132.920 145.600 132.960 ;
        RECT 4.000 131.560 145.600 132.920 ;
        RECT 4.000 130.240 146.000 131.560 ;
        RECT 4.400 128.880 146.000 130.240 ;
        RECT 4.400 128.840 145.600 128.880 ;
        RECT 4.000 127.480 145.600 128.840 ;
        RECT 4.000 126.160 146.000 127.480 ;
        RECT 4.400 124.800 146.000 126.160 ;
        RECT 4.400 124.760 145.600 124.800 ;
        RECT 4.000 123.400 145.600 124.760 ;
        RECT 4.000 122.080 146.000 123.400 ;
        RECT 4.400 120.720 146.000 122.080 ;
        RECT 4.400 120.680 145.600 120.720 ;
        RECT 4.000 119.320 145.600 120.680 ;
        RECT 4.000 118.000 146.000 119.320 ;
        RECT 4.400 116.640 146.000 118.000 ;
        RECT 4.400 116.600 145.600 116.640 ;
        RECT 4.000 115.240 145.600 116.600 ;
        RECT 4.000 113.920 146.000 115.240 ;
        RECT 4.400 112.560 146.000 113.920 ;
        RECT 4.400 112.520 145.600 112.560 ;
        RECT 4.000 111.160 145.600 112.520 ;
        RECT 4.000 109.840 146.000 111.160 ;
        RECT 4.400 108.480 146.000 109.840 ;
        RECT 4.400 108.440 145.600 108.480 ;
        RECT 4.000 107.080 145.600 108.440 ;
        RECT 4.000 105.760 146.000 107.080 ;
        RECT 4.400 104.400 146.000 105.760 ;
        RECT 4.400 104.360 145.600 104.400 ;
        RECT 4.000 103.000 145.600 104.360 ;
        RECT 4.000 101.680 146.000 103.000 ;
        RECT 4.400 100.320 146.000 101.680 ;
        RECT 4.400 100.280 145.600 100.320 ;
        RECT 4.000 98.920 145.600 100.280 ;
        RECT 4.000 97.600 146.000 98.920 ;
        RECT 4.400 96.240 146.000 97.600 ;
        RECT 4.400 96.200 145.600 96.240 ;
        RECT 4.000 94.840 145.600 96.200 ;
        RECT 4.000 93.520 146.000 94.840 ;
        RECT 4.400 92.160 146.000 93.520 ;
        RECT 4.400 92.120 145.600 92.160 ;
        RECT 4.000 90.760 145.600 92.120 ;
        RECT 4.000 89.440 146.000 90.760 ;
        RECT 4.400 88.080 146.000 89.440 ;
        RECT 4.400 88.040 145.600 88.080 ;
        RECT 4.000 86.680 145.600 88.040 ;
        RECT 4.000 85.360 146.000 86.680 ;
        RECT 4.400 84.000 146.000 85.360 ;
        RECT 4.400 83.960 145.600 84.000 ;
        RECT 4.000 82.600 145.600 83.960 ;
        RECT 4.000 81.280 146.000 82.600 ;
        RECT 4.400 79.920 146.000 81.280 ;
        RECT 4.400 79.880 145.600 79.920 ;
        RECT 4.000 78.520 145.600 79.880 ;
        RECT 4.000 77.200 146.000 78.520 ;
        RECT 4.400 75.840 146.000 77.200 ;
        RECT 4.400 75.800 145.600 75.840 ;
        RECT 4.000 74.440 145.600 75.800 ;
        RECT 4.000 73.120 146.000 74.440 ;
        RECT 4.400 71.760 146.000 73.120 ;
        RECT 4.400 71.720 145.600 71.760 ;
        RECT 4.000 70.360 145.600 71.720 ;
        RECT 4.000 69.040 146.000 70.360 ;
        RECT 4.400 67.680 146.000 69.040 ;
        RECT 4.400 67.640 145.600 67.680 ;
        RECT 4.000 66.280 145.600 67.640 ;
        RECT 4.000 64.960 146.000 66.280 ;
        RECT 4.400 63.600 146.000 64.960 ;
        RECT 4.400 63.560 145.600 63.600 ;
        RECT 4.000 62.200 145.600 63.560 ;
        RECT 4.000 60.880 146.000 62.200 ;
        RECT 4.400 59.520 146.000 60.880 ;
        RECT 4.400 59.480 145.600 59.520 ;
        RECT 4.000 58.120 145.600 59.480 ;
        RECT 4.000 56.800 146.000 58.120 ;
        RECT 4.400 55.440 146.000 56.800 ;
        RECT 4.400 55.400 145.600 55.440 ;
        RECT 4.000 54.040 145.600 55.400 ;
        RECT 4.000 52.720 146.000 54.040 ;
        RECT 4.400 51.360 146.000 52.720 ;
        RECT 4.400 51.320 145.600 51.360 ;
        RECT 4.000 49.960 145.600 51.320 ;
        RECT 4.000 48.640 146.000 49.960 ;
        RECT 4.400 47.280 146.000 48.640 ;
        RECT 4.400 47.240 145.600 47.280 ;
        RECT 4.000 45.880 145.600 47.240 ;
        RECT 4.000 44.560 146.000 45.880 ;
        RECT 4.400 43.200 146.000 44.560 ;
        RECT 4.400 43.160 145.600 43.200 ;
        RECT 4.000 41.800 145.600 43.160 ;
        RECT 4.000 40.480 146.000 41.800 ;
        RECT 4.400 39.120 146.000 40.480 ;
        RECT 4.400 39.080 145.600 39.120 ;
        RECT 4.000 37.720 145.600 39.080 ;
        RECT 4.000 36.400 146.000 37.720 ;
        RECT 4.400 35.040 146.000 36.400 ;
        RECT 4.400 35.000 145.600 35.040 ;
        RECT 4.000 33.640 145.600 35.000 ;
        RECT 4.000 32.320 146.000 33.640 ;
        RECT 4.400 30.960 146.000 32.320 ;
        RECT 4.400 30.920 145.600 30.960 ;
        RECT 4.000 29.560 145.600 30.920 ;
        RECT 4.000 28.240 146.000 29.560 ;
        RECT 4.400 26.880 146.000 28.240 ;
        RECT 4.400 26.840 145.600 26.880 ;
        RECT 4.000 25.480 145.600 26.840 ;
        RECT 4.000 24.160 146.000 25.480 ;
        RECT 4.400 22.800 146.000 24.160 ;
        RECT 4.400 22.760 145.600 22.800 ;
        RECT 4.000 21.400 145.600 22.760 ;
        RECT 4.000 20.080 146.000 21.400 ;
        RECT 4.400 18.720 146.000 20.080 ;
        RECT 4.400 18.680 145.600 18.720 ;
        RECT 4.000 17.320 145.600 18.680 ;
        RECT 4.000 16.000 146.000 17.320 ;
        RECT 4.400 14.640 146.000 16.000 ;
        RECT 4.400 14.600 145.600 14.640 ;
        RECT 4.000 13.240 145.600 14.600 ;
        RECT 4.000 11.920 146.000 13.240 ;
        RECT 4.400 10.560 146.000 11.920 ;
        RECT 4.400 10.520 145.600 10.560 ;
        RECT 4.000 9.160 145.600 10.520 ;
        RECT 4.000 7.840 146.000 9.160 ;
        RECT 4.400 6.480 146.000 7.840 ;
        RECT 4.400 6.440 145.600 6.480 ;
        RECT 4.000 5.080 145.600 6.440 ;
        RECT 4.000 3.760 146.000 5.080 ;
        RECT 4.400 2.400 146.000 3.760 ;
        RECT 4.400 2.360 145.600 2.400 ;
        RECT 4.000 1.535 145.600 2.360 ;
      LAYER met4 ;
        RECT 29.875 10.640 50.635 198.800 ;
        RECT 53.035 10.640 72.385 198.800 ;
  END
END wrapped_frequency_counter
END LIBRARY

