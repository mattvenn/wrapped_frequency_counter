magic
tech sky130A
magscale 1 2
timestamp 1647448631
<< viali >>
rect 1409 17221 1443 17255
rect 3985 17221 4019 17255
rect 9137 17221 9171 17255
rect 11989 17221 12023 17255
rect 23857 17221 23891 17255
rect 39129 17221 39163 17255
rect 47041 17221 47075 17255
rect 19993 17153 20027 17187
rect 3065 17085 3099 17119
rect 3249 17085 3283 17119
rect 5641 17085 5675 17119
rect 5825 17085 5859 17119
rect 6561 17085 6595 17119
rect 6745 17085 6779 17119
rect 7757 17085 7791 17119
rect 8953 17085 8987 17119
rect 9413 17085 9447 17119
rect 13001 17085 13035 17119
rect 14105 17085 14139 17119
rect 14289 17085 14323 17119
rect 15485 17085 15519 17119
rect 17877 17085 17911 17119
rect 18521 17085 18555 17119
rect 18705 17085 18739 17119
rect 19257 17085 19291 17119
rect 21281 17085 21315 17119
rect 22017 17085 22051 17119
rect 22201 17085 22235 17119
rect 24409 17085 24443 17119
rect 24593 17085 24627 17119
rect 24869 17085 24903 17119
rect 27169 17085 27203 17119
rect 27353 17085 27387 17119
rect 29009 17085 29043 17119
rect 29745 17085 29779 17119
rect 29929 17085 29963 17119
rect 30941 17085 30975 17119
rect 32137 17085 32171 17119
rect 32321 17085 32355 17119
rect 32597 17085 32631 17119
rect 34713 17085 34747 17119
rect 34897 17085 34931 17119
rect 35173 17085 35207 17119
rect 37289 17085 37323 17119
rect 37473 17085 37507 17119
rect 39957 17085 39991 17119
rect 40141 17085 40175 17119
rect 40601 17085 40635 17119
rect 42533 17085 42567 17119
rect 42717 17085 42751 17119
rect 43177 17085 43211 17119
rect 45201 17085 45235 17119
rect 45385 17085 45419 17119
rect 12173 17017 12207 17051
rect 20085 16949 20119 16983
rect 47777 16949 47811 16983
rect 3065 16745 3099 16779
rect 5181 16745 5215 16779
rect 6561 16745 6595 16779
rect 7389 16745 7423 16779
rect 17969 16745 18003 16779
rect 22385 16745 22419 16779
rect 24501 16745 24535 16779
rect 28181 16745 28215 16779
rect 30021 16745 30055 16779
rect 30573 16745 30607 16779
rect 31677 16745 31711 16779
rect 37473 16745 37507 16779
rect 40509 16745 40543 16779
rect 42165 16745 42199 16779
rect 45109 16745 45143 16779
rect 9689 16609 9723 16643
rect 10149 16609 10183 16643
rect 10609 16609 10643 16643
rect 15117 16609 15151 16643
rect 15577 16609 15611 16643
rect 16129 16609 16163 16643
rect 19533 16609 19567 16643
rect 19993 16609 20027 16643
rect 20177 16609 20211 16643
rect 23857 16609 23891 16643
rect 32689 16609 32723 16643
rect 35449 16609 35483 16643
rect 42625 16609 42659 16643
rect 43821 16609 43855 16643
rect 45845 16609 45879 16643
rect 46305 16609 46339 16643
rect 2421 16541 2455 16575
rect 4537 16541 4571 16575
rect 7849 16541 7883 16575
rect 7941 16541 7975 16575
rect 12449 16541 12483 16575
rect 13553 16541 13587 16575
rect 18061 16541 18095 16575
rect 18521 16541 18555 16575
rect 22477 16541 22511 16575
rect 24409 16541 24443 16575
rect 25237 16541 25271 16575
rect 27077 16541 27111 16575
rect 27537 16541 27571 16575
rect 27629 16541 27663 16575
rect 28825 16541 28859 16575
rect 30113 16541 30147 16575
rect 31585 16541 31619 16575
rect 32229 16541 32263 16575
rect 36921 16541 36955 16575
rect 37381 16541 37415 16575
rect 38485 16541 38519 16575
rect 39129 16541 39163 16575
rect 39865 16541 39899 16575
rect 39957 16541 39991 16575
rect 45017 16541 45051 16575
rect 48145 16541 48179 16575
rect 2329 16473 2363 16507
rect 4445 16473 4479 16507
rect 10333 16473 10367 16507
rect 13461 16473 13495 16507
rect 15761 16473 15795 16507
rect 21833 16473 21867 16507
rect 26893 16473 26927 16507
rect 32413 16473 32447 16507
rect 36737 16473 36771 16507
rect 42809 16473 42843 16507
rect 46489 16473 46523 16507
rect 38577 16405 38611 16439
rect 7941 16201 7975 16235
rect 10333 16201 10367 16235
rect 15761 16201 15795 16235
rect 24593 16201 24627 16235
rect 32413 16201 32447 16235
rect 33885 16201 33919 16235
rect 35265 16201 35299 16235
rect 42625 16201 42659 16235
rect 43453 16201 43487 16235
rect 47685 16201 47719 16235
rect 30665 16133 30699 16167
rect 8033 16065 8067 16099
rect 10241 16065 10275 16099
rect 12357 16065 12391 16099
rect 15669 16065 15703 16099
rect 18245 16065 18279 16099
rect 24041 16065 24075 16099
rect 24501 16065 24535 16099
rect 25145 16065 25179 16099
rect 26249 16065 26283 16099
rect 26985 16065 27019 16099
rect 28825 16065 28859 16099
rect 31585 16065 31619 16099
rect 32505 16065 32539 16099
rect 33793 16065 33827 16099
rect 34621 16065 34655 16099
rect 35173 16065 35207 16099
rect 36645 16065 36679 16099
rect 37289 16065 37323 16099
rect 38945 16065 38979 16099
rect 40785 16065 40819 16099
rect 42533 16065 42567 16099
rect 43545 16065 43579 16099
rect 44741 16065 44775 16099
rect 47593 16065 47627 16099
rect 12541 15997 12575 16031
rect 12909 15997 12943 16031
rect 18429 15997 18463 16031
rect 18705 15997 18739 16031
rect 25329 15997 25363 16031
rect 29009 15997 29043 16031
rect 32965 15997 32999 16031
rect 39129 15997 39163 16031
rect 45201 15997 45235 16031
rect 45385 15997 45419 16031
rect 46857 15997 46891 16031
rect 2053 15861 2087 15895
rect 11713 15861 11747 15895
rect 16681 15861 16715 15895
rect 26157 15861 26191 15895
rect 35817 15861 35851 15895
rect 41245 15861 41279 15895
rect 18521 15657 18555 15691
rect 28457 15657 28491 15691
rect 43269 15657 43303 15691
rect 45293 15657 45327 15691
rect 11713 15521 11747 15555
rect 12449 15521 12483 15555
rect 16129 15521 16163 15555
rect 16773 15521 16807 15555
rect 25237 15521 25271 15555
rect 25421 15521 25455 15555
rect 25789 15521 25823 15555
rect 35633 15521 35667 15555
rect 36093 15521 36127 15555
rect 40877 15521 40911 15555
rect 41889 15521 41923 15555
rect 46765 15521 46799 15555
rect 48145 15521 48179 15555
rect 2513 15453 2547 15487
rect 15669 15453 15703 15487
rect 18613 15453 18647 15487
rect 19901 15453 19935 15487
rect 28365 15453 28399 15487
rect 40233 15453 40267 15487
rect 45201 15453 45235 15487
rect 11897 15385 11931 15419
rect 15577 15385 15611 15419
rect 16313 15385 16347 15419
rect 19441 15385 19475 15419
rect 24593 15385 24627 15419
rect 35817 15385 35851 15419
rect 40325 15385 40359 15419
rect 41061 15385 41095 15419
rect 47961 15385 47995 15419
rect 2421 15317 2455 15351
rect 24685 15317 24719 15351
rect 11897 15113 11931 15147
rect 12541 15113 12575 15147
rect 35909 15113 35943 15147
rect 47685 15113 47719 15147
rect 2237 15045 2271 15079
rect 25881 15045 25915 15079
rect 2053 14977 2087 15011
rect 11805 14977 11839 15011
rect 12449 14977 12483 15011
rect 18521 14977 18555 15011
rect 18981 14977 19015 15011
rect 20361 14977 20395 15011
rect 24685 14977 24719 15011
rect 25145 14977 25179 15011
rect 27077 14977 27111 15011
rect 27261 14977 27295 15011
rect 28181 14977 28215 15011
rect 28733 14977 28767 15011
rect 30941 14977 30975 15011
rect 32137 14977 32171 15011
rect 36001 14977 36035 15011
rect 45569 14977 45603 15011
rect 46857 14977 46891 15011
rect 47593 14977 47627 15011
rect 2789 14909 2823 14943
rect 18337 14909 18371 14943
rect 19717 14909 19751 14943
rect 20637 14909 20671 14943
rect 24501 14909 24535 14943
rect 29009 14909 29043 14943
rect 31401 14909 31435 14943
rect 32413 14909 32447 14943
rect 27905 14773 27939 14807
rect 46397 14773 46431 14807
rect 46949 14773 46983 14807
rect 18521 14569 18555 14603
rect 19625 14433 19659 14467
rect 46305 14433 46339 14467
rect 46489 14433 46523 14467
rect 48145 14433 48179 14467
rect 1961 14365 1995 14399
rect 2605 14365 2639 14399
rect 19901 14365 19935 14399
rect 25237 14365 25271 14399
rect 25697 14365 25731 14399
rect 26985 14365 27019 14399
rect 27261 14365 27295 14399
rect 31401 14365 31435 14399
rect 31677 14365 31711 14399
rect 45661 14365 45695 14399
rect 18613 14297 18647 14331
rect 27813 14297 27847 14331
rect 27997 14297 28031 14331
rect 2513 14229 2547 14263
rect 2237 13957 2271 13991
rect 28181 13957 28215 13991
rect 45385 13957 45419 13991
rect 47685 13957 47719 13991
rect 2053 13889 2087 13923
rect 25237 13889 25271 13923
rect 27353 13889 27387 13923
rect 28733 13889 28767 13923
rect 45201 13889 45235 13923
rect 47593 13889 47627 13923
rect 2789 13821 2823 13855
rect 25513 13821 25547 13855
rect 29009 13821 29043 13855
rect 46857 13821 46891 13855
rect 27169 13345 27203 13379
rect 45201 13345 45235 13379
rect 46305 13345 46339 13379
rect 2145 13277 2179 13311
rect 3801 13277 3835 13311
rect 26893 13277 26927 13311
rect 45661 13277 45695 13311
rect 45753 13209 45787 13243
rect 46489 13209 46523 13243
rect 48145 13209 48179 13243
rect 45385 12869 45419 12903
rect 47685 12869 47719 12903
rect 2053 12801 2087 12835
rect 27629 12801 27663 12835
rect 47593 12801 47627 12835
rect 2237 12733 2271 12767
rect 2789 12733 2823 12767
rect 27353 12733 27387 12767
rect 45201 12733 45235 12767
rect 46857 12733 46891 12767
rect 2513 12393 2547 12427
rect 44465 12393 44499 12427
rect 3801 12257 3835 12291
rect 4261 12257 4295 12291
rect 47593 12257 47627 12291
rect 2605 12189 2639 12223
rect 45477 12189 45511 12223
rect 45937 12189 45971 12223
rect 3985 12121 4019 12155
rect 46121 12121 46155 12155
rect 3893 11849 3927 11883
rect 47685 11849 47719 11883
rect 3985 11713 4019 11747
rect 47593 11713 47627 11747
rect 44741 11645 44775 11679
rect 45201 11645 45235 11679
rect 45385 11645 45419 11679
rect 46857 11645 46891 11679
rect 2145 11101 2179 11135
rect 45845 11101 45879 11135
rect 46305 11101 46339 11135
rect 46489 11033 46523 11067
rect 48145 11033 48179 11067
rect 46581 10761 46615 10795
rect 47685 10761 47719 10795
rect 2053 10625 2087 10659
rect 46673 10625 46707 10659
rect 47593 10625 47627 10659
rect 2237 10557 2271 10591
rect 2789 10557 2823 10591
rect 11529 10421 11563 10455
rect 13001 10421 13035 10455
rect 46029 10421 46063 10455
rect 2513 10217 2547 10251
rect 11069 10081 11103 10115
rect 11529 10081 11563 10115
rect 46305 10081 46339 10115
rect 48145 10081 48179 10115
rect 2605 10013 2639 10047
rect 13553 10013 13587 10047
rect 40049 10013 40083 10047
rect 11253 9945 11287 9979
rect 46489 9945 46523 9979
rect 13461 9877 13495 9911
rect 11621 9673 11655 9707
rect 13185 9605 13219 9639
rect 47685 9605 47719 9639
rect 11713 9537 11747 9571
rect 13001 9537 13035 9571
rect 40049 9537 40083 9571
rect 47593 9537 47627 9571
rect 13553 9469 13587 9503
rect 40233 9469 40267 9503
rect 40601 9469 40635 9503
rect 40141 9129 40175 9163
rect 2053 8925 2087 8959
rect 40049 8925 40083 8959
rect 2053 8449 2087 8483
rect 2237 8381 2271 8415
rect 2789 8381 2823 8415
rect 10425 8245 10459 8279
rect 2329 8041 2363 8075
rect 10333 7905 10367 7939
rect 10977 7905 11011 7939
rect 2421 7837 2455 7871
rect 17693 7837 17727 7871
rect 29837 7837 29871 7871
rect 33241 7837 33275 7871
rect 10517 7769 10551 7803
rect 33333 7701 33367 7735
rect 10517 7497 10551 7531
rect 33885 7429 33919 7463
rect 10425 7361 10459 7395
rect 17693 7361 17727 7395
rect 29101 7361 29135 7395
rect 29745 7361 29779 7395
rect 17877 7293 17911 7327
rect 18153 7293 18187 7327
rect 29193 7293 29227 7327
rect 29929 7293 29963 7327
rect 31585 7293 31619 7327
rect 33701 7293 33735 7327
rect 34621 7293 34655 7327
rect 2237 7157 2271 7191
rect 33701 6953 33735 6987
rect 18245 6817 18279 6851
rect 2697 6749 2731 6783
rect 18337 6749 18371 6783
rect 46765 6749 46799 6783
rect 47685 6749 47719 6783
rect 2605 6613 2639 6647
rect 2329 6341 2363 6375
rect 2145 6273 2179 6307
rect 47593 6273 47627 6307
rect 2789 6205 2823 6239
rect 45201 6205 45235 6239
rect 45385 6205 45419 6239
rect 46581 6205 46615 6239
rect 47685 6069 47719 6103
rect 45201 5865 45235 5899
rect 46673 5729 46707 5763
rect 48145 5729 48179 5763
rect 1961 5661 1995 5695
rect 2605 5661 2639 5695
rect 3249 5661 3283 5695
rect 5733 5661 5767 5695
rect 45661 5661 45695 5695
rect 47961 5593 47995 5627
rect 2513 5525 2547 5559
rect 47685 5321 47719 5355
rect 2329 5253 2363 5287
rect 2145 5185 2179 5219
rect 5641 5185 5675 5219
rect 6929 5185 6963 5219
rect 27997 5185 28031 5219
rect 45201 5185 45235 5219
rect 47593 5185 47627 5219
rect 2789 5117 2823 5151
rect 45385 5117 45419 5151
rect 46857 5117 46891 5151
rect 1501 4981 1535 5015
rect 5549 4981 5583 5015
rect 6837 4981 6871 5015
rect 28089 4981 28123 5015
rect 33057 4981 33091 5015
rect 44097 4981 44131 5015
rect 44741 4981 44775 5015
rect 45293 4777 45327 4811
rect 1409 4641 1443 4675
rect 3249 4641 3283 4675
rect 5181 4641 5215 4675
rect 5549 4641 5583 4675
rect 46305 4641 46339 4675
rect 3985 4573 4019 4607
rect 4997 4573 5031 4607
rect 8953 4573 8987 4607
rect 15761 4573 15795 4607
rect 27905 4573 27939 4607
rect 28733 4573 28767 4607
rect 32045 4573 32079 4607
rect 33057 4573 33091 4607
rect 34161 4573 34195 4607
rect 34713 4573 34747 4607
rect 35909 4573 35943 4607
rect 37197 4573 37231 4607
rect 42349 4573 42383 4607
rect 43269 4573 43303 4607
rect 43729 4573 43763 4607
rect 45201 4573 45235 4607
rect 3065 4505 3099 4539
rect 3893 4505 3927 4539
rect 7849 4505 7883 4539
rect 8217 4505 8251 4539
rect 46489 4505 46523 4539
rect 48145 4505 48179 4539
rect 33149 4437 33183 4471
rect 34805 4437 34839 4471
rect 42441 4437 42475 4471
rect 43177 4437 43211 4471
rect 6561 4165 6595 4199
rect 28089 4165 28123 4199
rect 33149 4165 33183 4199
rect 2237 4097 2271 4131
rect 4997 4097 5031 4131
rect 9229 4097 9263 4131
rect 15853 4097 15887 4131
rect 26985 4097 27019 4131
rect 27905 4097 27939 4131
rect 32137 4097 32171 4131
rect 32965 4097 32999 4131
rect 35909 4097 35943 4131
rect 36553 4097 36587 4131
rect 37289 4097 37323 4131
rect 44741 4097 44775 4131
rect 47593 4097 47627 4131
rect 2881 4029 2915 4063
rect 4353 4029 4387 4063
rect 4537 4029 4571 4063
rect 6377 4029 6411 4063
rect 6837 4029 6871 4063
rect 18705 4029 18739 4063
rect 19901 4029 19935 4063
rect 20085 4029 20119 4063
rect 27261 4029 27295 4063
rect 28365 4029 28399 4063
rect 33517 4029 33551 4063
rect 36645 4029 36679 4063
rect 37473 4029 37507 4063
rect 37749 4029 37783 4063
rect 42441 4029 42475 4063
rect 42625 4029 42659 4063
rect 44281 4029 44315 4063
rect 44925 4029 44959 4063
rect 46581 4029 46615 4063
rect 13829 3961 13863 3995
rect 2145 3893 2179 3927
rect 5825 3893 5859 3927
rect 9321 3893 9355 3927
rect 9873 3893 9907 3927
rect 11713 3893 11747 3927
rect 12541 3893 12575 3927
rect 14289 3893 14323 3927
rect 15945 3893 15979 3927
rect 31585 3893 31619 3927
rect 32229 3893 32263 3927
rect 35265 3893 35299 3927
rect 36001 3893 36035 3927
rect 39957 3893 39991 3927
rect 41889 3893 41923 3927
rect 47685 3893 47719 3927
rect 3893 3689 3927 3723
rect 4445 3689 4479 3723
rect 5273 3689 5307 3723
rect 19349 3689 19383 3723
rect 20085 3689 20119 3723
rect 45109 3689 45143 3723
rect 1409 3553 1443 3587
rect 1593 3553 1627 3587
rect 2789 3553 2823 3587
rect 5733 3553 5767 3587
rect 6193 3553 6227 3587
rect 9137 3553 9171 3587
rect 9321 3553 9355 3587
rect 9689 3553 9723 3587
rect 11621 3553 11655 3587
rect 12265 3553 12299 3587
rect 15761 3553 15795 3587
rect 15945 3553 15979 3587
rect 16221 3553 16255 3587
rect 27721 3553 27755 3587
rect 32045 3553 32079 3587
rect 32229 3553 32263 3587
rect 32689 3553 32723 3587
rect 35909 3553 35943 3587
rect 36093 3553 36127 3587
rect 36737 3553 36771 3587
rect 41981 3553 42015 3587
rect 46489 3553 46523 3587
rect 3985 3485 4019 3519
rect 8217 3485 8251 3519
rect 14289 3485 14323 3519
rect 15117 3485 15151 3519
rect 18153 3485 18187 3519
rect 19257 3485 19291 3519
rect 23857 3485 23891 3519
rect 24869 3485 24903 3519
rect 25513 3485 25547 3519
rect 26433 3485 26467 3519
rect 26893 3485 26927 3519
rect 29561 3485 29595 3519
rect 31309 3485 31343 3519
rect 34713 3485 34747 3519
rect 38209 3485 38243 3519
rect 39129 3485 39163 3519
rect 39865 3485 39899 3519
rect 42441 3485 42475 3519
rect 45201 3485 45235 3519
rect 45845 3485 45879 3519
rect 46305 3485 46339 3519
rect 5917 3417 5951 3451
rect 11805 3417 11839 3451
rect 27077 3417 27111 3451
rect 41714 3417 41748 3451
rect 42625 3417 42659 3451
rect 44281 3417 44315 3451
rect 48145 3417 48179 3451
rect 8309 3349 8343 3383
rect 14381 3349 14415 3383
rect 15025 3349 15059 3383
rect 18245 3349 18279 3383
rect 24777 3349 24811 3383
rect 25421 3349 25455 3383
rect 34805 3349 34839 3383
rect 39957 3349 39991 3383
rect 40601 3349 40635 3383
rect 5733 3145 5767 3179
rect 11805 3145 11839 3179
rect 27077 3145 27111 3179
rect 41705 3145 41739 3179
rect 46673 3145 46707 3179
rect 8309 3077 8343 3111
rect 9045 3077 9079 3111
rect 15301 3077 15335 3111
rect 18337 3077 18371 3111
rect 24133 3077 24167 3111
rect 25789 3077 25823 3111
rect 28273 3077 28307 3111
rect 29009 3077 29043 3111
rect 31493 3077 31527 3111
rect 32321 3077 32355 3111
rect 35081 3077 35115 3111
rect 42625 3077 42659 3111
rect 43361 3077 43395 3111
rect 4629 3009 4663 3043
rect 5825 3009 5859 3043
rect 6929 3009 6963 3043
rect 8217 3009 8251 3043
rect 11713 3009 11747 3043
rect 12633 3009 12667 3043
rect 15485 3009 15519 3043
rect 15945 3009 15979 3043
rect 20453 3009 20487 3043
rect 22569 3009 22603 3043
rect 23949 3009 23983 3043
rect 26985 3009 27019 3043
rect 28181 3009 28215 3043
rect 28825 3009 28859 3043
rect 31401 3009 31435 3043
rect 32137 3009 32171 3043
rect 34897 3009 34931 3043
rect 37289 3009 37323 3043
rect 38485 3009 38519 3043
rect 39129 3009 39163 3043
rect 41889 3009 41923 3043
rect 42533 3009 42567 3043
rect 45477 3009 45511 3043
rect 46765 3009 46799 3043
rect 47593 3009 47627 3043
rect 1685 2941 1719 2975
rect 2145 2941 2179 2975
rect 2329 2941 2363 2975
rect 2605 2941 2639 2975
rect 7757 2941 7791 2975
rect 8861 2941 8895 2975
rect 9321 2941 9355 2975
rect 13829 2941 13863 2975
rect 17693 2941 17727 2975
rect 18153 2941 18187 2975
rect 19349 2941 19383 2975
rect 29653 2941 29687 2975
rect 33977 2941 34011 2975
rect 36093 2941 36127 2975
rect 38577 2941 38611 2975
rect 39313 2941 39347 2975
rect 40969 2941 41003 2975
rect 43177 2941 43211 2975
rect 43913 2941 43947 2975
rect 22477 2873 22511 2907
rect 4537 2805 4571 2839
rect 6837 2805 6871 2839
rect 12541 2805 12575 2839
rect 16037 2805 16071 2839
rect 16681 2805 16715 2839
rect 20545 2805 20579 2839
rect 21281 2805 21315 2839
rect 23213 2805 23247 2839
rect 26433 2805 26467 2839
rect 37381 2805 37415 2839
rect 45569 2805 45603 2839
rect 47685 2805 47719 2839
rect 2513 2601 2547 2635
rect 3985 2465 4019 2499
rect 4629 2465 4663 2499
rect 6377 2465 6411 2499
rect 6561 2465 6595 2499
rect 6837 2465 6871 2499
rect 8953 2465 8987 2499
rect 9413 2465 9447 2499
rect 11713 2465 11747 2499
rect 13369 2465 13403 2499
rect 13553 2465 13587 2499
rect 14197 2465 14231 2499
rect 14381 2465 14415 2499
rect 14841 2465 14875 2499
rect 16681 2465 16715 2499
rect 17141 2465 17175 2499
rect 20821 2465 20855 2499
rect 21097 2465 21131 2499
rect 21281 2465 21315 2499
rect 22477 2465 22511 2499
rect 23673 2465 23707 2499
rect 23857 2465 23891 2499
rect 26249 2465 26283 2499
rect 26433 2465 26467 2499
rect 28549 2465 28583 2499
rect 29009 2465 29043 2499
rect 32137 2465 32171 2499
rect 32597 2465 32631 2499
rect 34713 2465 34747 2499
rect 34897 2465 34931 2499
rect 37289 2465 37323 2499
rect 37473 2465 37507 2499
rect 39957 2465 39991 2499
rect 40141 2465 40175 2499
rect 43729 2465 43763 2499
rect 46581 2465 46615 2499
rect 46857 2465 46891 2499
rect 2605 2397 2639 2431
rect 3249 2397 3283 2431
rect 3801 2397 3835 2431
rect 29561 2397 29595 2431
rect 31125 2397 31159 2431
rect 44465 2397 44499 2431
rect 47041 2397 47075 2431
rect 47593 2397 47627 2431
rect 9137 2329 9171 2363
rect 16865 2329 16899 2363
rect 24593 2329 24627 2363
rect 28825 2329 28859 2363
rect 29653 2329 29687 2363
rect 31217 2329 31251 2363
rect 32321 2329 32355 2363
rect 36553 2329 36587 2363
rect 39129 2329 39163 2363
rect 41797 2329 41831 2363
rect 44281 2329 44315 2363
<< metal1 >>
rect 4614 17484 4620 17536
rect 4672 17524 4678 17536
rect 12342 17524 12348 17536
rect 4672 17496 12348 17524
rect 4672 17484 4678 17496
rect 12342 17484 12348 17496
rect 12400 17484 12406 17536
rect 1104 17434 48852 17456
rect 1104 17382 16880 17434
rect 16932 17382 16944 17434
rect 16996 17382 17008 17434
rect 17060 17382 17072 17434
rect 17124 17382 17136 17434
rect 17188 17382 32811 17434
rect 32863 17382 32875 17434
rect 32927 17382 32939 17434
rect 32991 17382 33003 17434
rect 33055 17382 33067 17434
rect 33119 17382 48852 17434
rect 1104 17360 48852 17382
rect 4062 17280 4068 17332
rect 4120 17320 4126 17332
rect 4120 17292 15516 17320
rect 4120 17280 4126 17292
rect 1394 17252 1400 17264
rect 1355 17224 1400 17252
rect 1394 17212 1400 17224
rect 1452 17212 1458 17264
rect 2590 17212 2596 17264
rect 2648 17252 2654 17264
rect 3973 17255 4031 17261
rect 3973 17252 3985 17255
rect 2648 17224 3985 17252
rect 2648 17212 2654 17224
rect 3973 17221 3985 17224
rect 4019 17221 4031 17255
rect 3973 17215 4031 17221
rect 8294 17212 8300 17264
rect 8352 17252 8358 17264
rect 9125 17255 9183 17261
rect 9125 17252 9137 17255
rect 8352 17224 9137 17252
rect 8352 17212 8358 17224
rect 9125 17221 9137 17224
rect 9171 17221 9183 17255
rect 9125 17215 9183 17221
rect 11606 17212 11612 17264
rect 11664 17252 11670 17264
rect 11977 17255 12035 17261
rect 11977 17252 11989 17255
rect 11664 17224 11989 17252
rect 11664 17212 11670 17224
rect 11977 17221 11989 17224
rect 12023 17221 12035 17255
rect 11977 17215 12035 17221
rect 3050 17116 3056 17128
rect 3011 17088 3056 17116
rect 3050 17076 3056 17088
rect 3108 17076 3114 17128
rect 3234 17116 3240 17128
rect 3195 17088 3240 17116
rect 3234 17076 3240 17088
rect 3292 17076 3298 17128
rect 5626 17116 5632 17128
rect 5587 17088 5632 17116
rect 5626 17076 5632 17088
rect 5684 17076 5690 17128
rect 5810 17116 5816 17128
rect 5771 17088 5816 17116
rect 5810 17076 5816 17088
rect 5868 17076 5874 17128
rect 6546 17116 6552 17128
rect 6507 17088 6552 17116
rect 6546 17076 6552 17088
rect 6604 17076 6610 17128
rect 6733 17119 6791 17125
rect 6733 17085 6745 17119
rect 6779 17116 6791 17119
rect 7558 17116 7564 17128
rect 6779 17088 7564 17116
rect 6779 17085 6791 17088
rect 6733 17079 6791 17085
rect 7558 17076 7564 17088
rect 7616 17076 7622 17128
rect 7742 17116 7748 17128
rect 7703 17088 7748 17116
rect 7742 17076 7748 17088
rect 7800 17076 7806 17128
rect 7926 17076 7932 17128
rect 7984 17116 7990 17128
rect 8941 17119 8999 17125
rect 8941 17116 8953 17119
rect 7984 17088 8953 17116
rect 7984 17076 7990 17088
rect 8941 17085 8953 17088
rect 8987 17085 8999 17119
rect 8941 17079 8999 17085
rect 9401 17119 9459 17125
rect 9401 17085 9413 17119
rect 9447 17085 9459 17119
rect 9401 17079 9459 17085
rect 12989 17119 13047 17125
rect 12989 17085 13001 17119
rect 13035 17116 13047 17119
rect 14093 17119 14151 17125
rect 14093 17116 14105 17119
rect 13035 17088 14105 17116
rect 13035 17085 13047 17088
rect 12989 17079 13047 17085
rect 14093 17085 14105 17088
rect 14139 17085 14151 17119
rect 14274 17116 14280 17128
rect 14235 17088 14280 17116
rect 14093 17079 14151 17085
rect 8386 17008 8392 17060
rect 8444 17048 8450 17060
rect 9416 17048 9444 17079
rect 14274 17076 14280 17088
rect 14332 17076 14338 17128
rect 15488 17125 15516 17292
rect 18138 17280 18144 17332
rect 18196 17320 18202 17332
rect 24486 17320 24492 17332
rect 18196 17292 24492 17320
rect 18196 17280 18202 17292
rect 24486 17280 24492 17292
rect 24544 17280 24550 17332
rect 15562 17212 15568 17264
rect 15620 17252 15626 17264
rect 23842 17252 23848 17264
rect 15620 17224 20024 17252
rect 23803 17224 23848 17252
rect 15620 17212 15626 17224
rect 19996 17193 20024 17224
rect 23842 17212 23848 17224
rect 23900 17212 23906 17264
rect 31386 17252 31392 17264
rect 28920 17224 31392 17252
rect 19981 17187 20039 17193
rect 19981 17153 19993 17187
rect 20027 17153 20039 17187
rect 19981 17147 20039 17153
rect 15473 17119 15531 17125
rect 15473 17085 15485 17119
rect 15519 17085 15531 17119
rect 15473 17079 15531 17085
rect 17865 17119 17923 17125
rect 17865 17085 17877 17119
rect 17911 17116 17923 17119
rect 18046 17116 18052 17128
rect 17911 17088 18052 17116
rect 17911 17085 17923 17088
rect 17865 17079 17923 17085
rect 18046 17076 18052 17088
rect 18104 17076 18110 17128
rect 18506 17116 18512 17128
rect 18467 17088 18512 17116
rect 18506 17076 18512 17088
rect 18564 17076 18570 17128
rect 18693 17119 18751 17125
rect 18693 17085 18705 17119
rect 18739 17116 18751 17119
rect 19245 17119 19303 17125
rect 19245 17116 19257 17119
rect 18739 17088 19257 17116
rect 18739 17085 18751 17088
rect 18693 17079 18751 17085
rect 19245 17085 19257 17088
rect 19291 17085 19303 17119
rect 19245 17079 19303 17085
rect 12158 17048 12164 17060
rect 8444 17020 9444 17048
rect 12119 17020 12164 17048
rect 8444 17008 8450 17020
rect 12158 17008 12164 17020
rect 12216 17008 12222 17060
rect 12342 17008 12348 17060
rect 12400 17048 12406 17060
rect 19886 17048 19892 17060
rect 12400 17020 19892 17048
rect 12400 17008 12406 17020
rect 19886 17008 19892 17020
rect 19944 17008 19950 17060
rect 19996 17048 20024 17147
rect 21269 17119 21327 17125
rect 21269 17085 21281 17119
rect 21315 17116 21327 17119
rect 22005 17119 22063 17125
rect 22005 17116 22017 17119
rect 21315 17088 22017 17116
rect 21315 17085 21327 17088
rect 21269 17079 21327 17085
rect 22005 17085 22017 17088
rect 22051 17085 22063 17119
rect 22186 17116 22192 17128
rect 22147 17088 22192 17116
rect 22005 17079 22063 17085
rect 22186 17076 22192 17088
rect 22244 17076 22250 17128
rect 24394 17116 24400 17128
rect 24355 17088 24400 17116
rect 24394 17076 24400 17088
rect 24452 17076 24458 17128
rect 24578 17116 24584 17128
rect 24539 17088 24584 17116
rect 24578 17076 24584 17088
rect 24636 17076 24642 17128
rect 24854 17116 24860 17128
rect 24815 17088 24860 17116
rect 24854 17076 24860 17088
rect 24912 17076 24918 17128
rect 27154 17116 27160 17128
rect 27115 17088 27160 17116
rect 27154 17076 27160 17088
rect 27212 17076 27218 17128
rect 27341 17119 27399 17125
rect 27341 17085 27353 17119
rect 27387 17116 27399 17119
rect 27614 17116 27620 17128
rect 27387 17088 27620 17116
rect 27387 17085 27399 17088
rect 27341 17079 27399 17085
rect 27614 17076 27620 17088
rect 27672 17076 27678 17128
rect 28920 17048 28948 17224
rect 31386 17212 31392 17224
rect 31444 17212 31450 17264
rect 39117 17255 39175 17261
rect 39117 17221 39129 17255
rect 39163 17252 39175 17255
rect 39942 17252 39948 17264
rect 39163 17224 39948 17252
rect 39163 17221 39175 17224
rect 39117 17215 39175 17221
rect 39942 17212 39948 17224
rect 40000 17212 40006 17264
rect 47026 17252 47032 17264
rect 46987 17224 47032 17252
rect 47026 17212 47032 17224
rect 47084 17212 47090 17264
rect 28997 17119 29055 17125
rect 28997 17085 29009 17119
rect 29043 17085 29055 17119
rect 28997 17079 29055 17085
rect 29733 17119 29791 17125
rect 29733 17085 29745 17119
rect 29779 17085 29791 17119
rect 29914 17116 29920 17128
rect 29875 17088 29920 17116
rect 29733 17079 29791 17085
rect 19996 17020 28948 17048
rect 7742 16940 7748 16992
rect 7800 16980 7806 16992
rect 15654 16980 15660 16992
rect 7800 16952 15660 16980
rect 7800 16940 7806 16952
rect 15654 16940 15660 16952
rect 15712 16940 15718 16992
rect 17126 16940 17132 16992
rect 17184 16980 17190 16992
rect 19702 16980 19708 16992
rect 17184 16952 19708 16980
rect 17184 16940 17190 16952
rect 19702 16940 19708 16952
rect 19760 16940 19766 16992
rect 20073 16983 20131 16989
rect 20073 16949 20085 16983
rect 20119 16980 20131 16983
rect 20162 16980 20168 16992
rect 20119 16952 20168 16980
rect 20119 16949 20131 16952
rect 20073 16943 20131 16949
rect 20162 16940 20168 16952
rect 20220 16940 20226 16992
rect 29012 16980 29040 17079
rect 29748 17048 29776 17079
rect 29914 17076 29920 17088
rect 29972 17076 29978 17128
rect 30926 17116 30932 17128
rect 30887 17088 30932 17116
rect 30926 17076 30932 17088
rect 30984 17076 30990 17128
rect 32122 17116 32128 17128
rect 32083 17088 32128 17116
rect 32122 17076 32128 17088
rect 32180 17076 32186 17128
rect 32306 17116 32312 17128
rect 32267 17088 32312 17116
rect 32306 17076 32312 17088
rect 32364 17076 32370 17128
rect 32398 17076 32404 17128
rect 32456 17116 32462 17128
rect 32585 17119 32643 17125
rect 32585 17116 32597 17119
rect 32456 17088 32597 17116
rect 32456 17076 32462 17088
rect 32585 17085 32597 17088
rect 32631 17085 32643 17119
rect 34698 17116 34704 17128
rect 34659 17088 34704 17116
rect 32585 17079 32643 17085
rect 34698 17076 34704 17088
rect 34756 17076 34762 17128
rect 34882 17116 34888 17128
rect 34843 17088 34888 17116
rect 34882 17076 34888 17088
rect 34940 17076 34946 17128
rect 35161 17119 35219 17125
rect 35161 17085 35173 17119
rect 35207 17085 35219 17119
rect 37274 17116 37280 17128
rect 37235 17088 37280 17116
rect 35161 17079 35219 17085
rect 30558 17048 30564 17060
rect 29748 17020 30564 17048
rect 30558 17008 30564 17020
rect 30616 17008 30622 17060
rect 33502 17008 33508 17060
rect 33560 17048 33566 17060
rect 35176 17048 35204 17079
rect 37274 17076 37280 17088
rect 37332 17076 37338 17128
rect 37458 17116 37464 17128
rect 37419 17088 37464 17116
rect 37458 17076 37464 17088
rect 37516 17076 37522 17128
rect 39942 17116 39948 17128
rect 39903 17088 39948 17116
rect 39942 17076 39948 17088
rect 40000 17076 40006 17128
rect 40126 17116 40132 17128
rect 40087 17088 40132 17116
rect 40126 17076 40132 17088
rect 40184 17076 40190 17128
rect 40586 17116 40592 17128
rect 40547 17088 40592 17116
rect 40586 17076 40592 17088
rect 40644 17076 40650 17128
rect 42150 17076 42156 17128
rect 42208 17116 42214 17128
rect 42521 17119 42579 17125
rect 42521 17116 42533 17119
rect 42208 17088 42533 17116
rect 42208 17076 42214 17088
rect 42521 17085 42533 17088
rect 42567 17085 42579 17119
rect 42702 17116 42708 17128
rect 42663 17088 42708 17116
rect 42521 17079 42579 17085
rect 42702 17076 42708 17088
rect 42760 17076 42766 17128
rect 43162 17116 43168 17128
rect 43123 17088 43168 17116
rect 43162 17076 43168 17088
rect 43220 17076 43226 17128
rect 44726 17076 44732 17128
rect 44784 17116 44790 17128
rect 45189 17119 45247 17125
rect 45189 17116 45201 17119
rect 44784 17088 45201 17116
rect 44784 17076 44790 17088
rect 45189 17085 45201 17088
rect 45235 17085 45247 17119
rect 45370 17116 45376 17128
rect 45331 17088 45376 17116
rect 45189 17079 45247 17085
rect 45370 17076 45376 17088
rect 45428 17076 45434 17128
rect 33560 17020 35204 17048
rect 33560 17008 33566 17020
rect 38010 16980 38016 16992
rect 29012 16952 38016 16980
rect 38010 16940 38016 16952
rect 38068 16940 38074 16992
rect 40678 16940 40684 16992
rect 40736 16980 40742 16992
rect 47486 16980 47492 16992
rect 40736 16952 47492 16980
rect 40736 16940 40742 16952
rect 47486 16940 47492 16952
rect 47544 16940 47550 16992
rect 47762 16980 47768 16992
rect 47723 16952 47768 16980
rect 47762 16940 47768 16952
rect 47820 16940 47826 16992
rect 1104 16890 48852 16912
rect 1104 16838 8915 16890
rect 8967 16838 8979 16890
rect 9031 16838 9043 16890
rect 9095 16838 9107 16890
rect 9159 16838 9171 16890
rect 9223 16838 24846 16890
rect 24898 16838 24910 16890
rect 24962 16838 24974 16890
rect 25026 16838 25038 16890
rect 25090 16838 25102 16890
rect 25154 16838 40776 16890
rect 40828 16838 40840 16890
rect 40892 16838 40904 16890
rect 40956 16838 40968 16890
rect 41020 16838 41032 16890
rect 41084 16838 48852 16890
rect 1104 16816 48852 16838
rect 3053 16779 3111 16785
rect 3053 16745 3065 16779
rect 3099 16776 3111 16779
rect 3234 16776 3240 16788
rect 3099 16748 3240 16776
rect 3099 16745 3111 16748
rect 3053 16739 3111 16745
rect 3234 16736 3240 16748
rect 3292 16736 3298 16788
rect 5169 16779 5227 16785
rect 5169 16745 5181 16779
rect 5215 16776 5227 16779
rect 5810 16776 5816 16788
rect 5215 16748 5816 16776
rect 5215 16745 5227 16748
rect 5169 16739 5227 16745
rect 5810 16736 5816 16748
rect 5868 16736 5874 16788
rect 6546 16776 6552 16788
rect 6507 16748 6552 16776
rect 6546 16736 6552 16748
rect 6604 16736 6610 16788
rect 7377 16779 7435 16785
rect 7377 16745 7389 16779
rect 7423 16776 7435 16779
rect 7926 16776 7932 16788
rect 7423 16748 7932 16776
rect 7423 16745 7435 16748
rect 7377 16739 7435 16745
rect 7926 16736 7932 16748
rect 7984 16736 7990 16788
rect 15562 16776 15568 16788
rect 12406 16748 15568 16776
rect 12406 16708 12434 16748
rect 15562 16736 15568 16748
rect 15620 16736 15626 16788
rect 15654 16736 15660 16788
rect 15712 16776 15718 16788
rect 17957 16779 18015 16785
rect 15712 16748 17264 16776
rect 15712 16736 15718 16748
rect 17126 16708 17132 16720
rect 2424 16680 12434 16708
rect 13556 16680 17132 16708
rect 2424 16584 2452 16680
rect 4614 16600 4620 16652
rect 4672 16600 4678 16652
rect 7742 16600 7748 16652
rect 7800 16640 7806 16652
rect 9677 16643 9735 16649
rect 7800 16612 7880 16640
rect 7800 16600 7806 16612
rect 2406 16572 2412 16584
rect 2367 16544 2412 16572
rect 2406 16532 2412 16544
rect 2464 16532 2470 16584
rect 4525 16575 4583 16581
rect 4525 16541 4537 16575
rect 4571 16572 4583 16575
rect 4632 16572 4660 16600
rect 7852 16581 7880 16612
rect 9677 16609 9689 16643
rect 9723 16640 9735 16643
rect 10137 16643 10195 16649
rect 10137 16640 10149 16643
rect 9723 16612 10149 16640
rect 9723 16609 9735 16612
rect 9677 16603 9735 16609
rect 10137 16609 10149 16612
rect 10183 16609 10195 16643
rect 10594 16640 10600 16652
rect 10555 16612 10600 16640
rect 10137 16603 10195 16609
rect 10594 16600 10600 16612
rect 10652 16600 10658 16652
rect 4571 16544 4660 16572
rect 7837 16575 7895 16581
rect 4571 16541 4583 16544
rect 4525 16535 4583 16541
rect 7837 16541 7849 16575
rect 7883 16541 7895 16575
rect 7837 16535 7895 16541
rect 7929 16575 7987 16581
rect 7929 16541 7941 16575
rect 7975 16572 7987 16575
rect 8294 16572 8300 16584
rect 7975 16544 8300 16572
rect 7975 16541 7987 16544
rect 7929 16535 7987 16541
rect 8294 16532 8300 16544
rect 8352 16532 8358 16584
rect 12434 16572 12440 16584
rect 12395 16544 12440 16572
rect 12434 16532 12440 16544
rect 12492 16532 12498 16584
rect 13556 16581 13584 16680
rect 17126 16668 17132 16680
rect 17184 16668 17190 16720
rect 17236 16708 17264 16748
rect 17957 16745 17969 16779
rect 18003 16776 18015 16779
rect 18506 16776 18512 16788
rect 18003 16748 18512 16776
rect 18003 16745 18015 16748
rect 17957 16739 18015 16745
rect 18506 16736 18512 16748
rect 18564 16736 18570 16788
rect 22186 16736 22192 16788
rect 22244 16776 22250 16788
rect 22373 16779 22431 16785
rect 22373 16776 22385 16779
rect 22244 16748 22385 16776
rect 22244 16736 22250 16748
rect 22373 16745 22385 16748
rect 22419 16745 22431 16779
rect 22373 16739 22431 16745
rect 24489 16779 24547 16785
rect 24489 16745 24501 16779
rect 24535 16776 24547 16779
rect 24578 16776 24584 16788
rect 24535 16748 24584 16776
rect 24535 16745 24547 16748
rect 24489 16739 24547 16745
rect 24578 16736 24584 16748
rect 24636 16736 24642 16788
rect 24670 16736 24676 16788
rect 24728 16776 24734 16788
rect 26786 16776 26792 16788
rect 24728 16748 26792 16776
rect 24728 16736 24734 16748
rect 26786 16736 26792 16748
rect 26844 16736 26850 16788
rect 27154 16736 27160 16788
rect 27212 16776 27218 16788
rect 28169 16779 28227 16785
rect 28169 16776 28181 16779
rect 27212 16748 28181 16776
rect 27212 16736 27218 16748
rect 28169 16745 28181 16748
rect 28215 16745 28227 16779
rect 28169 16739 28227 16745
rect 29914 16736 29920 16788
rect 29972 16776 29978 16788
rect 30009 16779 30067 16785
rect 30009 16776 30021 16779
rect 29972 16748 30021 16776
rect 29972 16736 29978 16748
rect 30009 16745 30021 16748
rect 30055 16745 30067 16779
rect 30558 16776 30564 16788
rect 30519 16748 30564 16776
rect 30009 16739 30067 16745
rect 30558 16736 30564 16748
rect 30616 16736 30622 16788
rect 31665 16779 31723 16785
rect 31665 16745 31677 16779
rect 31711 16776 31723 16779
rect 32306 16776 32312 16788
rect 31711 16748 32312 16776
rect 31711 16745 31723 16748
rect 31665 16739 31723 16745
rect 32306 16736 32312 16748
rect 32364 16736 32370 16788
rect 37458 16776 37464 16788
rect 37419 16748 37464 16776
rect 37458 16736 37464 16748
rect 37516 16736 37522 16788
rect 39942 16736 39948 16788
rect 40000 16776 40006 16788
rect 40497 16779 40555 16785
rect 40497 16776 40509 16779
rect 40000 16748 40509 16776
rect 40000 16736 40006 16748
rect 40497 16745 40509 16748
rect 40543 16745 40555 16779
rect 42150 16776 42156 16788
rect 42111 16748 42156 16776
rect 40497 16739 40555 16745
rect 42150 16736 42156 16748
rect 42208 16736 42214 16788
rect 45097 16779 45155 16785
rect 45097 16745 45109 16779
rect 45143 16776 45155 16779
rect 45370 16776 45376 16788
rect 45143 16748 45376 16776
rect 45143 16745 45155 16748
rect 45097 16739 45155 16745
rect 45370 16736 45376 16748
rect 45428 16736 45434 16788
rect 17236 16680 18000 16708
rect 17972 16652 18000 16680
rect 19886 16668 19892 16720
rect 19944 16708 19950 16720
rect 27890 16708 27896 16720
rect 19944 16680 22048 16708
rect 19944 16668 19950 16680
rect 15105 16643 15163 16649
rect 15105 16609 15117 16643
rect 15151 16640 15163 16643
rect 15565 16643 15623 16649
rect 15565 16640 15577 16643
rect 15151 16612 15577 16640
rect 15151 16609 15163 16612
rect 15105 16603 15163 16609
rect 15565 16609 15577 16612
rect 15611 16609 15623 16643
rect 16114 16640 16120 16652
rect 16075 16612 16120 16640
rect 15565 16603 15623 16609
rect 16114 16600 16120 16612
rect 16172 16600 16178 16652
rect 17954 16600 17960 16652
rect 18012 16600 18018 16652
rect 19521 16643 19579 16649
rect 19521 16609 19533 16643
rect 19567 16640 19579 16643
rect 19981 16643 20039 16649
rect 19981 16640 19993 16643
rect 19567 16612 19993 16640
rect 19567 16609 19579 16612
rect 19521 16603 19579 16609
rect 19981 16609 19993 16612
rect 20027 16609 20039 16643
rect 20162 16640 20168 16652
rect 20123 16612 20168 16640
rect 19981 16603 20039 16609
rect 20162 16600 20168 16612
rect 20220 16600 20226 16652
rect 22020 16640 22048 16680
rect 22480 16680 27896 16708
rect 22480 16640 22508 16680
rect 27890 16668 27896 16680
rect 27948 16668 27954 16720
rect 40678 16708 40684 16720
rect 30116 16680 40684 16708
rect 22020 16612 22508 16640
rect 13541 16575 13599 16581
rect 13541 16541 13553 16575
rect 13587 16541 13599 16575
rect 13541 16535 13599 16541
rect 18049 16575 18107 16581
rect 18049 16541 18061 16575
rect 18095 16572 18107 16575
rect 18138 16572 18144 16584
rect 18095 16544 18144 16572
rect 18095 16541 18107 16544
rect 18049 16535 18107 16541
rect 18138 16532 18144 16544
rect 18196 16532 18202 16584
rect 18230 16532 18236 16584
rect 18288 16572 18294 16584
rect 22480 16581 22508 16612
rect 23845 16643 23903 16649
rect 23845 16609 23857 16643
rect 23891 16640 23903 16643
rect 25130 16640 25136 16652
rect 23891 16612 25136 16640
rect 23891 16609 23903 16612
rect 23845 16603 23903 16609
rect 25130 16600 25136 16612
rect 25188 16600 25194 16652
rect 30006 16600 30012 16652
rect 30064 16640 30070 16652
rect 30116 16640 30144 16680
rect 40678 16668 40684 16680
rect 40736 16668 40742 16720
rect 42426 16668 42432 16720
rect 42484 16708 42490 16720
rect 46566 16708 46572 16720
rect 42484 16680 46572 16708
rect 42484 16668 42490 16680
rect 46566 16668 46572 16680
rect 46624 16668 46630 16720
rect 30064 16612 30144 16640
rect 30064 16600 30070 16612
rect 18509 16575 18567 16581
rect 18509 16572 18521 16575
rect 18288 16544 18521 16572
rect 18288 16532 18294 16544
rect 18509 16541 18521 16544
rect 18555 16541 18567 16575
rect 18509 16535 18567 16541
rect 22465 16575 22523 16581
rect 22465 16541 22477 16575
rect 22511 16541 22523 16575
rect 22465 16535 22523 16541
rect 24397 16575 24455 16581
rect 24397 16541 24409 16575
rect 24443 16572 24455 16575
rect 24670 16572 24676 16584
rect 24443 16544 24676 16572
rect 24443 16541 24455 16544
rect 24397 16535 24455 16541
rect 24670 16532 24676 16544
rect 24728 16532 24734 16584
rect 25222 16572 25228 16584
rect 25183 16544 25228 16572
rect 25222 16532 25228 16544
rect 25280 16532 25286 16584
rect 27062 16532 27068 16584
rect 27120 16572 27126 16584
rect 27522 16572 27528 16584
rect 27120 16544 27165 16572
rect 27483 16544 27528 16572
rect 27120 16532 27126 16544
rect 27522 16532 27528 16544
rect 27580 16532 27586 16584
rect 27614 16532 27620 16584
rect 27672 16572 27678 16584
rect 28810 16572 28816 16584
rect 27672 16544 27717 16572
rect 28771 16544 28816 16572
rect 27672 16532 27678 16544
rect 28810 16532 28816 16544
rect 28868 16532 28874 16584
rect 30116 16581 30144 16612
rect 31294 16600 31300 16652
rect 31352 16640 31358 16652
rect 32674 16640 32680 16652
rect 31352 16612 31524 16640
rect 32635 16612 32680 16640
rect 31352 16600 31358 16612
rect 30101 16575 30159 16581
rect 30101 16541 30113 16575
rect 30147 16541 30159 16575
rect 31496 16572 31524 16612
rect 32674 16600 32680 16612
rect 32732 16600 32738 16652
rect 35434 16640 35440 16652
rect 35395 16612 35440 16640
rect 35434 16600 35440 16612
rect 35492 16600 35498 16652
rect 42613 16643 42671 16649
rect 42613 16609 42625 16643
rect 42659 16640 42671 16643
rect 43254 16640 43260 16652
rect 42659 16612 43260 16640
rect 42659 16609 42671 16612
rect 42613 16603 42671 16609
rect 43254 16600 43260 16612
rect 43312 16600 43318 16652
rect 43806 16640 43812 16652
rect 43767 16612 43812 16640
rect 43806 16600 43812 16612
rect 43864 16600 43870 16652
rect 45833 16643 45891 16649
rect 45833 16609 45845 16643
rect 45879 16640 45891 16643
rect 46293 16643 46351 16649
rect 46293 16640 46305 16643
rect 45879 16612 46305 16640
rect 45879 16609 45891 16612
rect 45833 16603 45891 16609
rect 46293 16609 46305 16612
rect 46339 16609 46351 16643
rect 46293 16603 46351 16609
rect 31573 16575 31631 16581
rect 31573 16572 31585 16575
rect 31496 16544 31585 16572
rect 30101 16535 30159 16541
rect 31573 16541 31585 16544
rect 31619 16541 31631 16575
rect 32214 16572 32220 16584
rect 32175 16544 32220 16572
rect 31573 16535 31631 16541
rect 32214 16532 32220 16544
rect 32272 16532 32278 16584
rect 36906 16532 36912 16584
rect 36964 16572 36970 16584
rect 37366 16572 37372 16584
rect 36964 16544 37009 16572
rect 37327 16544 37372 16572
rect 36964 16532 36970 16544
rect 37366 16532 37372 16544
rect 37424 16532 37430 16584
rect 38473 16575 38531 16581
rect 38473 16541 38485 16575
rect 38519 16541 38531 16575
rect 38473 16535 38531 16541
rect 2317 16507 2375 16513
rect 2317 16473 2329 16507
rect 2363 16504 2375 16507
rect 3050 16504 3056 16516
rect 2363 16476 3056 16504
rect 2363 16473 2375 16476
rect 2317 16467 2375 16473
rect 3050 16464 3056 16476
rect 3108 16464 3114 16516
rect 4433 16507 4491 16513
rect 4433 16473 4445 16507
rect 4479 16504 4491 16507
rect 5626 16504 5632 16516
rect 4479 16476 5632 16504
rect 4479 16473 4491 16476
rect 4433 16467 4491 16473
rect 5626 16464 5632 16476
rect 5684 16464 5690 16516
rect 10318 16504 10324 16516
rect 10279 16476 10324 16504
rect 10318 16464 10324 16476
rect 10376 16464 10382 16516
rect 13449 16507 13507 16513
rect 13449 16473 13461 16507
rect 13495 16504 13507 16507
rect 14274 16504 14280 16516
rect 13495 16476 14280 16504
rect 13495 16473 13507 16476
rect 13449 16467 13507 16473
rect 14274 16464 14280 16476
rect 14332 16464 14338 16516
rect 15746 16504 15752 16516
rect 15707 16476 15752 16504
rect 15746 16464 15752 16476
rect 15804 16464 15810 16516
rect 21821 16507 21879 16513
rect 21821 16473 21833 16507
rect 21867 16504 21879 16507
rect 22554 16504 22560 16516
rect 21867 16476 22560 16504
rect 21867 16473 21879 16476
rect 21821 16467 21879 16473
rect 22554 16464 22560 16476
rect 22612 16464 22618 16516
rect 24578 16464 24584 16516
rect 24636 16504 24642 16516
rect 26881 16507 26939 16513
rect 26881 16504 26893 16507
rect 24636 16476 26893 16504
rect 24636 16464 24642 16476
rect 26881 16473 26893 16476
rect 26927 16473 26939 16507
rect 32398 16504 32404 16516
rect 32359 16476 32404 16504
rect 26881 16467 26939 16473
rect 32398 16464 32404 16476
rect 32456 16464 32462 16516
rect 35250 16464 35256 16516
rect 35308 16504 35314 16516
rect 36725 16507 36783 16513
rect 36725 16504 36737 16507
rect 35308 16476 36737 16504
rect 35308 16464 35314 16476
rect 36725 16473 36737 16476
rect 36771 16473 36783 16507
rect 36725 16467 36783 16473
rect 9674 16396 9680 16448
rect 9732 16436 9738 16448
rect 10594 16436 10600 16448
rect 9732 16408 10600 16436
rect 9732 16396 9738 16408
rect 10594 16396 10600 16408
rect 10652 16396 10658 16448
rect 33778 16396 33784 16448
rect 33836 16436 33842 16448
rect 38488 16436 38516 16535
rect 38930 16532 38936 16584
rect 38988 16572 38994 16584
rect 39117 16575 39175 16581
rect 39117 16572 39129 16575
rect 38988 16544 39129 16572
rect 38988 16532 38994 16544
rect 39117 16541 39129 16544
rect 39163 16541 39175 16575
rect 39850 16572 39856 16584
rect 39811 16544 39856 16572
rect 39117 16535 39175 16541
rect 39850 16532 39856 16544
rect 39908 16532 39914 16584
rect 39945 16575 40003 16581
rect 39945 16541 39957 16575
rect 39991 16572 40003 16575
rect 40126 16572 40132 16584
rect 39991 16544 40132 16572
rect 39991 16541 40003 16544
rect 39945 16535 40003 16541
rect 40126 16532 40132 16544
rect 40184 16532 40190 16584
rect 45005 16575 45063 16581
rect 45005 16541 45017 16575
rect 45051 16541 45063 16575
rect 45005 16535 45063 16541
rect 48133 16575 48191 16581
rect 48133 16541 48145 16575
rect 48179 16572 48191 16575
rect 48314 16572 48320 16584
rect 48179 16544 48320 16572
rect 48179 16541 48191 16544
rect 48133 16535 48191 16541
rect 42797 16507 42855 16513
rect 42797 16473 42809 16507
rect 42843 16504 42855 16507
rect 43438 16504 43444 16516
rect 42843 16476 43444 16504
rect 42843 16473 42855 16476
rect 42797 16467 42855 16473
rect 43438 16464 43444 16476
rect 43496 16464 43502 16516
rect 33836 16408 38516 16436
rect 38565 16439 38623 16445
rect 33836 16396 33842 16408
rect 38565 16405 38577 16439
rect 38611 16436 38623 16439
rect 39114 16436 39120 16448
rect 38611 16408 39120 16436
rect 38611 16405 38623 16408
rect 38565 16399 38623 16405
rect 39114 16396 39120 16408
rect 39172 16396 39178 16448
rect 43162 16396 43168 16448
rect 43220 16436 43226 16448
rect 45020 16436 45048 16535
rect 48314 16532 48320 16544
rect 48372 16532 48378 16584
rect 46477 16507 46535 16513
rect 46477 16473 46489 16507
rect 46523 16504 46535 16507
rect 47670 16504 47676 16516
rect 46523 16476 47676 16504
rect 46523 16473 46535 16476
rect 46477 16467 46535 16473
rect 47670 16464 47676 16476
rect 47728 16464 47734 16516
rect 43220 16408 45048 16436
rect 43220 16396 43226 16408
rect 1104 16346 48852 16368
rect 1104 16294 16880 16346
rect 16932 16294 16944 16346
rect 16996 16294 17008 16346
rect 17060 16294 17072 16346
rect 17124 16294 17136 16346
rect 17188 16294 32811 16346
rect 32863 16294 32875 16346
rect 32927 16294 32939 16346
rect 32991 16294 33003 16346
rect 33055 16294 33067 16346
rect 33119 16294 48852 16346
rect 1104 16272 48852 16294
rect 7558 16192 7564 16244
rect 7616 16232 7622 16244
rect 7929 16235 7987 16241
rect 7929 16232 7941 16235
rect 7616 16204 7941 16232
rect 7616 16192 7622 16204
rect 7929 16201 7941 16204
rect 7975 16201 7987 16235
rect 10318 16232 10324 16244
rect 10279 16204 10324 16232
rect 7929 16195 7987 16201
rect 10318 16192 10324 16204
rect 10376 16192 10382 16244
rect 12434 16232 12440 16244
rect 12360 16204 12440 16232
rect 8021 16099 8079 16105
rect 8021 16065 8033 16099
rect 8067 16065 8079 16099
rect 10226 16096 10232 16108
rect 10187 16068 10232 16096
rect 8021 16059 8079 16065
rect 8036 15960 8064 16059
rect 10226 16056 10232 16068
rect 10284 16056 10290 16108
rect 12360 16105 12388 16204
rect 12434 16192 12440 16204
rect 12492 16192 12498 16244
rect 15746 16232 15752 16244
rect 15707 16204 15752 16232
rect 15746 16192 15752 16204
rect 15804 16192 15810 16244
rect 24578 16232 24584 16244
rect 24539 16204 24584 16232
rect 24578 16192 24584 16204
rect 24636 16192 24642 16244
rect 32398 16232 32404 16244
rect 32359 16204 32404 16232
rect 32398 16192 32404 16204
rect 32456 16192 32462 16244
rect 33873 16235 33931 16241
rect 33873 16201 33885 16235
rect 33919 16232 33931 16235
rect 34882 16232 34888 16244
rect 33919 16204 34888 16232
rect 33919 16201 33931 16204
rect 33873 16195 33931 16201
rect 34882 16192 34888 16204
rect 34940 16192 34946 16244
rect 35250 16232 35256 16244
rect 35211 16204 35256 16232
rect 35250 16192 35256 16204
rect 35308 16192 35314 16244
rect 42613 16235 42671 16241
rect 42613 16201 42625 16235
rect 42659 16232 42671 16235
rect 42702 16232 42708 16244
rect 42659 16204 42708 16232
rect 42659 16201 42671 16204
rect 42613 16195 42671 16201
rect 42702 16192 42708 16204
rect 42760 16192 42766 16244
rect 43438 16232 43444 16244
rect 43399 16204 43444 16232
rect 43438 16192 43444 16204
rect 43496 16192 43502 16244
rect 47670 16232 47676 16244
rect 47631 16204 47676 16232
rect 47670 16192 47676 16204
rect 47728 16192 47734 16244
rect 22094 16124 22100 16176
rect 22152 16164 22158 16176
rect 28994 16164 29000 16176
rect 22152 16136 29000 16164
rect 22152 16124 22158 16136
rect 12345 16099 12403 16105
rect 12345 16065 12357 16099
rect 12391 16065 12403 16099
rect 12345 16059 12403 16065
rect 15562 16056 15568 16108
rect 15620 16096 15626 16108
rect 15657 16099 15715 16105
rect 15657 16096 15669 16099
rect 15620 16068 15669 16096
rect 15620 16056 15626 16068
rect 15657 16065 15669 16068
rect 15703 16065 15715 16099
rect 18230 16096 18236 16108
rect 18191 16068 18236 16096
rect 15657 16059 15715 16065
rect 18230 16056 18236 16068
rect 18288 16056 18294 16108
rect 24029 16099 24087 16105
rect 24029 16065 24041 16099
rect 24075 16096 24087 16099
rect 24394 16096 24400 16108
rect 24075 16068 24400 16096
rect 24075 16065 24087 16068
rect 24029 16059 24087 16065
rect 24394 16056 24400 16068
rect 24452 16056 24458 16108
rect 24504 16105 24532 16136
rect 28994 16124 29000 16136
rect 29052 16124 29058 16176
rect 30653 16167 30711 16173
rect 30653 16133 30665 16167
rect 30699 16164 30711 16167
rect 45554 16164 45560 16176
rect 30699 16136 45560 16164
rect 30699 16133 30711 16136
rect 30653 16127 30711 16133
rect 45554 16124 45560 16136
rect 45612 16124 45618 16176
rect 24489 16099 24547 16105
rect 24489 16065 24501 16099
rect 24535 16065 24547 16099
rect 24489 16059 24547 16065
rect 24670 16056 24676 16108
rect 24728 16096 24734 16108
rect 25133 16099 25191 16105
rect 25133 16096 25145 16099
rect 24728 16068 25145 16096
rect 24728 16056 24734 16068
rect 25133 16065 25145 16068
rect 25179 16065 25191 16099
rect 25133 16059 25191 16065
rect 26237 16099 26295 16105
rect 26237 16065 26249 16099
rect 26283 16096 26295 16099
rect 26973 16099 27031 16105
rect 26283 16068 26924 16096
rect 26283 16065 26295 16068
rect 26237 16059 26295 16065
rect 12526 16028 12532 16040
rect 12487 16000 12532 16028
rect 12526 15988 12532 16000
rect 12584 15988 12590 16040
rect 12894 16028 12900 16040
rect 12855 16000 12900 16028
rect 12894 15988 12900 16000
rect 12952 15988 12958 16040
rect 18417 16031 18475 16037
rect 18417 15997 18429 16031
rect 18463 16028 18475 16031
rect 18506 16028 18512 16040
rect 18463 16000 18512 16028
rect 18463 15997 18475 16000
rect 18417 15991 18475 15997
rect 18506 15988 18512 16000
rect 18564 15988 18570 16040
rect 18690 16028 18696 16040
rect 18651 16000 18696 16028
rect 18690 15988 18696 16000
rect 18748 15988 18754 16040
rect 19242 15988 19248 16040
rect 19300 16028 19306 16040
rect 25314 16028 25320 16040
rect 19300 16000 25320 16028
rect 19300 15988 19306 16000
rect 25314 15988 25320 16000
rect 25372 15988 25378 16040
rect 19610 15960 19616 15972
rect 8036 15932 19616 15960
rect 19610 15920 19616 15932
rect 19668 15920 19674 15972
rect 26896 15960 26924 16068
rect 26973 16065 26985 16099
rect 27019 16096 27031 16099
rect 27062 16096 27068 16108
rect 27019 16068 27068 16096
rect 27019 16065 27031 16068
rect 26973 16059 27031 16065
rect 27062 16056 27068 16068
rect 27120 16056 27126 16108
rect 28810 16096 28816 16108
rect 28771 16068 28816 16096
rect 28810 16056 28816 16068
rect 28868 16056 28874 16108
rect 31573 16099 31631 16105
rect 31573 16065 31585 16099
rect 31619 16096 31631 16099
rect 32122 16096 32128 16108
rect 31619 16068 32128 16096
rect 31619 16065 31631 16068
rect 31573 16059 31631 16065
rect 32122 16056 32128 16068
rect 32180 16056 32186 16108
rect 32493 16099 32551 16105
rect 32493 16065 32505 16099
rect 32539 16096 32551 16099
rect 32674 16096 32680 16108
rect 32539 16068 32680 16096
rect 32539 16065 32551 16068
rect 32493 16059 32551 16065
rect 32674 16056 32680 16068
rect 32732 16096 32738 16108
rect 32732 16068 33732 16096
rect 32732 16056 32738 16068
rect 28442 15988 28448 16040
rect 28500 16028 28506 16040
rect 28997 16031 29055 16037
rect 28997 16028 29009 16031
rect 28500 16000 29009 16028
rect 28500 15988 28506 16000
rect 28997 15997 29009 16000
rect 29043 15997 29055 16031
rect 28997 15991 29055 15997
rect 32214 15988 32220 16040
rect 32272 16028 32278 16040
rect 32953 16031 33011 16037
rect 32953 16028 32965 16031
rect 32272 16000 32965 16028
rect 32272 15988 32278 16000
rect 32953 15997 32965 16000
rect 32999 15997 33011 16031
rect 33704 16028 33732 16068
rect 33778 16056 33784 16108
rect 33836 16096 33842 16108
rect 34609 16099 34667 16105
rect 33836 16068 33881 16096
rect 33836 16056 33842 16068
rect 34609 16065 34621 16099
rect 34655 16096 34667 16099
rect 34698 16096 34704 16108
rect 34655 16068 34704 16096
rect 34655 16065 34667 16068
rect 34609 16059 34667 16065
rect 34698 16056 34704 16068
rect 34756 16056 34762 16108
rect 35161 16099 35219 16105
rect 35161 16065 35173 16099
rect 35207 16065 35219 16099
rect 35161 16059 35219 16065
rect 36633 16099 36691 16105
rect 36633 16065 36645 16099
rect 36679 16096 36691 16099
rect 36906 16096 36912 16108
rect 36679 16068 36912 16096
rect 36679 16065 36691 16068
rect 36633 16059 36691 16065
rect 35176 16028 35204 16059
rect 36906 16056 36912 16068
rect 36964 16056 36970 16108
rect 37274 16096 37280 16108
rect 37235 16068 37280 16096
rect 37274 16056 37280 16068
rect 37332 16056 37338 16108
rect 38930 16096 38936 16108
rect 38891 16068 38936 16096
rect 38930 16056 38936 16068
rect 38988 16056 38994 16108
rect 40773 16099 40831 16105
rect 40773 16065 40785 16099
rect 40819 16096 40831 16099
rect 42426 16096 42432 16108
rect 40819 16068 42432 16096
rect 40819 16065 40831 16068
rect 40773 16059 40831 16065
rect 42426 16056 42432 16068
rect 42484 16056 42490 16108
rect 42521 16099 42579 16105
rect 42521 16065 42533 16099
rect 42567 16096 42579 16099
rect 43162 16096 43168 16108
rect 42567 16068 43168 16096
rect 42567 16065 42579 16068
rect 42521 16059 42579 16065
rect 43162 16056 43168 16068
rect 43220 16056 43226 16108
rect 43533 16099 43591 16105
rect 43533 16065 43545 16099
rect 43579 16065 43591 16099
rect 44726 16096 44732 16108
rect 44687 16068 44732 16096
rect 43533 16059 43591 16065
rect 39114 16028 39120 16040
rect 33704 16000 35204 16028
rect 39075 16000 39120 16028
rect 32953 15991 33011 15997
rect 39114 15988 39120 16000
rect 39172 15988 39178 16040
rect 42794 15988 42800 16040
rect 42852 16028 42858 16040
rect 43548 16028 43576 16059
rect 44726 16056 44732 16068
rect 44784 16056 44790 16108
rect 47302 16056 47308 16108
rect 47360 16096 47366 16108
rect 47581 16099 47639 16105
rect 47581 16096 47593 16099
rect 47360 16068 47593 16096
rect 47360 16056 47366 16068
rect 47581 16065 47593 16068
rect 47627 16065 47639 16099
rect 47581 16059 47639 16065
rect 42852 16000 43576 16028
rect 45189 16031 45247 16037
rect 42852 15988 42858 16000
rect 45189 15997 45201 16031
rect 45235 15997 45247 16031
rect 45370 16028 45376 16040
rect 45331 16000 45376 16028
rect 45189 15991 45247 15997
rect 26970 15960 26976 15972
rect 26883 15932 26976 15960
rect 26970 15920 26976 15932
rect 27028 15960 27034 15972
rect 28534 15960 28540 15972
rect 27028 15932 28540 15960
rect 27028 15920 27034 15932
rect 28534 15920 28540 15932
rect 28592 15920 28598 15972
rect 45204 15960 45232 15991
rect 45370 15988 45376 16000
rect 45428 15988 45434 16040
rect 46842 16028 46848 16040
rect 46803 16000 46848 16028
rect 46842 15988 46848 16000
rect 46900 15988 46906 16040
rect 45554 15960 45560 15972
rect 45204 15932 45560 15960
rect 45554 15920 45560 15932
rect 45612 15920 45618 15972
rect 2038 15892 2044 15904
rect 1999 15864 2044 15892
rect 2038 15852 2044 15864
rect 2096 15852 2102 15904
rect 11698 15892 11704 15904
rect 11659 15864 11704 15892
rect 11698 15852 11704 15864
rect 11756 15852 11762 15904
rect 16114 15852 16120 15904
rect 16172 15892 16178 15904
rect 16669 15895 16727 15901
rect 16669 15892 16681 15895
rect 16172 15864 16681 15892
rect 16172 15852 16178 15864
rect 16669 15861 16681 15864
rect 16715 15861 16727 15895
rect 16669 15855 16727 15861
rect 25406 15852 25412 15904
rect 25464 15892 25470 15904
rect 26145 15895 26203 15901
rect 26145 15892 26157 15895
rect 25464 15864 26157 15892
rect 25464 15852 25470 15864
rect 26145 15861 26157 15864
rect 26191 15861 26203 15895
rect 26145 15855 26203 15861
rect 35618 15852 35624 15904
rect 35676 15892 35682 15904
rect 35805 15895 35863 15901
rect 35805 15892 35817 15895
rect 35676 15864 35817 15892
rect 35676 15852 35682 15864
rect 35805 15861 35817 15864
rect 35851 15861 35863 15895
rect 41230 15892 41236 15904
rect 41191 15864 41236 15892
rect 35805 15855 35863 15861
rect 41230 15852 41236 15864
rect 41288 15852 41294 15904
rect 1104 15802 48852 15824
rect 1104 15750 8915 15802
rect 8967 15750 8979 15802
rect 9031 15750 9043 15802
rect 9095 15750 9107 15802
rect 9159 15750 9171 15802
rect 9223 15750 24846 15802
rect 24898 15750 24910 15802
rect 24962 15750 24974 15802
rect 25026 15750 25038 15802
rect 25090 15750 25102 15802
rect 25154 15750 40776 15802
rect 40828 15750 40840 15802
rect 40892 15750 40904 15802
rect 40956 15750 40968 15802
rect 41020 15750 41032 15802
rect 41084 15750 48852 15802
rect 1104 15728 48852 15750
rect 18506 15688 18512 15700
rect 18467 15660 18512 15688
rect 18506 15648 18512 15660
rect 18564 15648 18570 15700
rect 28442 15688 28448 15700
rect 28403 15660 28448 15688
rect 28442 15648 28448 15660
rect 28500 15648 28506 15700
rect 28534 15648 28540 15700
rect 28592 15688 28598 15700
rect 42794 15688 42800 15700
rect 28592 15660 42800 15688
rect 28592 15648 28598 15660
rect 42794 15648 42800 15660
rect 42852 15648 42858 15700
rect 43254 15688 43260 15700
rect 43215 15660 43260 15688
rect 43254 15648 43260 15660
rect 43312 15648 43318 15700
rect 45281 15691 45339 15697
rect 45281 15657 45293 15691
rect 45327 15688 45339 15691
rect 45370 15688 45376 15700
rect 45327 15660 45376 15688
rect 45327 15657 45339 15660
rect 45281 15651 45339 15657
rect 45370 15648 45376 15660
rect 45428 15648 45434 15700
rect 15562 15580 15568 15632
rect 15620 15620 15626 15632
rect 22094 15620 22100 15632
rect 15620 15592 22100 15620
rect 15620 15580 15626 15592
rect 22094 15580 22100 15592
rect 22152 15580 22158 15632
rect 22204 15592 40172 15620
rect 11698 15552 11704 15564
rect 11659 15524 11704 15552
rect 11698 15512 11704 15524
rect 11756 15512 11762 15564
rect 12250 15512 12256 15564
rect 12308 15552 12314 15564
rect 12437 15555 12495 15561
rect 12437 15552 12449 15555
rect 12308 15524 12449 15552
rect 12308 15512 12314 15524
rect 12437 15521 12449 15524
rect 12483 15521 12495 15555
rect 16114 15552 16120 15564
rect 16075 15524 16120 15552
rect 12437 15515 12495 15521
rect 16114 15512 16120 15524
rect 16172 15512 16178 15564
rect 16758 15552 16764 15564
rect 16719 15524 16764 15552
rect 16758 15512 16764 15524
rect 16816 15512 16822 15564
rect 22204 15552 22232 15592
rect 25222 15552 25228 15564
rect 22066 15524 22232 15552
rect 25183 15524 25228 15552
rect 2406 15444 2412 15496
rect 2464 15484 2470 15496
rect 2501 15487 2559 15493
rect 2501 15484 2513 15487
rect 2464 15456 2513 15484
rect 2464 15444 2470 15456
rect 2501 15453 2513 15456
rect 2547 15453 2559 15487
rect 15654 15484 15660 15496
rect 15615 15456 15660 15484
rect 2501 15447 2559 15453
rect 15654 15444 15660 15456
rect 15712 15444 15718 15496
rect 18414 15444 18420 15496
rect 18472 15484 18478 15496
rect 18601 15487 18659 15493
rect 18601 15484 18613 15487
rect 18472 15456 18613 15484
rect 18472 15444 18478 15456
rect 18601 15453 18613 15456
rect 18647 15484 18659 15487
rect 19242 15484 19248 15496
rect 18647 15456 19248 15484
rect 18647 15453 18659 15456
rect 18601 15447 18659 15453
rect 19242 15444 19248 15456
rect 19300 15444 19306 15496
rect 19886 15484 19892 15496
rect 19847 15456 19892 15484
rect 19886 15444 19892 15456
rect 19944 15444 19950 15496
rect 11882 15416 11888 15428
rect 11843 15388 11888 15416
rect 11882 15376 11888 15388
rect 11940 15376 11946 15428
rect 15565 15419 15623 15425
rect 15565 15385 15577 15419
rect 15611 15416 15623 15419
rect 16301 15419 16359 15425
rect 16301 15416 16313 15419
rect 15611 15388 16313 15416
rect 15611 15385 15623 15388
rect 15565 15379 15623 15385
rect 16301 15385 16313 15388
rect 16347 15385 16359 15419
rect 19426 15416 19432 15428
rect 19387 15388 19432 15416
rect 16301 15379 16359 15385
rect 19426 15376 19432 15388
rect 19484 15416 19490 15428
rect 22066 15416 22094 15524
rect 25222 15512 25228 15524
rect 25280 15512 25286 15564
rect 25406 15552 25412 15564
rect 25367 15524 25412 15552
rect 25406 15512 25412 15524
rect 25464 15512 25470 15564
rect 25774 15552 25780 15564
rect 25735 15524 25780 15552
rect 25774 15512 25780 15524
rect 25832 15512 25838 15564
rect 35618 15552 35624 15564
rect 35579 15524 35624 15552
rect 35618 15512 35624 15524
rect 35676 15512 35682 15564
rect 36078 15552 36084 15564
rect 36039 15524 36084 15552
rect 36078 15512 36084 15524
rect 36136 15512 36142 15564
rect 40144 15496 40172 15592
rect 40865 15555 40923 15561
rect 40865 15521 40877 15555
rect 40911 15552 40923 15555
rect 41230 15552 41236 15564
rect 40911 15524 41236 15552
rect 40911 15521 40923 15524
rect 40865 15515 40923 15521
rect 41230 15512 41236 15524
rect 41288 15512 41294 15564
rect 41874 15552 41880 15564
rect 41835 15524 41880 15552
rect 41874 15512 41880 15524
rect 41932 15512 41938 15564
rect 27706 15444 27712 15496
rect 27764 15484 27770 15496
rect 28353 15487 28411 15493
rect 28353 15484 28365 15487
rect 27764 15456 28365 15484
rect 27764 15444 27770 15456
rect 28353 15453 28365 15456
rect 28399 15453 28411 15487
rect 28353 15447 28411 15453
rect 40126 15444 40132 15496
rect 40184 15484 40190 15496
rect 40221 15487 40279 15493
rect 40221 15484 40233 15487
rect 40184 15456 40233 15484
rect 40184 15444 40190 15456
rect 40221 15453 40233 15456
rect 40267 15453 40279 15487
rect 42812 15484 42840 15648
rect 46750 15552 46756 15564
rect 46711 15524 46756 15552
rect 46750 15512 46756 15524
rect 46808 15512 46814 15564
rect 47762 15512 47768 15564
rect 47820 15552 47826 15564
rect 48133 15555 48191 15561
rect 48133 15552 48145 15555
rect 47820 15524 48145 15552
rect 47820 15512 47826 15524
rect 48133 15521 48145 15524
rect 48179 15521 48191 15555
rect 48133 15515 48191 15521
rect 45189 15487 45247 15493
rect 45189 15484 45201 15487
rect 42812 15456 45201 15484
rect 40221 15447 40279 15453
rect 45189 15453 45201 15456
rect 45235 15453 45247 15487
rect 45189 15447 45247 15453
rect 24578 15416 24584 15428
rect 19484 15388 22094 15416
rect 24539 15388 24584 15416
rect 19484 15376 19490 15388
rect 24578 15376 24584 15388
rect 24636 15376 24642 15428
rect 35805 15419 35863 15425
rect 35805 15385 35817 15419
rect 35851 15416 35863 15419
rect 35894 15416 35900 15428
rect 35851 15388 35900 15416
rect 35851 15385 35863 15388
rect 35805 15379 35863 15385
rect 35894 15376 35900 15388
rect 35952 15376 35958 15428
rect 40313 15419 40371 15425
rect 40313 15385 40325 15419
rect 40359 15416 40371 15419
rect 41049 15419 41107 15425
rect 41049 15416 41061 15419
rect 40359 15388 41061 15416
rect 40359 15385 40371 15388
rect 40313 15379 40371 15385
rect 41049 15385 41061 15388
rect 41095 15385 41107 15419
rect 47946 15416 47952 15428
rect 47907 15388 47952 15416
rect 41049 15379 41107 15385
rect 47946 15376 47952 15388
rect 48004 15376 48010 15428
rect 2222 15308 2228 15360
rect 2280 15348 2286 15360
rect 2409 15351 2467 15357
rect 2409 15348 2421 15351
rect 2280 15320 2421 15348
rect 2280 15308 2286 15320
rect 2409 15317 2421 15320
rect 2455 15317 2467 15351
rect 24670 15348 24676 15360
rect 24631 15320 24676 15348
rect 2409 15311 2467 15317
rect 24670 15308 24676 15320
rect 24728 15308 24734 15360
rect 1104 15258 48852 15280
rect 1104 15206 16880 15258
rect 16932 15206 16944 15258
rect 16996 15206 17008 15258
rect 17060 15206 17072 15258
rect 17124 15206 17136 15258
rect 17188 15206 32811 15258
rect 32863 15206 32875 15258
rect 32927 15206 32939 15258
rect 32991 15206 33003 15258
rect 33055 15206 33067 15258
rect 33119 15206 48852 15258
rect 1104 15184 48852 15206
rect 11882 15144 11888 15156
rect 11843 15116 11888 15144
rect 11882 15104 11888 15116
rect 11940 15104 11946 15156
rect 12526 15144 12532 15156
rect 12487 15116 12532 15144
rect 12526 15104 12532 15116
rect 12584 15104 12590 15156
rect 17954 15104 17960 15156
rect 18012 15144 18018 15156
rect 18322 15144 18328 15156
rect 18012 15116 18328 15144
rect 18012 15104 18018 15116
rect 18322 15104 18328 15116
rect 18380 15144 18386 15156
rect 27522 15144 27528 15156
rect 18380 15116 27528 15144
rect 18380 15104 18386 15116
rect 27522 15104 27528 15116
rect 27580 15104 27586 15156
rect 27614 15104 27620 15156
rect 27672 15144 27678 15156
rect 33778 15144 33784 15156
rect 27672 15116 33784 15144
rect 27672 15104 27678 15116
rect 33778 15104 33784 15116
rect 33836 15104 33842 15156
rect 35894 15104 35900 15156
rect 35952 15144 35958 15156
rect 47673 15147 47731 15153
rect 35952 15116 35997 15144
rect 35952 15104 35958 15116
rect 47673 15113 47685 15147
rect 47719 15144 47731 15147
rect 47946 15144 47952 15156
rect 47719 15116 47952 15144
rect 47719 15113 47731 15116
rect 47673 15107 47731 15113
rect 47946 15104 47952 15116
rect 48004 15104 48010 15156
rect 2222 15076 2228 15088
rect 2183 15048 2228 15076
rect 2222 15036 2228 15048
rect 2280 15036 2286 15088
rect 18046 15036 18052 15088
rect 18104 15076 18110 15088
rect 25866 15076 25872 15088
rect 18104 15048 25872 15076
rect 18104 15036 18110 15048
rect 25866 15036 25872 15048
rect 25924 15036 25930 15088
rect 36004 15048 46796 15076
rect 36004 15020 36032 15048
rect 46768 15020 46796 15048
rect 2038 15008 2044 15020
rect 1999 14980 2044 15008
rect 2038 14968 2044 14980
rect 2096 14968 2102 15020
rect 11790 15008 11796 15020
rect 11751 14980 11796 15008
rect 11790 14968 11796 14980
rect 11848 14968 11854 15020
rect 12434 15008 12440 15020
rect 12395 14980 12440 15008
rect 12434 14968 12440 14980
rect 12492 14968 12498 15020
rect 18506 15008 18512 15020
rect 18467 14980 18512 15008
rect 18506 14968 18512 14980
rect 18564 15008 18570 15020
rect 18969 15011 19027 15017
rect 18969 15008 18981 15011
rect 18564 14980 18981 15008
rect 18564 14968 18570 14980
rect 18969 14977 18981 14980
rect 19015 15008 19027 15011
rect 19886 15008 19892 15020
rect 19015 14980 19892 15008
rect 19015 14977 19027 14980
rect 18969 14971 19027 14977
rect 19886 14968 19892 14980
rect 19944 15008 19950 15020
rect 20349 15011 20407 15017
rect 20349 15008 20361 15011
rect 19944 14980 20361 15008
rect 19944 14968 19950 14980
rect 20349 14977 20361 14980
rect 20395 14977 20407 15011
rect 24670 15008 24676 15020
rect 24583 14980 24676 15008
rect 20349 14971 20407 14977
rect 24670 14968 24676 14980
rect 24728 15008 24734 15020
rect 25133 15011 25191 15017
rect 25133 15008 25145 15011
rect 24728 14980 25145 15008
rect 24728 14968 24734 14980
rect 25133 14977 25145 14980
rect 25179 15008 25191 15011
rect 25222 15008 25228 15020
rect 25179 14980 25228 15008
rect 25179 14977 25191 14980
rect 25133 14971 25191 14977
rect 25222 14968 25228 14980
rect 25280 14968 25286 15020
rect 27065 15011 27123 15017
rect 27065 14977 27077 15011
rect 27111 14977 27123 15011
rect 27065 14971 27123 14977
rect 27249 15011 27307 15017
rect 27249 14977 27261 15011
rect 27295 15008 27307 15011
rect 28169 15011 28227 15017
rect 28169 15008 28181 15011
rect 27295 14980 28181 15008
rect 27295 14977 27307 14980
rect 27249 14971 27307 14977
rect 28169 14977 28181 14980
rect 28215 15008 28227 15011
rect 28721 15011 28779 15017
rect 28721 15008 28733 15011
rect 28215 14980 28733 15008
rect 28215 14977 28227 14980
rect 28169 14971 28227 14977
rect 28721 14977 28733 14980
rect 28767 15008 28779 15011
rect 30929 15011 30987 15017
rect 30929 15008 30941 15011
rect 28767 14980 30941 15008
rect 28767 14977 28779 14980
rect 28721 14971 28779 14977
rect 30929 14977 30941 14980
rect 30975 15008 30987 15011
rect 31662 15008 31668 15020
rect 30975 14980 31668 15008
rect 30975 14977 30987 14980
rect 30929 14971 30987 14977
rect 2774 14900 2780 14952
rect 2832 14940 2838 14952
rect 2832 14912 2877 14940
rect 2832 14900 2838 14912
rect 15654 14900 15660 14952
rect 15712 14940 15718 14952
rect 15712 14912 18276 14940
rect 15712 14900 15718 14912
rect 11790 14832 11796 14884
rect 11848 14872 11854 14884
rect 18248 14872 18276 14912
rect 18322 14900 18328 14952
rect 18380 14940 18386 14952
rect 19702 14940 19708 14952
rect 18380 14912 18425 14940
rect 19663 14912 19708 14940
rect 18380 14900 18386 14912
rect 19702 14900 19708 14912
rect 19760 14900 19766 14952
rect 20622 14940 20628 14952
rect 20583 14912 20628 14940
rect 20622 14900 20628 14912
rect 20680 14900 20686 14952
rect 24486 14940 24492 14952
rect 24447 14912 24492 14940
rect 24486 14900 24492 14912
rect 24544 14900 24550 14952
rect 24578 14900 24584 14952
rect 24636 14940 24642 14952
rect 27080 14940 27108 14971
rect 31662 14968 31668 14980
rect 31720 15008 31726 15020
rect 32125 15011 32183 15017
rect 32125 15008 32137 15011
rect 31720 14980 32137 15008
rect 31720 14968 31726 14980
rect 32125 14977 32137 14980
rect 32171 14977 32183 15011
rect 35986 15008 35992 15020
rect 35899 14980 35992 15008
rect 32125 14971 32183 14977
rect 35986 14968 35992 14980
rect 36044 14968 36050 15020
rect 45554 14968 45560 15020
rect 45612 15008 45618 15020
rect 45612 14980 45657 15008
rect 45612 14968 45618 14980
rect 46750 14968 46756 15020
rect 46808 15008 46814 15020
rect 46845 15011 46903 15017
rect 46845 15008 46857 15011
rect 46808 14980 46857 15008
rect 46808 14968 46814 14980
rect 46845 14977 46857 14980
rect 46891 14977 46903 15011
rect 46845 14971 46903 14977
rect 47581 15011 47639 15017
rect 47581 14977 47593 15011
rect 47627 14977 47639 15011
rect 47581 14971 47639 14977
rect 27798 14940 27804 14952
rect 24636 14912 27804 14940
rect 24636 14900 24642 14912
rect 27798 14900 27804 14912
rect 27856 14900 27862 14952
rect 28997 14943 29055 14949
rect 28997 14909 29009 14943
rect 29043 14909 29055 14943
rect 28997 14903 29055 14909
rect 31389 14943 31447 14949
rect 31389 14909 31401 14943
rect 31435 14909 31447 14943
rect 31389 14903 31447 14909
rect 32401 14943 32459 14949
rect 32401 14909 32413 14943
rect 32447 14940 32459 14943
rect 32674 14940 32680 14952
rect 32447 14912 32680 14940
rect 32447 14909 32459 14912
rect 32401 14903 32459 14909
rect 29012 14872 29040 14903
rect 29086 14872 29092 14884
rect 11848 14844 18184 14872
rect 18248 14844 29092 14872
rect 11848 14832 11854 14844
rect 12434 14764 12440 14816
rect 12492 14804 12498 14816
rect 18046 14804 18052 14816
rect 12492 14776 18052 14804
rect 12492 14764 12498 14776
rect 18046 14764 18052 14776
rect 18104 14764 18110 14816
rect 18156 14804 18184 14844
rect 29086 14832 29092 14844
rect 29144 14832 29150 14884
rect 20622 14804 20628 14816
rect 18156 14776 20628 14804
rect 20622 14764 20628 14776
rect 20680 14764 20686 14816
rect 24486 14764 24492 14816
rect 24544 14804 24550 14816
rect 27614 14804 27620 14816
rect 24544 14776 27620 14804
rect 24544 14764 24550 14776
rect 27614 14764 27620 14776
rect 27672 14764 27678 14816
rect 27706 14764 27712 14816
rect 27764 14804 27770 14816
rect 27893 14807 27951 14813
rect 27893 14804 27905 14807
rect 27764 14776 27905 14804
rect 27764 14764 27770 14776
rect 27893 14773 27905 14776
rect 27939 14773 27951 14807
rect 31404 14804 31432 14903
rect 32674 14900 32680 14912
rect 32732 14900 32738 14952
rect 46934 14940 46940 14952
rect 35866 14912 46940 14940
rect 35866 14872 35894 14912
rect 46934 14900 46940 14912
rect 46992 14940 46998 14952
rect 47596 14940 47624 14971
rect 46992 14912 47624 14940
rect 46992 14900 46998 14912
rect 31726 14844 35894 14872
rect 31478 14804 31484 14816
rect 31404 14776 31484 14804
rect 27893 14767 27951 14773
rect 31478 14764 31484 14776
rect 31536 14804 31542 14816
rect 31726 14804 31754 14844
rect 31536 14776 31754 14804
rect 31536 14764 31542 14776
rect 46290 14764 46296 14816
rect 46348 14804 46354 14816
rect 46385 14807 46443 14813
rect 46385 14804 46397 14807
rect 46348 14776 46397 14804
rect 46348 14764 46354 14776
rect 46385 14773 46397 14776
rect 46431 14773 46443 14807
rect 46385 14767 46443 14773
rect 46474 14764 46480 14816
rect 46532 14804 46538 14816
rect 46937 14807 46995 14813
rect 46937 14804 46949 14807
rect 46532 14776 46949 14804
rect 46532 14764 46538 14776
rect 46937 14773 46949 14776
rect 46983 14773 46995 14807
rect 46937 14767 46995 14773
rect 1104 14714 48852 14736
rect 1104 14662 8915 14714
rect 8967 14662 8979 14714
rect 9031 14662 9043 14714
rect 9095 14662 9107 14714
rect 9159 14662 9171 14714
rect 9223 14662 24846 14714
rect 24898 14662 24910 14714
rect 24962 14662 24974 14714
rect 25026 14662 25038 14714
rect 25090 14662 25102 14714
rect 25154 14662 40776 14714
rect 40828 14662 40840 14714
rect 40892 14662 40904 14714
rect 40956 14662 40968 14714
rect 41020 14662 41032 14714
rect 41084 14662 48852 14714
rect 1104 14640 48852 14662
rect 18506 14600 18512 14612
rect 18467 14572 18512 14600
rect 18506 14560 18512 14572
rect 18564 14560 18570 14612
rect 1949 14399 2007 14405
rect 1949 14365 1961 14399
rect 1995 14396 2007 14399
rect 2038 14396 2044 14408
rect 1995 14368 2044 14396
rect 1995 14365 2007 14368
rect 1949 14359 2007 14365
rect 2038 14356 2044 14368
rect 2096 14356 2102 14408
rect 2593 14399 2651 14405
rect 2593 14365 2605 14399
rect 2639 14396 2651 14399
rect 2682 14396 2688 14408
rect 2639 14368 2688 14396
rect 2639 14365 2651 14368
rect 2593 14359 2651 14365
rect 2682 14356 2688 14368
rect 2740 14396 2746 14408
rect 7742 14396 7748 14408
rect 2740 14368 7748 14396
rect 2740 14356 2746 14368
rect 7742 14356 7748 14368
rect 7800 14356 7806 14408
rect 18524 14396 18552 14560
rect 19610 14464 19616 14476
rect 19523 14436 19616 14464
rect 19610 14424 19616 14436
rect 19668 14464 19674 14476
rect 39850 14464 39856 14476
rect 19668 14436 39856 14464
rect 19668 14424 19674 14436
rect 39850 14424 39856 14436
rect 39908 14424 39914 14476
rect 46290 14464 46296 14476
rect 46251 14436 46296 14464
rect 46290 14424 46296 14436
rect 46348 14424 46354 14476
rect 46474 14464 46480 14476
rect 46435 14436 46480 14464
rect 46474 14424 46480 14436
rect 46532 14424 46538 14476
rect 48130 14464 48136 14476
rect 48091 14436 48136 14464
rect 48130 14424 48136 14436
rect 48188 14424 48194 14476
rect 19889 14399 19947 14405
rect 19889 14396 19901 14399
rect 18524 14368 19901 14396
rect 19889 14365 19901 14368
rect 19935 14365 19947 14399
rect 25222 14396 25228 14408
rect 25183 14368 25228 14396
rect 19889 14359 19947 14365
rect 25222 14356 25228 14368
rect 25280 14356 25286 14408
rect 25685 14399 25743 14405
rect 25685 14365 25697 14399
rect 25731 14396 25743 14399
rect 25774 14396 25780 14408
rect 25731 14368 25780 14396
rect 25731 14365 25743 14368
rect 25685 14359 25743 14365
rect 25774 14356 25780 14368
rect 25832 14396 25838 14408
rect 26970 14396 26976 14408
rect 25832 14368 26004 14396
rect 26931 14368 26976 14396
rect 25832 14356 25838 14368
rect 12158 14288 12164 14340
rect 12216 14328 12222 14340
rect 18601 14331 18659 14337
rect 18601 14328 18613 14331
rect 12216 14300 18613 14328
rect 12216 14288 12222 14300
rect 18601 14297 18613 14300
rect 18647 14297 18659 14331
rect 18601 14291 18659 14297
rect 2222 14220 2228 14272
rect 2280 14260 2286 14272
rect 2501 14263 2559 14269
rect 2501 14260 2513 14263
rect 2280 14232 2513 14260
rect 2280 14220 2286 14232
rect 2501 14229 2513 14232
rect 2547 14229 2559 14263
rect 18616 14260 18644 14291
rect 24578 14260 24584 14272
rect 18616 14232 24584 14260
rect 2501 14223 2559 14229
rect 24578 14220 24584 14232
rect 24636 14220 24642 14272
rect 25976 14260 26004 14368
rect 26970 14356 26976 14368
rect 27028 14356 27034 14408
rect 27249 14399 27307 14405
rect 27249 14365 27261 14399
rect 27295 14396 27307 14399
rect 31386 14396 31392 14408
rect 27295 14368 28028 14396
rect 31347 14368 31392 14396
rect 27295 14365 27307 14368
rect 27249 14359 27307 14365
rect 28000 14340 28028 14368
rect 31386 14356 31392 14368
rect 31444 14356 31450 14408
rect 31662 14396 31668 14408
rect 31623 14368 31668 14396
rect 31662 14356 31668 14368
rect 31720 14356 31726 14408
rect 45186 14356 45192 14408
rect 45244 14396 45250 14408
rect 45649 14399 45707 14405
rect 45649 14396 45661 14399
rect 45244 14368 45661 14396
rect 45244 14356 45250 14368
rect 45649 14365 45661 14368
rect 45695 14365 45707 14399
rect 45649 14359 45707 14365
rect 27798 14328 27804 14340
rect 27759 14300 27804 14328
rect 27798 14288 27804 14300
rect 27856 14288 27862 14340
rect 27982 14328 27988 14340
rect 27943 14300 27988 14328
rect 27982 14288 27988 14300
rect 28040 14288 28046 14340
rect 31404 14328 31432 14356
rect 33226 14328 33232 14340
rect 31404 14300 33232 14328
rect 33226 14288 33232 14300
rect 33284 14288 33290 14340
rect 35986 14260 35992 14272
rect 25976 14232 35992 14260
rect 35986 14220 35992 14232
rect 36044 14220 36050 14272
rect 1104 14170 48852 14192
rect 1104 14118 16880 14170
rect 16932 14118 16944 14170
rect 16996 14118 17008 14170
rect 17060 14118 17072 14170
rect 17124 14118 17136 14170
rect 17188 14118 32811 14170
rect 32863 14118 32875 14170
rect 32927 14118 32939 14170
rect 32991 14118 33003 14170
rect 33055 14118 33067 14170
rect 33119 14118 48852 14170
rect 1104 14096 48852 14118
rect 2222 13988 2228 14000
rect 2183 13960 2228 13988
rect 2222 13948 2228 13960
rect 2280 13948 2286 14000
rect 27890 13948 27896 14000
rect 27948 13988 27954 14000
rect 28169 13991 28227 13997
rect 28169 13988 28181 13991
rect 27948 13960 28181 13988
rect 27948 13948 27954 13960
rect 28169 13957 28181 13960
rect 28215 13988 28227 13991
rect 45373 13991 45431 13997
rect 28215 13960 31754 13988
rect 28215 13957 28227 13960
rect 28169 13951 28227 13957
rect 2038 13920 2044 13932
rect 1999 13892 2044 13920
rect 2038 13880 2044 13892
rect 2096 13880 2102 13932
rect 25222 13920 25228 13932
rect 25183 13892 25228 13920
rect 25222 13880 25228 13892
rect 25280 13880 25286 13932
rect 27341 13923 27399 13929
rect 27341 13889 27353 13923
rect 27387 13920 27399 13923
rect 27982 13920 27988 13932
rect 27387 13892 27988 13920
rect 27387 13889 27399 13892
rect 27341 13883 27399 13889
rect 27982 13880 27988 13892
rect 28040 13920 28046 13932
rect 28721 13923 28779 13929
rect 28721 13920 28733 13923
rect 28040 13892 28733 13920
rect 28040 13880 28046 13892
rect 28721 13889 28733 13892
rect 28767 13889 28779 13923
rect 30006 13920 30012 13932
rect 28721 13883 28779 13889
rect 28828 13892 30012 13920
rect 2774 13812 2780 13864
rect 2832 13852 2838 13864
rect 2832 13824 2877 13852
rect 2832 13812 2838 13824
rect 10226 13812 10232 13864
rect 10284 13852 10290 13864
rect 25501 13855 25559 13861
rect 25501 13852 25513 13855
rect 10284 13824 25513 13852
rect 10284 13812 10290 13824
rect 25501 13821 25513 13824
rect 25547 13852 25559 13855
rect 28828 13852 28856 13892
rect 30006 13880 30012 13892
rect 30064 13880 30070 13932
rect 31726 13920 31754 13960
rect 45373 13957 45385 13991
rect 45419 13988 45431 13991
rect 47673 13991 47731 13997
rect 47673 13988 47685 13991
rect 45419 13960 47685 13988
rect 45419 13957 45431 13960
rect 45373 13951 45431 13957
rect 47673 13957 47685 13960
rect 47719 13957 47731 13991
rect 47673 13951 47731 13957
rect 34698 13920 34704 13932
rect 31726 13892 34704 13920
rect 34698 13880 34704 13892
rect 34756 13880 34762 13932
rect 45186 13920 45192 13932
rect 45147 13892 45192 13920
rect 45186 13880 45192 13892
rect 45244 13880 45250 13932
rect 47026 13880 47032 13932
rect 47084 13920 47090 13932
rect 47581 13923 47639 13929
rect 47581 13920 47593 13923
rect 47084 13892 47593 13920
rect 47084 13880 47090 13892
rect 47581 13889 47593 13892
rect 47627 13889 47639 13923
rect 47581 13883 47639 13889
rect 25547 13824 28856 13852
rect 25547 13821 25559 13824
rect 25501 13815 25559 13821
rect 28994 13812 29000 13864
rect 29052 13852 29058 13864
rect 31386 13852 31392 13864
rect 29052 13824 31392 13852
rect 29052 13812 29058 13824
rect 31386 13812 31392 13824
rect 31444 13812 31450 13864
rect 46842 13852 46848 13864
rect 46803 13824 46848 13852
rect 46842 13812 46848 13824
rect 46900 13812 46906 13864
rect 1104 13626 48852 13648
rect 1104 13574 8915 13626
rect 8967 13574 8979 13626
rect 9031 13574 9043 13626
rect 9095 13574 9107 13626
rect 9159 13574 9171 13626
rect 9223 13574 24846 13626
rect 24898 13574 24910 13626
rect 24962 13574 24974 13626
rect 25026 13574 25038 13626
rect 25090 13574 25102 13626
rect 25154 13574 40776 13626
rect 40828 13574 40840 13626
rect 40892 13574 40904 13626
rect 40956 13574 40968 13626
rect 41020 13574 41032 13626
rect 41084 13574 48852 13626
rect 1104 13552 48852 13574
rect 26786 13336 26792 13388
rect 26844 13376 26850 13388
rect 27157 13379 27215 13385
rect 27157 13376 27169 13379
rect 26844 13348 27169 13376
rect 26844 13336 26850 13348
rect 27157 13345 27169 13348
rect 27203 13376 27215 13379
rect 27430 13376 27436 13388
rect 27203 13348 27436 13376
rect 27203 13345 27215 13348
rect 27157 13339 27215 13345
rect 27430 13336 27436 13348
rect 27488 13336 27494 13388
rect 45189 13379 45247 13385
rect 45189 13345 45201 13379
rect 45235 13376 45247 13379
rect 46293 13379 46351 13385
rect 46293 13376 46305 13379
rect 45235 13348 46305 13376
rect 45235 13345 45247 13348
rect 45189 13339 45247 13345
rect 46293 13345 46305 13348
rect 46339 13345 46351 13379
rect 46293 13339 46351 13345
rect 2038 13268 2044 13320
rect 2096 13308 2102 13320
rect 2133 13311 2191 13317
rect 2133 13308 2145 13311
rect 2096 13280 2145 13308
rect 2096 13268 2102 13280
rect 2133 13277 2145 13280
rect 2179 13277 2191 13311
rect 3786 13308 3792 13320
rect 3747 13280 3792 13308
rect 2133 13271 2191 13277
rect 3786 13268 3792 13280
rect 3844 13268 3850 13320
rect 26881 13311 26939 13317
rect 26881 13277 26893 13311
rect 26927 13308 26939 13311
rect 27614 13308 27620 13320
rect 26927 13280 27620 13308
rect 26927 13277 26939 13280
rect 26881 13271 26939 13277
rect 27614 13268 27620 13280
rect 27672 13308 27678 13320
rect 27982 13308 27988 13320
rect 27672 13280 27988 13308
rect 27672 13268 27678 13280
rect 27982 13268 27988 13280
rect 28040 13268 28046 13320
rect 45649 13311 45707 13317
rect 45649 13277 45661 13311
rect 45695 13277 45707 13311
rect 45649 13271 45707 13277
rect 27430 13200 27436 13252
rect 27488 13240 27494 13252
rect 27488 13212 35894 13240
rect 27488 13200 27494 13212
rect 35866 13172 35894 13212
rect 36538 13172 36544 13184
rect 35866 13144 36544 13172
rect 36538 13132 36544 13144
rect 36596 13172 36602 13184
rect 37366 13172 37372 13184
rect 36596 13144 37372 13172
rect 36596 13132 36602 13144
rect 37366 13132 37372 13144
rect 37424 13132 37430 13184
rect 45664 13172 45692 13271
rect 45741 13243 45799 13249
rect 45741 13209 45753 13243
rect 45787 13240 45799 13243
rect 46477 13243 46535 13249
rect 46477 13240 46489 13243
rect 45787 13212 46489 13240
rect 45787 13209 45799 13212
rect 45741 13203 45799 13209
rect 46477 13209 46489 13212
rect 46523 13209 46535 13243
rect 48130 13240 48136 13252
rect 48091 13212 48136 13240
rect 46477 13203 46535 13209
rect 48130 13200 48136 13212
rect 48188 13200 48194 13252
rect 46934 13172 46940 13184
rect 45664 13144 46940 13172
rect 46934 13132 46940 13144
rect 46992 13132 46998 13184
rect 1104 13082 48852 13104
rect 1104 13030 16880 13082
rect 16932 13030 16944 13082
rect 16996 13030 17008 13082
rect 17060 13030 17072 13082
rect 17124 13030 17136 13082
rect 17188 13030 32811 13082
rect 32863 13030 32875 13082
rect 32927 13030 32939 13082
rect 32991 13030 33003 13082
rect 33055 13030 33067 13082
rect 33119 13030 48852 13082
rect 1104 13008 48852 13030
rect 45373 12903 45431 12909
rect 45373 12869 45385 12903
rect 45419 12900 45431 12903
rect 47673 12903 47731 12909
rect 47673 12900 47685 12903
rect 45419 12872 47685 12900
rect 45419 12869 45431 12872
rect 45373 12863 45431 12869
rect 47673 12869 47685 12872
rect 47719 12869 47731 12903
rect 47673 12863 47731 12869
rect 2038 12832 2044 12844
rect 1999 12804 2044 12832
rect 2038 12792 2044 12804
rect 2096 12792 2102 12844
rect 27614 12832 27620 12844
rect 27575 12804 27620 12832
rect 27614 12792 27620 12804
rect 27672 12792 27678 12844
rect 47486 12792 47492 12844
rect 47544 12832 47550 12844
rect 47581 12835 47639 12841
rect 47581 12832 47593 12835
rect 47544 12804 47593 12832
rect 47544 12792 47550 12804
rect 47581 12801 47593 12804
rect 47627 12801 47639 12835
rect 47581 12795 47639 12801
rect 2222 12764 2228 12776
rect 2183 12736 2228 12764
rect 2222 12724 2228 12736
rect 2280 12724 2286 12776
rect 2774 12724 2780 12776
rect 2832 12764 2838 12776
rect 27338 12764 27344 12776
rect 2832 12736 2877 12764
rect 27251 12736 27344 12764
rect 2832 12724 2838 12736
rect 27338 12724 27344 12736
rect 27396 12764 27402 12776
rect 42334 12764 42340 12776
rect 27396 12736 42340 12764
rect 27396 12724 27402 12736
rect 42334 12724 42340 12736
rect 42392 12724 42398 12776
rect 45186 12764 45192 12776
rect 45147 12736 45192 12764
rect 45186 12724 45192 12736
rect 45244 12724 45250 12776
rect 46842 12764 46848 12776
rect 46803 12736 46848 12764
rect 46842 12724 46848 12736
rect 46900 12724 46906 12776
rect 32674 12656 32680 12708
rect 32732 12696 32738 12708
rect 47486 12696 47492 12708
rect 32732 12668 47492 12696
rect 32732 12656 32738 12668
rect 47486 12656 47492 12668
rect 47544 12656 47550 12708
rect 1104 12538 48852 12560
rect 1104 12486 8915 12538
rect 8967 12486 8979 12538
rect 9031 12486 9043 12538
rect 9095 12486 9107 12538
rect 9159 12486 9171 12538
rect 9223 12486 24846 12538
rect 24898 12486 24910 12538
rect 24962 12486 24974 12538
rect 25026 12486 25038 12538
rect 25090 12486 25102 12538
rect 25154 12486 40776 12538
rect 40828 12486 40840 12538
rect 40892 12486 40904 12538
rect 40956 12486 40968 12538
rect 41020 12486 41032 12538
rect 41084 12486 48852 12538
rect 1104 12464 48852 12486
rect 2222 12384 2228 12436
rect 2280 12424 2286 12436
rect 2501 12427 2559 12433
rect 2501 12424 2513 12427
rect 2280 12396 2513 12424
rect 2280 12384 2286 12396
rect 2501 12393 2513 12396
rect 2547 12393 2559 12427
rect 2501 12387 2559 12393
rect 44453 12427 44511 12433
rect 44453 12393 44465 12427
rect 44499 12424 44511 12427
rect 45186 12424 45192 12436
rect 44499 12396 45192 12424
rect 44499 12393 44511 12396
rect 44453 12387 44511 12393
rect 45186 12384 45192 12396
rect 45244 12384 45250 12436
rect 3786 12288 3792 12300
rect 3747 12260 3792 12288
rect 3786 12248 3792 12260
rect 3844 12248 3850 12300
rect 4062 12248 4068 12300
rect 4120 12288 4126 12300
rect 4249 12291 4307 12297
rect 4249 12288 4261 12291
rect 4120 12260 4261 12288
rect 4120 12248 4126 12260
rect 4249 12257 4261 12260
rect 4295 12257 4307 12291
rect 47578 12288 47584 12300
rect 47539 12260 47584 12288
rect 4249 12251 4307 12257
rect 47578 12248 47584 12260
rect 47636 12248 47642 12300
rect 2590 12220 2596 12232
rect 2551 12192 2596 12220
rect 2590 12180 2596 12192
rect 2648 12180 2654 12232
rect 45465 12223 45523 12229
rect 45465 12189 45477 12223
rect 45511 12220 45523 12223
rect 45925 12223 45983 12229
rect 45925 12220 45937 12223
rect 45511 12192 45937 12220
rect 45511 12189 45523 12192
rect 45465 12183 45523 12189
rect 45925 12189 45937 12192
rect 45971 12189 45983 12223
rect 45925 12183 45983 12189
rect 3970 12152 3976 12164
rect 3931 12124 3976 12152
rect 3970 12112 3976 12124
rect 4028 12112 4034 12164
rect 46109 12155 46167 12161
rect 46109 12121 46121 12155
rect 46155 12152 46167 12155
rect 47670 12152 47676 12164
rect 46155 12124 47676 12152
rect 46155 12121 46167 12124
rect 46109 12115 46167 12121
rect 47670 12112 47676 12124
rect 47728 12112 47734 12164
rect 1104 11994 48852 12016
rect 1104 11942 16880 11994
rect 16932 11942 16944 11994
rect 16996 11942 17008 11994
rect 17060 11942 17072 11994
rect 17124 11942 17136 11994
rect 17188 11942 32811 11994
rect 32863 11942 32875 11994
rect 32927 11942 32939 11994
rect 32991 11942 33003 11994
rect 33055 11942 33067 11994
rect 33119 11942 48852 11994
rect 1104 11920 48852 11942
rect 3881 11883 3939 11889
rect 3881 11849 3893 11883
rect 3927 11880 3939 11883
rect 3970 11880 3976 11892
rect 3927 11852 3976 11880
rect 3927 11849 3939 11852
rect 3881 11843 3939 11849
rect 3970 11840 3976 11852
rect 4028 11840 4034 11892
rect 47670 11880 47676 11892
rect 47631 11852 47676 11880
rect 47670 11840 47676 11852
rect 47728 11840 47734 11892
rect 3973 11747 4031 11753
rect 3973 11713 3985 11747
rect 4019 11744 4031 11747
rect 8202 11744 8208 11756
rect 4019 11716 8208 11744
rect 4019 11713 4031 11716
rect 3973 11707 4031 11713
rect 8202 11704 8208 11716
rect 8260 11744 8266 11756
rect 27338 11744 27344 11756
rect 8260 11716 27344 11744
rect 8260 11704 8266 11716
rect 27338 11704 27344 11716
rect 27396 11704 27402 11756
rect 47394 11704 47400 11756
rect 47452 11744 47458 11756
rect 47581 11747 47639 11753
rect 47581 11744 47593 11747
rect 47452 11716 47593 11744
rect 47452 11704 47458 11716
rect 47581 11713 47593 11716
rect 47627 11713 47639 11747
rect 47581 11707 47639 11713
rect 44729 11679 44787 11685
rect 44729 11645 44741 11679
rect 44775 11676 44787 11679
rect 45189 11679 45247 11685
rect 45189 11676 45201 11679
rect 44775 11648 45201 11676
rect 44775 11645 44787 11648
rect 44729 11639 44787 11645
rect 45189 11645 45201 11648
rect 45235 11645 45247 11679
rect 45189 11639 45247 11645
rect 45373 11679 45431 11685
rect 45373 11645 45385 11679
rect 45419 11676 45431 11679
rect 46566 11676 46572 11688
rect 45419 11648 46572 11676
rect 45419 11645 45431 11648
rect 45373 11639 45431 11645
rect 46566 11636 46572 11648
rect 46624 11636 46630 11688
rect 46842 11676 46848 11688
rect 46803 11648 46848 11676
rect 46842 11636 46848 11648
rect 46900 11636 46906 11688
rect 1104 11450 48852 11472
rect 1104 11398 8915 11450
rect 8967 11398 8979 11450
rect 9031 11398 9043 11450
rect 9095 11398 9107 11450
rect 9159 11398 9171 11450
rect 9223 11398 24846 11450
rect 24898 11398 24910 11450
rect 24962 11398 24974 11450
rect 25026 11398 25038 11450
rect 25090 11398 25102 11450
rect 25154 11398 40776 11450
rect 40828 11398 40840 11450
rect 40892 11398 40904 11450
rect 40956 11398 40968 11450
rect 41020 11398 41032 11450
rect 41084 11398 48852 11450
rect 1104 11376 48852 11398
rect 2038 11092 2044 11144
rect 2096 11132 2102 11144
rect 2133 11135 2191 11141
rect 2133 11132 2145 11135
rect 2096 11104 2145 11132
rect 2096 11092 2102 11104
rect 2133 11101 2145 11104
rect 2179 11101 2191 11135
rect 2133 11095 2191 11101
rect 45833 11135 45891 11141
rect 45833 11101 45845 11135
rect 45879 11132 45891 11135
rect 46293 11135 46351 11141
rect 46293 11132 46305 11135
rect 45879 11104 46305 11132
rect 45879 11101 45891 11104
rect 45833 11095 45891 11101
rect 46293 11101 46305 11104
rect 46339 11101 46351 11135
rect 46293 11095 46351 11101
rect 46477 11067 46535 11073
rect 46477 11033 46489 11067
rect 46523 11064 46535 11067
rect 47670 11064 47676 11076
rect 46523 11036 47676 11064
rect 46523 11033 46535 11036
rect 46477 11027 46535 11033
rect 47670 11024 47676 11036
rect 47728 11024 47734 11076
rect 48130 11064 48136 11076
rect 48091 11036 48136 11064
rect 48130 11024 48136 11036
rect 48188 11024 48194 11076
rect 1104 10906 48852 10928
rect 1104 10854 16880 10906
rect 16932 10854 16944 10906
rect 16996 10854 17008 10906
rect 17060 10854 17072 10906
rect 17124 10854 17136 10906
rect 17188 10854 32811 10906
rect 32863 10854 32875 10906
rect 32927 10854 32939 10906
rect 32991 10854 33003 10906
rect 33055 10854 33067 10906
rect 33119 10854 48852 10906
rect 1104 10832 48852 10854
rect 46566 10792 46572 10804
rect 46527 10764 46572 10792
rect 46566 10752 46572 10764
rect 46624 10752 46630 10804
rect 47670 10792 47676 10804
rect 47631 10764 47676 10792
rect 47670 10752 47676 10764
rect 47728 10752 47734 10804
rect 2038 10656 2044 10668
rect 1999 10628 2044 10656
rect 2038 10616 2044 10628
rect 2096 10616 2102 10668
rect 46658 10656 46664 10668
rect 46571 10628 46664 10656
rect 46658 10616 46664 10628
rect 46716 10656 46722 10668
rect 47026 10656 47032 10668
rect 46716 10628 47032 10656
rect 46716 10616 46722 10628
rect 47026 10616 47032 10628
rect 47084 10616 47090 10668
rect 47394 10616 47400 10668
rect 47452 10656 47458 10668
rect 47581 10659 47639 10665
rect 47581 10656 47593 10659
rect 47452 10628 47593 10656
rect 47452 10616 47458 10628
rect 47581 10625 47593 10628
rect 47627 10625 47639 10659
rect 47581 10619 47639 10625
rect 2225 10591 2283 10597
rect 2225 10557 2237 10591
rect 2271 10588 2283 10591
rect 2498 10588 2504 10600
rect 2271 10560 2504 10588
rect 2271 10557 2283 10560
rect 2225 10551 2283 10557
rect 2498 10548 2504 10560
rect 2556 10548 2562 10600
rect 2774 10588 2780 10600
rect 2735 10560 2780 10588
rect 2774 10548 2780 10560
rect 2832 10548 2838 10600
rect 11054 10412 11060 10464
rect 11112 10452 11118 10464
rect 11517 10455 11575 10461
rect 11517 10452 11529 10455
rect 11112 10424 11529 10452
rect 11112 10412 11118 10424
rect 11517 10421 11529 10424
rect 11563 10421 11575 10455
rect 12986 10452 12992 10464
rect 12947 10424 12992 10452
rect 11517 10415 11575 10421
rect 12986 10412 12992 10424
rect 13044 10412 13050 10464
rect 46017 10455 46075 10461
rect 46017 10421 46029 10455
rect 46063 10452 46075 10455
rect 46290 10452 46296 10464
rect 46063 10424 46296 10452
rect 46063 10421 46075 10424
rect 46017 10415 46075 10421
rect 46290 10412 46296 10424
rect 46348 10412 46354 10464
rect 1104 10362 48852 10384
rect 1104 10310 8915 10362
rect 8967 10310 8979 10362
rect 9031 10310 9043 10362
rect 9095 10310 9107 10362
rect 9159 10310 9171 10362
rect 9223 10310 24846 10362
rect 24898 10310 24910 10362
rect 24962 10310 24974 10362
rect 25026 10310 25038 10362
rect 25090 10310 25102 10362
rect 25154 10310 40776 10362
rect 40828 10310 40840 10362
rect 40892 10310 40904 10362
rect 40956 10310 40968 10362
rect 41020 10310 41032 10362
rect 41084 10310 48852 10362
rect 1104 10288 48852 10310
rect 2498 10248 2504 10260
rect 2459 10220 2504 10248
rect 2498 10208 2504 10220
rect 2556 10208 2562 10260
rect 6886 10152 11560 10180
rect 2593 10047 2651 10053
rect 2593 10013 2605 10047
rect 2639 10044 2651 10047
rect 2682 10044 2688 10056
rect 2639 10016 2688 10044
rect 2639 10013 2651 10016
rect 2593 10007 2651 10013
rect 2682 10004 2688 10016
rect 2740 10004 2746 10056
rect 3418 9936 3424 9988
rect 3476 9976 3482 9988
rect 6886 9976 6914 10152
rect 11054 10112 11060 10124
rect 11015 10084 11060 10112
rect 11054 10072 11060 10084
rect 11112 10072 11118 10124
rect 11532 10121 11560 10152
rect 11517 10115 11575 10121
rect 11517 10081 11529 10115
rect 11563 10081 11575 10115
rect 46290 10112 46296 10124
rect 46251 10084 46296 10112
rect 11517 10075 11575 10081
rect 46290 10072 46296 10084
rect 46348 10072 46354 10124
rect 48130 10112 48136 10124
rect 48091 10084 48136 10112
rect 48130 10072 48136 10084
rect 48188 10072 48194 10124
rect 13541 10047 13599 10053
rect 13541 10013 13553 10047
rect 13587 10044 13599 10047
rect 18322 10044 18328 10056
rect 13587 10016 18328 10044
rect 13587 10013 13599 10016
rect 13541 10007 13599 10013
rect 18322 10004 18328 10016
rect 18380 10004 18386 10056
rect 40034 10044 40040 10056
rect 39995 10016 40040 10044
rect 40034 10004 40040 10016
rect 40092 10004 40098 10056
rect 11238 9976 11244 9988
rect 3476 9948 6914 9976
rect 11199 9948 11244 9976
rect 3476 9936 3482 9948
rect 11238 9936 11244 9948
rect 11296 9936 11302 9988
rect 46477 9979 46535 9985
rect 46477 9945 46489 9979
rect 46523 9976 46535 9979
rect 47670 9976 47676 9988
rect 46523 9948 47676 9976
rect 46523 9945 46535 9948
rect 46477 9939 46535 9945
rect 47670 9936 47676 9948
rect 47728 9936 47734 9988
rect 13170 9868 13176 9920
rect 13228 9908 13234 9920
rect 13449 9911 13507 9917
rect 13449 9908 13461 9911
rect 13228 9880 13461 9908
rect 13228 9868 13234 9880
rect 13449 9877 13461 9880
rect 13495 9877 13507 9911
rect 13449 9871 13507 9877
rect 1104 9818 48852 9840
rect 1104 9766 16880 9818
rect 16932 9766 16944 9818
rect 16996 9766 17008 9818
rect 17060 9766 17072 9818
rect 17124 9766 17136 9818
rect 17188 9766 32811 9818
rect 32863 9766 32875 9818
rect 32927 9766 32939 9818
rect 32991 9766 33003 9818
rect 33055 9766 33067 9818
rect 33119 9766 48852 9818
rect 1104 9744 48852 9766
rect 11238 9664 11244 9716
rect 11296 9704 11302 9716
rect 11609 9707 11667 9713
rect 11609 9704 11621 9707
rect 11296 9676 11621 9704
rect 11296 9664 11302 9676
rect 11609 9673 11621 9676
rect 11655 9673 11667 9707
rect 11609 9667 11667 9673
rect 13170 9636 13176 9648
rect 13131 9608 13176 9636
rect 13170 9596 13176 9608
rect 13228 9596 13234 9648
rect 25314 9596 25320 9648
rect 25372 9636 25378 9648
rect 47670 9636 47676 9648
rect 25372 9608 45554 9636
rect 47631 9608 47676 9636
rect 25372 9596 25378 9608
rect 11701 9571 11759 9577
rect 11701 9537 11713 9571
rect 11747 9568 11759 9571
rect 11790 9568 11796 9580
rect 11747 9540 11796 9568
rect 11747 9537 11759 9540
rect 11701 9531 11759 9537
rect 11790 9528 11796 9540
rect 11848 9528 11854 9580
rect 12986 9568 12992 9580
rect 12947 9540 12992 9568
rect 12986 9528 12992 9540
rect 13044 9528 13050 9580
rect 40034 9568 40040 9580
rect 39995 9540 40040 9568
rect 40034 9528 40040 9540
rect 40092 9528 40098 9580
rect 45526 9568 45554 9608
rect 47670 9596 47676 9608
rect 47728 9596 47734 9648
rect 47578 9568 47584 9580
rect 45526 9540 47584 9568
rect 47578 9528 47584 9540
rect 47636 9528 47642 9580
rect 13538 9500 13544 9512
rect 13499 9472 13544 9500
rect 13538 9460 13544 9472
rect 13596 9460 13602 9512
rect 40218 9500 40224 9512
rect 40179 9472 40224 9500
rect 40218 9460 40224 9472
rect 40276 9460 40282 9512
rect 40586 9500 40592 9512
rect 40547 9472 40592 9500
rect 40586 9460 40592 9472
rect 40644 9460 40650 9512
rect 1104 9274 48852 9296
rect 1104 9222 8915 9274
rect 8967 9222 8979 9274
rect 9031 9222 9043 9274
rect 9095 9222 9107 9274
rect 9159 9222 9171 9274
rect 9223 9222 24846 9274
rect 24898 9222 24910 9274
rect 24962 9222 24974 9274
rect 25026 9222 25038 9274
rect 25090 9222 25102 9274
rect 25154 9222 40776 9274
rect 40828 9222 40840 9274
rect 40892 9222 40904 9274
rect 40956 9222 40968 9274
rect 41020 9222 41032 9274
rect 41084 9222 48852 9274
rect 1104 9200 48852 9222
rect 40129 9163 40187 9169
rect 40129 9129 40141 9163
rect 40175 9160 40187 9163
rect 40218 9160 40224 9172
rect 40175 9132 40224 9160
rect 40175 9129 40187 9132
rect 40129 9123 40187 9129
rect 40218 9120 40224 9132
rect 40276 9120 40282 9172
rect 2038 8956 2044 8968
rect 1999 8928 2044 8956
rect 2038 8916 2044 8928
rect 2096 8916 2102 8968
rect 20622 8916 20628 8968
rect 20680 8956 20686 8968
rect 40037 8959 40095 8965
rect 40037 8956 40049 8959
rect 20680 8928 40049 8956
rect 20680 8916 20686 8928
rect 40037 8925 40049 8928
rect 40083 8956 40095 8959
rect 46658 8956 46664 8968
rect 40083 8928 46664 8956
rect 40083 8925 40095 8928
rect 40037 8919 40095 8925
rect 46658 8916 46664 8928
rect 46716 8916 46722 8968
rect 1104 8730 48852 8752
rect 1104 8678 16880 8730
rect 16932 8678 16944 8730
rect 16996 8678 17008 8730
rect 17060 8678 17072 8730
rect 17124 8678 17136 8730
rect 17188 8678 32811 8730
rect 32863 8678 32875 8730
rect 32927 8678 32939 8730
rect 32991 8678 33003 8730
rect 33055 8678 33067 8730
rect 33119 8678 48852 8730
rect 1104 8656 48852 8678
rect 2038 8480 2044 8492
rect 1999 8452 2044 8480
rect 2038 8440 2044 8452
rect 2096 8440 2102 8492
rect 2222 8412 2228 8424
rect 2183 8384 2228 8412
rect 2222 8372 2228 8384
rect 2280 8372 2286 8424
rect 2774 8412 2780 8424
rect 2735 8384 2780 8412
rect 2774 8372 2780 8384
rect 2832 8372 2838 8424
rect 10318 8236 10324 8288
rect 10376 8276 10382 8288
rect 10413 8279 10471 8285
rect 10413 8276 10425 8279
rect 10376 8248 10425 8276
rect 10376 8236 10382 8248
rect 10413 8245 10425 8248
rect 10459 8245 10471 8279
rect 10413 8239 10471 8245
rect 1104 8186 48852 8208
rect 1104 8134 8915 8186
rect 8967 8134 8979 8186
rect 9031 8134 9043 8186
rect 9095 8134 9107 8186
rect 9159 8134 9171 8186
rect 9223 8134 24846 8186
rect 24898 8134 24910 8186
rect 24962 8134 24974 8186
rect 25026 8134 25038 8186
rect 25090 8134 25102 8186
rect 25154 8134 40776 8186
rect 40828 8134 40840 8186
rect 40892 8134 40904 8186
rect 40956 8134 40968 8186
rect 41020 8134 41032 8186
rect 41084 8134 48852 8186
rect 1104 8112 48852 8134
rect 2222 8032 2228 8084
rect 2280 8072 2286 8084
rect 2317 8075 2375 8081
rect 2317 8072 2329 8075
rect 2280 8044 2329 8072
rect 2280 8032 2286 8044
rect 2317 8041 2329 8044
rect 2363 8041 2375 8075
rect 2317 8035 2375 8041
rect 10318 7936 10324 7948
rect 10279 7908 10324 7936
rect 10318 7896 10324 7908
rect 10376 7896 10382 7948
rect 10962 7936 10968 7948
rect 10923 7908 10968 7936
rect 10962 7896 10968 7908
rect 11020 7896 11026 7948
rect 2406 7868 2412 7880
rect 2367 7840 2412 7868
rect 2406 7828 2412 7840
rect 2464 7828 2470 7880
rect 17678 7868 17684 7880
rect 17639 7840 17684 7868
rect 17678 7828 17684 7840
rect 17736 7828 17742 7880
rect 29730 7828 29736 7880
rect 29788 7868 29794 7880
rect 29825 7871 29883 7877
rect 29825 7868 29837 7871
rect 29788 7840 29837 7868
rect 29788 7828 29794 7840
rect 29825 7837 29837 7840
rect 29871 7837 29883 7871
rect 33226 7868 33232 7880
rect 33187 7840 33232 7868
rect 29825 7831 29883 7837
rect 33226 7828 33232 7840
rect 33284 7828 33290 7880
rect 10502 7800 10508 7812
rect 10463 7772 10508 7800
rect 10502 7760 10508 7772
rect 10560 7760 10566 7812
rect 33321 7735 33379 7741
rect 33321 7701 33333 7735
rect 33367 7732 33379 7735
rect 33870 7732 33876 7744
rect 33367 7704 33876 7732
rect 33367 7701 33379 7704
rect 33321 7695 33379 7701
rect 33870 7692 33876 7704
rect 33928 7692 33934 7744
rect 1104 7642 48852 7664
rect 1104 7590 16880 7642
rect 16932 7590 16944 7642
rect 16996 7590 17008 7642
rect 17060 7590 17072 7642
rect 17124 7590 17136 7642
rect 17188 7590 32811 7642
rect 32863 7590 32875 7642
rect 32927 7590 32939 7642
rect 32991 7590 33003 7642
rect 33055 7590 33067 7642
rect 33119 7590 48852 7642
rect 1104 7568 48852 7590
rect 10502 7528 10508 7540
rect 10463 7500 10508 7528
rect 10502 7488 10508 7500
rect 10560 7488 10566 7540
rect 33870 7460 33876 7472
rect 33831 7432 33876 7460
rect 33870 7420 33876 7432
rect 33928 7420 33934 7472
rect 10410 7392 10416 7404
rect 10371 7364 10416 7392
rect 10410 7352 10416 7364
rect 10468 7352 10474 7404
rect 17678 7392 17684 7404
rect 17639 7364 17684 7392
rect 17678 7352 17684 7364
rect 17736 7352 17742 7404
rect 29086 7392 29092 7404
rect 29047 7364 29092 7392
rect 29086 7352 29092 7364
rect 29144 7352 29150 7404
rect 29730 7392 29736 7404
rect 29691 7364 29736 7392
rect 29730 7352 29736 7364
rect 29788 7352 29794 7404
rect 17865 7327 17923 7333
rect 17865 7293 17877 7327
rect 17911 7324 17923 7327
rect 18046 7324 18052 7336
rect 17911 7296 18052 7324
rect 17911 7293 17923 7296
rect 17865 7287 17923 7293
rect 18046 7284 18052 7296
rect 18104 7284 18110 7336
rect 18141 7327 18199 7333
rect 18141 7293 18153 7327
rect 18187 7293 18199 7327
rect 18141 7287 18199 7293
rect 29181 7327 29239 7333
rect 29181 7293 29193 7327
rect 29227 7324 29239 7327
rect 29917 7327 29975 7333
rect 29917 7324 29929 7327
rect 29227 7296 29929 7324
rect 29227 7293 29239 7296
rect 29181 7287 29239 7293
rect 29917 7293 29929 7296
rect 29963 7293 29975 7327
rect 29917 7287 29975 7293
rect 31573 7327 31631 7333
rect 31573 7293 31585 7327
rect 31619 7293 31631 7327
rect 33686 7324 33692 7336
rect 33647 7296 33692 7324
rect 31573 7287 31631 7293
rect 3418 7216 3424 7268
rect 3476 7256 3482 7268
rect 18156 7256 18184 7287
rect 3476 7228 18184 7256
rect 31588 7256 31616 7287
rect 33686 7284 33692 7296
rect 33744 7284 33750 7336
rect 34606 7324 34612 7336
rect 34567 7296 34612 7324
rect 34606 7284 34612 7296
rect 34664 7284 34670 7336
rect 46750 7324 46756 7336
rect 35866 7296 46756 7324
rect 35866 7256 35894 7296
rect 46750 7284 46756 7296
rect 46808 7284 46814 7336
rect 31588 7228 35894 7256
rect 3476 7216 3482 7228
rect 2130 7148 2136 7200
rect 2188 7188 2194 7200
rect 2225 7191 2283 7197
rect 2225 7188 2237 7191
rect 2188 7160 2237 7188
rect 2188 7148 2194 7160
rect 2225 7157 2237 7160
rect 2271 7157 2283 7191
rect 2225 7151 2283 7157
rect 1104 7098 48852 7120
rect 1104 7046 8915 7098
rect 8967 7046 8979 7098
rect 9031 7046 9043 7098
rect 9095 7046 9107 7098
rect 9159 7046 9171 7098
rect 9223 7046 24846 7098
rect 24898 7046 24910 7098
rect 24962 7046 24974 7098
rect 25026 7046 25038 7098
rect 25090 7046 25102 7098
rect 25154 7046 40776 7098
rect 40828 7046 40840 7098
rect 40892 7046 40904 7098
rect 40956 7046 40968 7098
rect 41020 7046 41032 7098
rect 41084 7046 48852 7098
rect 1104 7024 48852 7046
rect 33686 6984 33692 6996
rect 33647 6956 33692 6984
rect 33686 6944 33692 6956
rect 33744 6944 33750 6996
rect 18046 6808 18052 6860
rect 18104 6848 18110 6860
rect 18233 6851 18291 6857
rect 18233 6848 18245 6851
rect 18104 6820 18245 6848
rect 18104 6808 18110 6820
rect 18233 6817 18245 6820
rect 18279 6817 18291 6851
rect 18233 6811 18291 6817
rect 2682 6780 2688 6792
rect 2643 6752 2688 6780
rect 2682 6740 2688 6752
rect 2740 6740 2746 6792
rect 18325 6783 18383 6789
rect 18325 6749 18337 6783
rect 18371 6780 18383 6783
rect 18414 6780 18420 6792
rect 18371 6752 18420 6780
rect 18371 6749 18383 6752
rect 18325 6743 18383 6749
rect 18414 6740 18420 6752
rect 18472 6740 18478 6792
rect 46290 6740 46296 6792
rect 46348 6780 46354 6792
rect 46753 6783 46811 6789
rect 46753 6780 46765 6783
rect 46348 6752 46765 6780
rect 46348 6740 46354 6752
rect 46753 6749 46765 6752
rect 46799 6749 46811 6783
rect 46753 6743 46811 6749
rect 47673 6783 47731 6789
rect 47673 6749 47685 6783
rect 47719 6780 47731 6783
rect 48130 6780 48136 6792
rect 47719 6752 48136 6780
rect 47719 6749 47731 6752
rect 47673 6743 47731 6749
rect 48130 6740 48136 6752
rect 48188 6740 48194 6792
rect 2314 6604 2320 6656
rect 2372 6644 2378 6656
rect 2593 6647 2651 6653
rect 2593 6644 2605 6647
rect 2372 6616 2605 6644
rect 2372 6604 2378 6616
rect 2593 6613 2605 6616
rect 2639 6613 2651 6647
rect 2593 6607 2651 6613
rect 1104 6554 48852 6576
rect 1104 6502 16880 6554
rect 16932 6502 16944 6554
rect 16996 6502 17008 6554
rect 17060 6502 17072 6554
rect 17124 6502 17136 6554
rect 17188 6502 32811 6554
rect 32863 6502 32875 6554
rect 32927 6502 32939 6554
rect 32991 6502 33003 6554
rect 33055 6502 33067 6554
rect 33119 6502 48852 6554
rect 1104 6480 48852 6502
rect 2314 6372 2320 6384
rect 2275 6344 2320 6372
rect 2314 6332 2320 6344
rect 2372 6332 2378 6384
rect 2130 6304 2136 6316
rect 2091 6276 2136 6304
rect 2130 6264 2136 6276
rect 2188 6264 2194 6316
rect 47486 6264 47492 6316
rect 47544 6304 47550 6316
rect 47581 6307 47639 6313
rect 47581 6304 47593 6307
rect 47544 6276 47593 6304
rect 47544 6264 47550 6276
rect 47581 6273 47593 6276
rect 47627 6273 47639 6307
rect 47581 6267 47639 6273
rect 2774 6236 2780 6248
rect 2735 6208 2780 6236
rect 2774 6196 2780 6208
rect 2832 6196 2838 6248
rect 45186 6236 45192 6248
rect 45147 6208 45192 6236
rect 45186 6196 45192 6208
rect 45244 6196 45250 6248
rect 45370 6236 45376 6248
rect 45331 6208 45376 6236
rect 45370 6196 45376 6208
rect 45428 6196 45434 6248
rect 46566 6236 46572 6248
rect 46527 6208 46572 6236
rect 46566 6196 46572 6208
rect 46624 6196 46630 6248
rect 46382 6060 46388 6112
rect 46440 6100 46446 6112
rect 47673 6103 47731 6109
rect 47673 6100 47685 6103
rect 46440 6072 47685 6100
rect 46440 6060 46446 6072
rect 47673 6069 47685 6072
rect 47719 6069 47731 6103
rect 47673 6063 47731 6069
rect 1104 6010 48852 6032
rect 1104 5958 8915 6010
rect 8967 5958 8979 6010
rect 9031 5958 9043 6010
rect 9095 5958 9107 6010
rect 9159 5958 9171 6010
rect 9223 5958 24846 6010
rect 24898 5958 24910 6010
rect 24962 5958 24974 6010
rect 25026 5958 25038 6010
rect 25090 5958 25102 6010
rect 25154 5958 40776 6010
rect 40828 5958 40840 6010
rect 40892 5958 40904 6010
rect 40956 5958 40968 6010
rect 41020 5958 41032 6010
rect 41084 5958 48852 6010
rect 1104 5936 48852 5958
rect 45186 5896 45192 5908
rect 45147 5868 45192 5896
rect 45186 5856 45192 5868
rect 45244 5856 45250 5908
rect 46658 5760 46664 5772
rect 46619 5732 46664 5760
rect 46658 5720 46664 5732
rect 46716 5720 46722 5772
rect 48130 5760 48136 5772
rect 48091 5732 48136 5760
rect 48130 5720 48136 5732
rect 48188 5720 48194 5772
rect 1946 5692 1952 5704
rect 1907 5664 1952 5692
rect 1946 5652 1952 5664
rect 2004 5652 2010 5704
rect 2498 5652 2504 5704
rect 2556 5692 2562 5704
rect 2593 5695 2651 5701
rect 2593 5692 2605 5695
rect 2556 5664 2605 5692
rect 2556 5652 2562 5664
rect 2593 5661 2605 5664
rect 2639 5661 2651 5695
rect 3234 5692 3240 5704
rect 3195 5664 3240 5692
rect 2593 5655 2651 5661
rect 2608 5624 2636 5655
rect 3234 5652 3240 5664
rect 3292 5652 3298 5704
rect 5718 5692 5724 5704
rect 5679 5664 5724 5692
rect 5718 5652 5724 5664
rect 5776 5652 5782 5704
rect 45646 5692 45652 5704
rect 45607 5664 45652 5692
rect 45646 5652 45652 5664
rect 45704 5652 45710 5704
rect 27982 5624 27988 5636
rect 2608 5596 27988 5624
rect 27982 5584 27988 5596
rect 28040 5584 28046 5636
rect 47946 5624 47952 5636
rect 47907 5596 47952 5624
rect 47946 5584 47952 5596
rect 48004 5584 48010 5636
rect 2314 5516 2320 5568
rect 2372 5556 2378 5568
rect 2501 5559 2559 5565
rect 2501 5556 2513 5559
rect 2372 5528 2513 5556
rect 2372 5516 2378 5528
rect 2501 5525 2513 5528
rect 2547 5525 2559 5559
rect 2501 5519 2559 5525
rect 1104 5466 48852 5488
rect 1104 5414 16880 5466
rect 16932 5414 16944 5466
rect 16996 5414 17008 5466
rect 17060 5414 17072 5466
rect 17124 5414 17136 5466
rect 17188 5414 32811 5466
rect 32863 5414 32875 5466
rect 32927 5414 32939 5466
rect 32991 5414 33003 5466
rect 33055 5414 33067 5466
rect 33119 5414 48852 5466
rect 1104 5392 48852 5414
rect 47673 5355 47731 5361
rect 47673 5321 47685 5355
rect 47719 5352 47731 5355
rect 47946 5352 47952 5364
rect 47719 5324 47952 5352
rect 47719 5321 47731 5324
rect 47673 5315 47731 5321
rect 47946 5312 47952 5324
rect 48004 5312 48010 5364
rect 2314 5284 2320 5296
rect 2275 5256 2320 5284
rect 2314 5244 2320 5256
rect 2372 5244 2378 5296
rect 10226 5284 10232 5296
rect 5644 5256 10232 5284
rect 1946 5176 1952 5228
rect 2004 5216 2010 5228
rect 5644 5225 5672 5256
rect 10226 5244 10232 5256
rect 10284 5244 10290 5296
rect 45646 5284 45652 5296
rect 45204 5256 45652 5284
rect 2133 5219 2191 5225
rect 2133 5216 2145 5219
rect 2004 5188 2145 5216
rect 2004 5176 2010 5188
rect 2133 5185 2145 5188
rect 2179 5185 2191 5219
rect 2133 5179 2191 5185
rect 5629 5219 5687 5225
rect 5629 5185 5641 5219
rect 5675 5185 5687 5219
rect 5629 5179 5687 5185
rect 6917 5219 6975 5225
rect 6917 5185 6929 5219
rect 6963 5216 6975 5219
rect 8294 5216 8300 5228
rect 6963 5188 8300 5216
rect 6963 5185 6975 5188
rect 6917 5179 6975 5185
rect 8294 5176 8300 5188
rect 8352 5176 8358 5228
rect 27982 5216 27988 5228
rect 27895 5188 27988 5216
rect 27982 5176 27988 5188
rect 28040 5216 28046 5228
rect 31478 5216 31484 5228
rect 28040 5188 31484 5216
rect 28040 5176 28046 5188
rect 31478 5176 31484 5188
rect 31536 5176 31542 5228
rect 45204 5225 45232 5256
rect 45646 5244 45652 5256
rect 45704 5244 45710 5296
rect 45189 5219 45247 5225
rect 45189 5185 45201 5219
rect 45235 5185 45247 5219
rect 45189 5179 45247 5185
rect 47302 5176 47308 5228
rect 47360 5216 47366 5228
rect 47581 5219 47639 5225
rect 47581 5216 47593 5219
rect 47360 5188 47593 5216
rect 47360 5176 47366 5188
rect 47581 5185 47593 5188
rect 47627 5185 47639 5219
rect 47581 5179 47639 5185
rect 2774 5148 2780 5160
rect 2735 5120 2780 5148
rect 2774 5108 2780 5120
rect 2832 5108 2838 5160
rect 45373 5151 45431 5157
rect 45373 5117 45385 5151
rect 45419 5148 45431 5151
rect 46382 5148 46388 5160
rect 45419 5120 46388 5148
rect 45419 5117 45431 5120
rect 45373 5111 45431 5117
rect 46382 5108 46388 5120
rect 46440 5108 46446 5160
rect 46842 5148 46848 5160
rect 46803 5120 46848 5148
rect 46842 5108 46848 5120
rect 46900 5108 46906 5160
rect 1486 5012 1492 5024
rect 1447 4984 1492 5012
rect 1486 4972 1492 4984
rect 1544 4972 1550 5024
rect 5166 4972 5172 5024
rect 5224 5012 5230 5024
rect 5537 5015 5595 5021
rect 5537 5012 5549 5015
rect 5224 4984 5549 5012
rect 5224 4972 5230 4984
rect 5537 4981 5549 4984
rect 5583 4981 5595 5015
rect 5537 4975 5595 4981
rect 6546 4972 6552 5024
rect 6604 5012 6610 5024
rect 6825 5015 6883 5021
rect 6825 5012 6837 5015
rect 6604 4984 6837 5012
rect 6604 4972 6610 4984
rect 6825 4981 6837 4984
rect 6871 4981 6883 5015
rect 28074 5012 28080 5024
rect 28035 4984 28080 5012
rect 6825 4975 6883 4981
rect 28074 4972 28080 4984
rect 28132 4972 28138 5024
rect 32674 4972 32680 5024
rect 32732 5012 32738 5024
rect 33045 5015 33103 5021
rect 33045 5012 33057 5015
rect 32732 4984 33057 5012
rect 32732 4972 32738 4984
rect 33045 4981 33057 4984
rect 33091 4981 33103 5015
rect 33045 4975 33103 4981
rect 44085 5015 44143 5021
rect 44085 4981 44097 5015
rect 44131 5012 44143 5015
rect 44450 5012 44456 5024
rect 44131 4984 44456 5012
rect 44131 4981 44143 4984
rect 44085 4975 44143 4981
rect 44450 4972 44456 4984
rect 44508 4972 44514 5024
rect 44726 5012 44732 5024
rect 44687 4984 44732 5012
rect 44726 4972 44732 4984
rect 44784 4972 44790 5024
rect 1104 4922 48852 4944
rect 1104 4870 8915 4922
rect 8967 4870 8979 4922
rect 9031 4870 9043 4922
rect 9095 4870 9107 4922
rect 9159 4870 9171 4922
rect 9223 4870 24846 4922
rect 24898 4870 24910 4922
rect 24962 4870 24974 4922
rect 25026 4870 25038 4922
rect 25090 4870 25102 4922
rect 25154 4870 40776 4922
rect 40828 4870 40840 4922
rect 40892 4870 40904 4922
rect 40956 4870 40968 4922
rect 41020 4870 41032 4922
rect 41084 4870 48852 4922
rect 1104 4848 48852 4870
rect 45281 4811 45339 4817
rect 45281 4777 45293 4811
rect 45327 4808 45339 4811
rect 45370 4808 45376 4820
rect 45327 4780 45376 4808
rect 45327 4777 45339 4780
rect 45281 4771 45339 4777
rect 45370 4768 45376 4780
rect 45428 4768 45434 4820
rect 1394 4672 1400 4684
rect 1355 4644 1400 4672
rect 1394 4632 1400 4644
rect 1452 4632 1458 4684
rect 3234 4672 3240 4684
rect 3195 4644 3240 4672
rect 3234 4632 3240 4644
rect 3292 4632 3298 4684
rect 5166 4672 5172 4684
rect 5127 4644 5172 4672
rect 5166 4632 5172 4644
rect 5224 4632 5230 4684
rect 5534 4672 5540 4684
rect 5495 4644 5540 4672
rect 5534 4632 5540 4644
rect 5592 4632 5598 4684
rect 46290 4672 46296 4684
rect 42352 4644 45232 4672
rect 46251 4644 46296 4672
rect 42352 4616 42380 4644
rect 3973 4607 4031 4613
rect 3973 4573 3985 4607
rect 4019 4604 4031 4607
rect 4062 4604 4068 4616
rect 4019 4576 4068 4604
rect 4019 4573 4031 4576
rect 3973 4567 4031 4573
rect 4062 4564 4068 4576
rect 4120 4564 4126 4616
rect 4982 4604 4988 4616
rect 4943 4576 4988 4604
rect 4982 4564 4988 4576
rect 5040 4564 5046 4616
rect 8754 4564 8760 4616
rect 8812 4604 8818 4616
rect 8941 4607 8999 4613
rect 8941 4604 8953 4607
rect 8812 4576 8953 4604
rect 8812 4564 8818 4576
rect 8941 4573 8953 4576
rect 8987 4573 8999 4607
rect 15746 4604 15752 4616
rect 15707 4576 15752 4604
rect 8941 4567 8999 4573
rect 15746 4564 15752 4576
rect 15804 4564 15810 4616
rect 27890 4604 27896 4616
rect 27851 4576 27896 4604
rect 27890 4564 27896 4576
rect 27948 4564 27954 4616
rect 28721 4607 28779 4613
rect 28721 4573 28733 4607
rect 28767 4604 28779 4607
rect 28994 4604 29000 4616
rect 28767 4576 29000 4604
rect 28767 4573 28779 4576
rect 28721 4567 28779 4573
rect 28994 4564 29000 4576
rect 29052 4564 29058 4616
rect 32030 4604 32036 4616
rect 31991 4576 32036 4604
rect 32030 4564 32036 4576
rect 32088 4564 32094 4616
rect 32766 4564 32772 4616
rect 32824 4604 32830 4616
rect 33045 4607 33103 4613
rect 33045 4604 33057 4607
rect 32824 4576 33057 4604
rect 32824 4564 32830 4576
rect 33045 4573 33057 4576
rect 33091 4573 33103 4607
rect 33045 4567 33103 4573
rect 34149 4607 34207 4613
rect 34149 4573 34161 4607
rect 34195 4604 34207 4607
rect 34514 4604 34520 4616
rect 34195 4576 34520 4604
rect 34195 4573 34207 4576
rect 34149 4567 34207 4573
rect 34514 4564 34520 4576
rect 34572 4564 34578 4616
rect 34698 4604 34704 4616
rect 34659 4576 34704 4604
rect 34698 4564 34704 4576
rect 34756 4564 34762 4616
rect 35894 4564 35900 4616
rect 35952 4604 35958 4616
rect 37185 4607 37243 4613
rect 35952 4576 35997 4604
rect 35952 4564 35958 4576
rect 37185 4573 37197 4607
rect 37231 4604 37243 4607
rect 37274 4604 37280 4616
rect 37231 4576 37280 4604
rect 37231 4573 37243 4576
rect 37185 4567 37243 4573
rect 37274 4564 37280 4576
rect 37332 4564 37338 4616
rect 42334 4604 42340 4616
rect 42295 4576 42340 4604
rect 42334 4564 42340 4576
rect 42392 4564 42398 4616
rect 43254 4604 43260 4616
rect 43215 4576 43260 4604
rect 43254 4564 43260 4576
rect 43312 4564 43318 4616
rect 43714 4604 43720 4616
rect 43675 4576 43720 4604
rect 43714 4564 43720 4576
rect 43772 4564 43778 4616
rect 45204 4613 45232 4644
rect 46290 4632 46296 4644
rect 46348 4632 46354 4684
rect 45189 4607 45247 4613
rect 45189 4573 45201 4607
rect 45235 4604 45247 4607
rect 45462 4604 45468 4616
rect 45235 4576 45468 4604
rect 45235 4573 45247 4576
rect 45189 4567 45247 4573
rect 45462 4564 45468 4576
rect 45520 4564 45526 4616
rect 3053 4539 3111 4545
rect 3053 4505 3065 4539
rect 3099 4536 3111 4539
rect 3881 4539 3939 4545
rect 3881 4536 3893 4539
rect 3099 4508 3893 4536
rect 3099 4505 3111 4508
rect 3053 4499 3111 4505
rect 3881 4505 3893 4508
rect 3927 4505 3939 4539
rect 7834 4536 7840 4548
rect 7795 4508 7840 4536
rect 3881 4499 3939 4505
rect 7834 4496 7840 4508
rect 7892 4496 7898 4548
rect 8205 4539 8263 4545
rect 8205 4505 8217 4539
rect 8251 4536 8263 4539
rect 9950 4536 9956 4548
rect 8251 4508 9956 4536
rect 8251 4505 8263 4508
rect 8205 4499 8263 4505
rect 2682 4428 2688 4480
rect 2740 4468 2746 4480
rect 8220 4468 8248 4499
rect 9950 4496 9956 4508
rect 10008 4536 10014 4548
rect 10410 4536 10416 4548
rect 10008 4508 10416 4536
rect 10008 4496 10014 4508
rect 10410 4496 10416 4508
rect 10468 4496 10474 4548
rect 46477 4539 46535 4545
rect 46477 4505 46489 4539
rect 46523 4536 46535 4539
rect 46658 4536 46664 4548
rect 46523 4508 46664 4536
rect 46523 4505 46535 4508
rect 46477 4499 46535 4505
rect 46658 4496 46664 4508
rect 46716 4496 46722 4548
rect 48133 4539 48191 4545
rect 48133 4505 48145 4539
rect 48179 4536 48191 4539
rect 48314 4536 48320 4548
rect 48179 4508 48320 4536
rect 48179 4505 48191 4508
rect 48133 4499 48191 4505
rect 48314 4496 48320 4508
rect 48372 4496 48378 4548
rect 33134 4468 33140 4480
rect 2740 4440 8248 4468
rect 33095 4440 33140 4468
rect 2740 4428 2746 4440
rect 33134 4428 33140 4440
rect 33192 4428 33198 4480
rect 34790 4468 34796 4480
rect 34751 4440 34796 4468
rect 34790 4428 34796 4440
rect 34848 4428 34854 4480
rect 42429 4471 42487 4477
rect 42429 4437 42441 4471
rect 42475 4468 42487 4471
rect 42610 4468 42616 4480
rect 42475 4440 42616 4468
rect 42475 4437 42487 4440
rect 42429 4431 42487 4437
rect 42610 4428 42616 4440
rect 42668 4428 42674 4480
rect 43162 4468 43168 4480
rect 43123 4440 43168 4468
rect 43162 4428 43168 4440
rect 43220 4428 43226 4480
rect 1104 4378 48852 4400
rect 1104 4326 16880 4378
rect 16932 4326 16944 4378
rect 16996 4326 17008 4378
rect 17060 4326 17072 4378
rect 17124 4326 17136 4378
rect 17188 4326 32811 4378
rect 32863 4326 32875 4378
rect 32927 4326 32939 4378
rect 32991 4326 33003 4378
rect 33055 4326 33067 4378
rect 33119 4326 48852 4378
rect 1104 4304 48852 4326
rect 4062 4196 4068 4208
rect 3160 4168 4068 4196
rect 2225 4131 2283 4137
rect 2225 4097 2237 4131
rect 2271 4128 2283 4131
rect 3160 4128 3188 4168
rect 4062 4156 4068 4168
rect 4120 4156 4126 4208
rect 6546 4196 6552 4208
rect 6507 4168 6552 4196
rect 6546 4156 6552 4168
rect 6604 4156 6610 4208
rect 28074 4196 28080 4208
rect 28035 4168 28080 4196
rect 28074 4156 28080 4168
rect 28132 4156 28138 4208
rect 33134 4196 33140 4208
rect 33095 4168 33140 4196
rect 33134 4156 33140 4168
rect 33192 4156 33198 4208
rect 4982 4128 4988 4140
rect 2271 4100 3188 4128
rect 4943 4100 4988 4128
rect 2271 4097 2283 4100
rect 2225 4091 2283 4097
rect 4982 4088 4988 4100
rect 5040 4088 5046 4140
rect 8294 4088 8300 4140
rect 8352 4128 8358 4140
rect 9217 4131 9275 4137
rect 9217 4128 9229 4131
rect 8352 4100 9229 4128
rect 8352 4088 8358 4100
rect 9217 4097 9229 4100
rect 9263 4097 9275 4131
rect 9217 4091 9275 4097
rect 2866 4060 2872 4072
rect 2827 4032 2872 4060
rect 2866 4020 2872 4032
rect 2924 4020 2930 4072
rect 3878 4020 3884 4072
rect 3936 4060 3942 4072
rect 4341 4063 4399 4069
rect 4341 4060 4353 4063
rect 3936 4032 4353 4060
rect 3936 4020 3942 4032
rect 4341 4029 4353 4032
rect 4387 4029 4399 4063
rect 4522 4060 4528 4072
rect 4483 4032 4528 4060
rect 4341 4023 4399 4029
rect 4522 4020 4528 4032
rect 4580 4020 4586 4072
rect 5258 4020 5264 4072
rect 5316 4060 5322 4072
rect 6365 4063 6423 4069
rect 6365 4060 6377 4063
rect 5316 4032 6377 4060
rect 5316 4020 5322 4032
rect 6365 4029 6377 4032
rect 6411 4029 6423 4063
rect 6365 4023 6423 4029
rect 6825 4063 6883 4069
rect 6825 4029 6837 4063
rect 6871 4029 6883 4063
rect 9232 4060 9260 4091
rect 15102 4088 15108 4140
rect 15160 4128 15166 4140
rect 15841 4131 15899 4137
rect 15841 4128 15853 4131
rect 15160 4100 15853 4128
rect 15160 4088 15166 4100
rect 15841 4097 15853 4100
rect 15887 4128 15899 4131
rect 17954 4128 17960 4140
rect 15887 4100 17960 4128
rect 15887 4097 15899 4100
rect 15841 4091 15899 4097
rect 17954 4088 17960 4100
rect 18012 4088 18018 4140
rect 20162 4088 20168 4140
rect 20220 4128 20226 4140
rect 26973 4131 27031 4137
rect 26973 4128 26985 4131
rect 20220 4100 26985 4128
rect 20220 4088 20226 4100
rect 26973 4097 26985 4100
rect 27019 4128 27031 4131
rect 27706 4128 27712 4140
rect 27019 4100 27712 4128
rect 27019 4097 27031 4100
rect 26973 4091 27031 4097
rect 27706 4088 27712 4100
rect 27764 4088 27770 4140
rect 27890 4128 27896 4140
rect 27851 4100 27896 4128
rect 27890 4088 27896 4100
rect 27948 4088 27954 4140
rect 32122 4128 32128 4140
rect 32083 4100 32128 4128
rect 32122 4088 32128 4100
rect 32180 4088 32186 4140
rect 32674 4088 32680 4140
rect 32732 4128 32738 4140
rect 32953 4131 33011 4137
rect 32953 4128 32965 4131
rect 32732 4100 32965 4128
rect 32732 4088 32738 4100
rect 32953 4097 32965 4100
rect 32999 4097 33011 4131
rect 32953 4091 33011 4097
rect 35897 4131 35955 4137
rect 35897 4097 35909 4131
rect 35943 4097 35955 4131
rect 36538 4128 36544 4140
rect 36499 4100 36544 4128
rect 35897 4091 35955 4097
rect 18690 4060 18696 4072
rect 9232 4032 16574 4060
rect 18651 4032 18696 4060
rect 6825 4023 6883 4029
rect 3970 3952 3976 4004
rect 4028 3992 4034 4004
rect 6840 3992 6868 4023
rect 4028 3964 6868 3992
rect 4028 3952 4034 3964
rect 7466 3952 7472 4004
rect 7524 3992 7530 4004
rect 7834 3992 7840 4004
rect 7524 3964 7840 3992
rect 7524 3952 7530 3964
rect 7834 3952 7840 3964
rect 7892 3992 7898 4004
rect 13170 3992 13176 4004
rect 7892 3964 13176 3992
rect 7892 3952 7898 3964
rect 13170 3952 13176 3964
rect 13228 3952 13234 4004
rect 13817 3995 13875 4001
rect 13817 3961 13829 3995
rect 13863 3992 13875 3995
rect 15470 3992 15476 4004
rect 13863 3964 15476 3992
rect 13863 3961 13875 3964
rect 13817 3955 13875 3961
rect 15470 3952 15476 3964
rect 15528 3952 15534 4004
rect 16546 3992 16574 4032
rect 18690 4020 18696 4032
rect 18748 4020 18754 4072
rect 19334 4020 19340 4072
rect 19392 4060 19398 4072
rect 19889 4063 19947 4069
rect 19889 4060 19901 4063
rect 19392 4032 19901 4060
rect 19392 4020 19398 4032
rect 19889 4029 19901 4032
rect 19935 4029 19947 4063
rect 20070 4060 20076 4072
rect 20031 4032 20076 4060
rect 19889 4023 19947 4029
rect 20070 4020 20076 4032
rect 20128 4020 20134 4072
rect 25498 4020 25504 4072
rect 25556 4060 25562 4072
rect 27246 4060 27252 4072
rect 25556 4032 27252 4060
rect 25556 4020 25562 4032
rect 27246 4020 27252 4032
rect 27304 4020 27310 4072
rect 28350 4060 28356 4072
rect 28311 4032 28356 4060
rect 28350 4020 28356 4032
rect 28408 4020 28414 4072
rect 33502 4060 33508 4072
rect 33463 4032 33508 4060
rect 33502 4020 33508 4032
rect 33560 4020 33566 4072
rect 35912 4060 35940 4091
rect 36538 4088 36544 4100
rect 36596 4088 36602 4140
rect 37274 4128 37280 4140
rect 37235 4100 37280 4128
rect 37274 4088 37280 4100
rect 37332 4088 37338 4140
rect 40126 4128 40132 4140
rect 39684 4100 40132 4128
rect 36633 4063 36691 4069
rect 35912 4032 36584 4060
rect 27430 3992 27436 4004
rect 16546 3964 27436 3992
rect 27430 3952 27436 3964
rect 27488 3952 27494 4004
rect 32122 3952 32128 4004
rect 32180 3992 32186 4004
rect 36556 3992 36584 4032
rect 36633 4029 36645 4063
rect 36679 4060 36691 4063
rect 37461 4063 37519 4069
rect 37461 4060 37473 4063
rect 36679 4032 37473 4060
rect 36679 4029 36691 4032
rect 36633 4023 36691 4029
rect 37461 4029 37473 4032
rect 37507 4029 37519 4063
rect 37461 4023 37519 4029
rect 37550 4020 37556 4072
rect 37608 4060 37614 4072
rect 37737 4063 37795 4069
rect 37737 4060 37749 4063
rect 37608 4032 37749 4060
rect 37608 4020 37614 4032
rect 37737 4029 37749 4032
rect 37783 4029 37795 4063
rect 37737 4023 37795 4029
rect 39684 3992 39712 4100
rect 40126 4088 40132 4100
rect 40184 4088 40190 4140
rect 44726 4128 44732 4140
rect 44687 4100 44732 4128
rect 44726 4088 44732 4100
rect 44784 4088 44790 4140
rect 47578 4128 47584 4140
rect 47539 4100 47584 4128
rect 47578 4088 47584 4100
rect 47636 4088 47642 4140
rect 32180 3964 36492 3992
rect 36556 3964 39712 3992
rect 39776 4032 41828 4060
rect 32180 3952 32186 3964
rect 1578 3884 1584 3936
rect 1636 3924 1642 3936
rect 2133 3927 2191 3933
rect 2133 3924 2145 3927
rect 1636 3896 2145 3924
rect 1636 3884 1642 3896
rect 2133 3893 2145 3896
rect 2179 3893 2191 3927
rect 5810 3924 5816 3936
rect 5771 3896 5816 3924
rect 2133 3887 2191 3893
rect 5810 3884 5816 3896
rect 5868 3884 5874 3936
rect 9306 3924 9312 3936
rect 9267 3896 9312 3924
rect 9306 3884 9312 3896
rect 9364 3884 9370 3936
rect 9858 3924 9864 3936
rect 9819 3896 9864 3924
rect 9858 3884 9864 3896
rect 9916 3884 9922 3936
rect 11606 3884 11612 3936
rect 11664 3924 11670 3936
rect 11701 3927 11759 3933
rect 11701 3924 11713 3927
rect 11664 3896 11713 3924
rect 11664 3884 11670 3896
rect 11701 3893 11713 3896
rect 11747 3893 11759 3927
rect 12526 3924 12532 3936
rect 12487 3896 12532 3924
rect 11701 3887 11759 3893
rect 12526 3884 12532 3896
rect 12584 3884 12590 3936
rect 14182 3884 14188 3936
rect 14240 3924 14246 3936
rect 14277 3927 14335 3933
rect 14277 3924 14289 3927
rect 14240 3896 14289 3924
rect 14240 3884 14246 3896
rect 14277 3893 14289 3896
rect 14323 3893 14335 3927
rect 15930 3924 15936 3936
rect 15891 3896 15936 3924
rect 14277 3887 14335 3893
rect 15930 3884 15936 3896
rect 15988 3884 15994 3936
rect 18138 3884 18144 3936
rect 18196 3924 18202 3936
rect 25774 3924 25780 3936
rect 18196 3896 25780 3924
rect 18196 3884 18202 3896
rect 25774 3884 25780 3896
rect 25832 3884 25838 3936
rect 31570 3924 31576 3936
rect 31531 3896 31576 3924
rect 31570 3884 31576 3896
rect 31628 3884 31634 3936
rect 32214 3924 32220 3936
rect 32175 3896 32220 3924
rect 32214 3884 32220 3896
rect 32272 3884 32278 3936
rect 34882 3884 34888 3936
rect 34940 3924 34946 3936
rect 35253 3927 35311 3933
rect 35253 3924 35265 3927
rect 34940 3896 35265 3924
rect 34940 3884 34946 3896
rect 35253 3893 35265 3896
rect 35299 3893 35311 3927
rect 35253 3887 35311 3893
rect 35989 3927 36047 3933
rect 35989 3893 36001 3927
rect 36035 3924 36047 3927
rect 36078 3924 36084 3936
rect 36035 3896 36084 3924
rect 36035 3893 36047 3896
rect 35989 3887 36047 3893
rect 36078 3884 36084 3896
rect 36136 3884 36142 3936
rect 36464 3924 36492 3964
rect 39776 3924 39804 4032
rect 41800 3992 41828 4032
rect 41874 4020 41880 4072
rect 41932 4060 41938 4072
rect 42429 4063 42487 4069
rect 42429 4060 42441 4063
rect 41932 4032 42441 4060
rect 41932 4020 41938 4032
rect 42429 4029 42441 4032
rect 42475 4029 42487 4063
rect 42429 4023 42487 4029
rect 42613 4063 42671 4069
rect 42613 4029 42625 4063
rect 42659 4060 42671 4063
rect 43162 4060 43168 4072
rect 42659 4032 43168 4060
rect 42659 4029 42671 4032
rect 42613 4023 42671 4029
rect 43162 4020 43168 4032
rect 43220 4020 43226 4072
rect 44269 4063 44327 4069
rect 44269 4029 44281 4063
rect 44315 4029 44327 4063
rect 44269 4023 44327 4029
rect 44913 4063 44971 4069
rect 44913 4029 44925 4063
rect 44959 4060 44971 4063
rect 45094 4060 45100 4072
rect 44959 4032 45100 4060
rect 44959 4029 44971 4032
rect 44913 4023 44971 4029
rect 43254 3992 43260 4004
rect 41800 3964 43260 3992
rect 43254 3952 43260 3964
rect 43312 3952 43318 4004
rect 44284 3992 44312 4023
rect 45094 4020 45100 4032
rect 45152 4020 45158 4072
rect 46569 4063 46627 4069
rect 46569 4029 46581 4063
rect 46615 4060 46627 4063
rect 47026 4060 47032 4072
rect 46615 4032 47032 4060
rect 46615 4029 46627 4032
rect 46569 4023 46627 4029
rect 47026 4020 47032 4032
rect 47084 4020 47090 4072
rect 46842 3992 46848 4004
rect 44284 3964 46848 3992
rect 46842 3952 46848 3964
rect 46900 3952 46906 4004
rect 39942 3924 39948 3936
rect 36464 3896 39804 3924
rect 39903 3896 39948 3924
rect 39942 3884 39948 3896
rect 40000 3884 40006 3936
rect 41877 3927 41935 3933
rect 41877 3893 41889 3927
rect 41923 3924 41935 3927
rect 42426 3924 42432 3936
rect 41923 3896 42432 3924
rect 41923 3893 41935 3896
rect 41877 3887 41935 3893
rect 42426 3884 42432 3896
rect 42484 3884 42490 3936
rect 46474 3884 46480 3936
rect 46532 3924 46538 3936
rect 47673 3927 47731 3933
rect 47673 3924 47685 3927
rect 46532 3896 47685 3924
rect 46532 3884 46538 3896
rect 47673 3893 47685 3896
rect 47719 3893 47731 3927
rect 47673 3887 47731 3893
rect 1104 3834 48852 3856
rect 1104 3782 8915 3834
rect 8967 3782 8979 3834
rect 9031 3782 9043 3834
rect 9095 3782 9107 3834
rect 9159 3782 9171 3834
rect 9223 3782 24846 3834
rect 24898 3782 24910 3834
rect 24962 3782 24974 3834
rect 25026 3782 25038 3834
rect 25090 3782 25102 3834
rect 25154 3782 40776 3834
rect 40828 3782 40840 3834
rect 40892 3782 40904 3834
rect 40956 3782 40968 3834
rect 41020 3782 41032 3834
rect 41084 3782 48852 3834
rect 1104 3760 48852 3782
rect 3878 3720 3884 3732
rect 3839 3692 3884 3720
rect 3878 3680 3884 3692
rect 3936 3680 3942 3732
rect 4433 3723 4491 3729
rect 4433 3689 4445 3723
rect 4479 3720 4491 3723
rect 4522 3720 4528 3732
rect 4479 3692 4528 3720
rect 4479 3689 4491 3692
rect 4433 3683 4491 3689
rect 4522 3680 4528 3692
rect 4580 3680 4586 3732
rect 5258 3720 5264 3732
rect 5219 3692 5264 3720
rect 5258 3680 5264 3692
rect 5316 3680 5322 3732
rect 11698 3720 11704 3732
rect 6886 3692 11704 3720
rect 1486 3652 1492 3664
rect 1412 3624 1492 3652
rect 1412 3593 1440 3624
rect 1486 3612 1492 3624
rect 1544 3612 1550 3664
rect 4062 3612 4068 3664
rect 4120 3652 4126 3664
rect 6886 3652 6914 3692
rect 11698 3680 11704 3692
rect 11756 3720 11762 3732
rect 19334 3720 19340 3732
rect 11756 3692 18000 3720
rect 19295 3692 19340 3720
rect 11756 3680 11762 3692
rect 9858 3652 9864 3664
rect 4120 3624 6914 3652
rect 9140 3624 9864 3652
rect 4120 3612 4126 3624
rect 1397 3587 1455 3593
rect 1397 3553 1409 3587
rect 1443 3553 1455 3587
rect 1578 3584 1584 3596
rect 1539 3556 1584 3584
rect 1397 3547 1455 3553
rect 1578 3544 1584 3556
rect 1636 3544 1642 3596
rect 2774 3584 2780 3596
rect 2735 3556 2780 3584
rect 2774 3544 2780 3556
rect 2832 3544 2838 3596
rect 5718 3584 5724 3596
rect 5679 3556 5724 3584
rect 5718 3544 5724 3556
rect 5776 3544 5782 3596
rect 5902 3544 5908 3596
rect 5960 3584 5966 3596
rect 9140 3593 9168 3624
rect 9858 3612 9864 3624
rect 9916 3612 9922 3664
rect 9950 3612 9956 3664
rect 10008 3652 10014 3664
rect 10008 3624 13032 3652
rect 10008 3612 10014 3624
rect 6181 3587 6239 3593
rect 6181 3584 6193 3587
rect 5960 3556 6193 3584
rect 5960 3544 5966 3556
rect 6181 3553 6193 3556
rect 6227 3553 6239 3587
rect 6181 3547 6239 3553
rect 9125 3587 9183 3593
rect 9125 3553 9137 3587
rect 9171 3553 9183 3587
rect 9306 3584 9312 3596
rect 9267 3556 9312 3584
rect 9125 3547 9183 3553
rect 9306 3544 9312 3556
rect 9364 3544 9370 3596
rect 9674 3584 9680 3596
rect 9635 3556 9680 3584
rect 9674 3544 9680 3556
rect 9732 3544 9738 3596
rect 11606 3584 11612 3596
rect 11567 3556 11612 3584
rect 11606 3544 11612 3556
rect 11664 3544 11670 3596
rect 12250 3584 12256 3596
rect 12211 3556 12256 3584
rect 12250 3544 12256 3556
rect 12308 3544 12314 3596
rect 3973 3519 4031 3525
rect 3973 3485 3985 3519
rect 4019 3485 4031 3519
rect 8202 3516 8208 3528
rect 8163 3488 8208 3516
rect 3973 3479 4031 3485
rect 3988 3380 4016 3479
rect 8202 3476 8208 3488
rect 8260 3476 8266 3528
rect 13004 3516 13032 3624
rect 13170 3612 13176 3664
rect 13228 3652 13234 3664
rect 17972 3652 18000 3692
rect 19334 3680 19340 3692
rect 19392 3680 19398 3732
rect 20070 3720 20076 3732
rect 20031 3692 20076 3720
rect 20070 3680 20076 3692
rect 20128 3680 20134 3732
rect 32122 3720 32128 3732
rect 26206 3692 32128 3720
rect 19426 3652 19432 3664
rect 13228 3624 16574 3652
rect 17972 3624 19432 3652
rect 13228 3612 13234 3624
rect 15746 3584 15752 3596
rect 15707 3556 15752 3584
rect 15746 3544 15752 3556
rect 15804 3544 15810 3596
rect 15930 3584 15936 3596
rect 15891 3556 15936 3584
rect 15930 3544 15936 3556
rect 15988 3544 15994 3596
rect 16114 3544 16120 3596
rect 16172 3584 16178 3596
rect 16209 3587 16267 3593
rect 16209 3584 16221 3587
rect 16172 3556 16221 3584
rect 16172 3544 16178 3556
rect 16209 3553 16221 3556
rect 16255 3553 16267 3587
rect 16546 3584 16574 3624
rect 19426 3612 19432 3624
rect 19484 3612 19490 3664
rect 19702 3612 19708 3664
rect 19760 3652 19766 3664
rect 26206 3652 26234 3692
rect 32122 3680 32128 3692
rect 32180 3680 32186 3732
rect 45094 3720 45100 3732
rect 45055 3692 45100 3720
rect 45094 3680 45100 3692
rect 45152 3680 45158 3732
rect 19760 3624 26234 3652
rect 19760 3612 19766 3624
rect 26970 3612 26976 3664
rect 27028 3612 27034 3664
rect 47578 3652 47584 3664
rect 45526 3624 47584 3652
rect 26988 3584 27016 3612
rect 27706 3584 27712 3596
rect 16546 3556 19288 3584
rect 16209 3547 16267 3553
rect 14277 3519 14335 3525
rect 14277 3516 14289 3519
rect 13004 3488 14289 3516
rect 14277 3485 14289 3488
rect 14323 3485 14335 3519
rect 15102 3516 15108 3528
rect 15063 3488 15108 3516
rect 14277 3479 14335 3485
rect 5718 3408 5724 3460
rect 5776 3448 5782 3460
rect 5905 3451 5963 3457
rect 5905 3448 5917 3451
rect 5776 3420 5917 3448
rect 5776 3408 5782 3420
rect 5905 3417 5917 3420
rect 5951 3417 5963 3451
rect 11790 3448 11796 3460
rect 11751 3420 11796 3448
rect 5905 3411 5963 3417
rect 11790 3408 11796 3420
rect 11848 3408 11854 3460
rect 14292 3448 14320 3479
rect 15102 3476 15108 3488
rect 15160 3476 15166 3528
rect 18141 3519 18199 3525
rect 18141 3485 18153 3519
rect 18187 3516 18199 3519
rect 19150 3516 19156 3528
rect 18187 3488 19156 3516
rect 18187 3485 18199 3488
rect 18141 3479 18199 3485
rect 19150 3476 19156 3488
rect 19208 3476 19214 3528
rect 19260 3525 19288 3556
rect 24872 3556 27016 3584
rect 27667 3556 27712 3584
rect 19245 3519 19303 3525
rect 19245 3485 19257 3519
rect 19291 3516 19303 3519
rect 20162 3516 20168 3528
rect 19291 3488 20168 3516
rect 19291 3485 19303 3488
rect 19245 3479 19303 3485
rect 20162 3476 20168 3488
rect 20220 3476 20226 3528
rect 23845 3519 23903 3525
rect 23845 3485 23857 3519
rect 23891 3516 23903 3519
rect 23934 3516 23940 3528
rect 23891 3488 23940 3516
rect 23891 3485 23903 3488
rect 23845 3479 23903 3485
rect 23934 3476 23940 3488
rect 23992 3476 23998 3528
rect 24872 3525 24900 3556
rect 27706 3544 27712 3556
rect 27764 3544 27770 3596
rect 32030 3584 32036 3596
rect 31991 3556 32036 3584
rect 32030 3544 32036 3556
rect 32088 3544 32094 3596
rect 32214 3584 32220 3596
rect 32175 3556 32220 3584
rect 32214 3544 32220 3556
rect 32272 3544 32278 3596
rect 32674 3584 32680 3596
rect 32635 3556 32680 3584
rect 32674 3544 32680 3556
rect 32732 3544 32738 3596
rect 35894 3544 35900 3596
rect 35952 3584 35958 3596
rect 36078 3584 36084 3596
rect 35952 3556 35997 3584
rect 36039 3556 36084 3584
rect 35952 3544 35958 3556
rect 36078 3544 36084 3556
rect 36136 3544 36142 3596
rect 36722 3584 36728 3596
rect 36683 3556 36728 3584
rect 36722 3544 36728 3556
rect 36780 3544 36786 3596
rect 41969 3587 42027 3593
rect 41969 3553 41981 3587
rect 42015 3584 42027 3587
rect 43806 3584 43812 3596
rect 42015 3556 43812 3584
rect 42015 3553 42027 3556
rect 41969 3547 42027 3553
rect 43806 3544 43812 3556
rect 43864 3544 43870 3596
rect 24857 3519 24915 3525
rect 24857 3485 24869 3519
rect 24903 3485 24915 3519
rect 25498 3516 25504 3528
rect 25459 3488 25504 3516
rect 24857 3479 24915 3485
rect 25498 3476 25504 3488
rect 25556 3476 25562 3528
rect 26421 3519 26479 3525
rect 26421 3485 26433 3519
rect 26467 3516 26479 3519
rect 26881 3519 26939 3525
rect 26881 3516 26893 3519
rect 26467 3488 26893 3516
rect 26467 3485 26479 3488
rect 26421 3479 26479 3485
rect 26881 3485 26893 3488
rect 26927 3485 26939 3519
rect 26881 3479 26939 3485
rect 28810 3476 28816 3528
rect 28868 3516 28874 3528
rect 29549 3519 29607 3525
rect 29549 3516 29561 3519
rect 28868 3488 29561 3516
rect 28868 3476 28874 3488
rect 29549 3485 29561 3488
rect 29595 3485 29607 3519
rect 29549 3479 29607 3485
rect 31297 3519 31355 3525
rect 31297 3485 31309 3519
rect 31343 3516 31355 3519
rect 31938 3516 31944 3528
rect 31343 3488 31944 3516
rect 31343 3485 31355 3488
rect 31297 3479 31355 3485
rect 31938 3476 31944 3488
rect 31996 3476 32002 3528
rect 34698 3516 34704 3528
rect 34659 3488 34704 3516
rect 34698 3476 34704 3488
rect 34756 3476 34762 3528
rect 37274 3476 37280 3528
rect 37332 3516 37338 3528
rect 38197 3519 38255 3525
rect 38197 3516 38209 3519
rect 37332 3488 38209 3516
rect 37332 3476 37338 3488
rect 38197 3485 38209 3488
rect 38243 3485 38255 3519
rect 39114 3516 39120 3528
rect 39075 3488 39120 3516
rect 38197 3479 38255 3485
rect 39114 3476 39120 3488
rect 39172 3476 39178 3528
rect 39850 3516 39856 3528
rect 39811 3488 39856 3516
rect 39850 3476 39856 3488
rect 39908 3476 39914 3528
rect 42426 3516 42432 3528
rect 42387 3488 42432 3516
rect 42426 3476 42432 3488
rect 42484 3476 42490 3528
rect 45189 3519 45247 3525
rect 45189 3485 45201 3519
rect 45235 3516 45247 3519
rect 45526 3516 45554 3624
rect 47578 3612 47584 3624
rect 47636 3612 47642 3664
rect 46474 3584 46480 3596
rect 46435 3556 46480 3584
rect 46474 3544 46480 3556
rect 46532 3544 46538 3596
rect 45235 3488 45554 3516
rect 45833 3519 45891 3525
rect 45235 3485 45247 3488
rect 45189 3479 45247 3485
rect 45833 3485 45845 3519
rect 45879 3516 45891 3519
rect 46293 3519 46351 3525
rect 46293 3516 46305 3519
rect 45879 3488 46305 3516
rect 45879 3485 45891 3488
rect 45833 3479 45891 3485
rect 46293 3485 46305 3488
rect 46339 3485 46351 3519
rect 46293 3479 46351 3485
rect 20438 3448 20444 3460
rect 14292 3420 20444 3448
rect 20438 3408 20444 3420
rect 20496 3408 20502 3460
rect 27062 3448 27068 3460
rect 27023 3420 27068 3448
rect 27062 3408 27068 3420
rect 27120 3408 27126 3460
rect 27246 3408 27252 3460
rect 27304 3448 27310 3460
rect 35158 3448 35164 3460
rect 27304 3420 35164 3448
rect 27304 3408 27310 3420
rect 35158 3408 35164 3420
rect 35216 3408 35222 3460
rect 41690 3408 41696 3460
rect 41748 3457 41754 3460
rect 41748 3448 41760 3457
rect 42610 3448 42616 3460
rect 41748 3420 41793 3448
rect 42571 3420 42616 3448
rect 41748 3411 41760 3420
rect 41748 3408 41754 3411
rect 42610 3408 42616 3420
rect 42668 3408 42674 3460
rect 44269 3451 44327 3457
rect 44269 3417 44281 3451
rect 44315 3448 44327 3451
rect 45094 3448 45100 3460
rect 44315 3420 45100 3448
rect 44315 3417 44327 3420
rect 44269 3411 44327 3417
rect 45094 3408 45100 3420
rect 45152 3408 45158 3460
rect 48130 3448 48136 3460
rect 48091 3420 48136 3448
rect 48130 3408 48136 3420
rect 48188 3408 48194 3460
rect 8110 3380 8116 3392
rect 3988 3352 8116 3380
rect 8110 3340 8116 3352
rect 8168 3340 8174 3392
rect 8294 3380 8300 3392
rect 8255 3352 8300 3380
rect 8294 3340 8300 3352
rect 8352 3340 8358 3392
rect 14366 3380 14372 3392
rect 14327 3352 14372 3380
rect 14366 3340 14372 3352
rect 14424 3340 14430 3392
rect 15013 3383 15071 3389
rect 15013 3349 15025 3383
rect 15059 3380 15071 3383
rect 15286 3380 15292 3392
rect 15059 3352 15292 3380
rect 15059 3349 15071 3352
rect 15013 3343 15071 3349
rect 15286 3340 15292 3352
rect 15344 3340 15350 3392
rect 18233 3383 18291 3389
rect 18233 3349 18245 3383
rect 18279 3380 18291 3383
rect 18322 3380 18328 3392
rect 18279 3352 18328 3380
rect 18279 3349 18291 3352
rect 18233 3343 18291 3349
rect 18322 3340 18328 3352
rect 18380 3340 18386 3392
rect 24118 3340 24124 3392
rect 24176 3380 24182 3392
rect 24765 3383 24823 3389
rect 24765 3380 24777 3383
rect 24176 3352 24777 3380
rect 24176 3340 24182 3352
rect 24765 3349 24777 3352
rect 24811 3349 24823 3383
rect 24765 3343 24823 3349
rect 25409 3383 25467 3389
rect 25409 3349 25421 3383
rect 25455 3380 25467 3383
rect 26234 3380 26240 3392
rect 25455 3352 26240 3380
rect 25455 3349 25467 3352
rect 25409 3343 25467 3349
rect 26234 3340 26240 3352
rect 26292 3340 26298 3392
rect 34793 3383 34851 3389
rect 34793 3349 34805 3383
rect 34839 3380 34851 3383
rect 35066 3380 35072 3392
rect 34839 3352 35072 3380
rect 34839 3349 34851 3352
rect 34793 3343 34851 3349
rect 35066 3340 35072 3352
rect 35124 3340 35130 3392
rect 39945 3383 40003 3389
rect 39945 3349 39957 3383
rect 39991 3380 40003 3383
rect 40126 3380 40132 3392
rect 39991 3352 40132 3380
rect 39991 3349 40003 3352
rect 39945 3343 40003 3349
rect 40126 3340 40132 3352
rect 40184 3340 40190 3392
rect 40589 3383 40647 3389
rect 40589 3349 40601 3383
rect 40635 3380 40647 3383
rect 41874 3380 41880 3392
rect 40635 3352 41880 3380
rect 40635 3349 40647 3352
rect 40589 3343 40647 3349
rect 41874 3340 41880 3352
rect 41932 3340 41938 3392
rect 1104 3290 48852 3312
rect 1104 3238 16880 3290
rect 16932 3238 16944 3290
rect 16996 3238 17008 3290
rect 17060 3238 17072 3290
rect 17124 3238 17136 3290
rect 17188 3238 32811 3290
rect 32863 3238 32875 3290
rect 32927 3238 32939 3290
rect 32991 3238 33003 3290
rect 33055 3238 33067 3290
rect 33119 3238 48852 3290
rect 1104 3216 48852 3238
rect 5718 3176 5724 3188
rect 5679 3148 5724 3176
rect 5718 3136 5724 3148
rect 5776 3136 5782 3188
rect 8110 3136 8116 3188
rect 8168 3176 8174 3188
rect 11790 3176 11796 3188
rect 8168 3148 9168 3176
rect 11751 3148 11796 3176
rect 8168 3136 8174 3148
rect 4614 3040 4620 3052
rect 4575 3012 4620 3040
rect 4614 3000 4620 3012
rect 4672 3000 4678 3052
rect 8220 3049 8248 3148
rect 8297 3111 8355 3117
rect 8297 3077 8309 3111
rect 8343 3108 8355 3111
rect 9033 3111 9091 3117
rect 9033 3108 9045 3111
rect 8343 3080 9045 3108
rect 8343 3077 8355 3080
rect 8297 3071 8355 3077
rect 9033 3077 9045 3080
rect 9079 3077 9091 3111
rect 9140 3108 9168 3148
rect 11790 3136 11796 3148
rect 11848 3136 11854 3188
rect 11900 3148 16574 3176
rect 11900 3108 11928 3148
rect 15286 3108 15292 3120
rect 9140 3080 11928 3108
rect 15247 3080 15292 3108
rect 9033 3071 9091 3077
rect 15286 3068 15292 3080
rect 15344 3068 15350 3120
rect 16546 3108 16574 3148
rect 18046 3136 18052 3188
rect 18104 3176 18110 3188
rect 27062 3176 27068 3188
rect 18104 3148 25820 3176
rect 27023 3148 27068 3176
rect 18104 3136 18110 3148
rect 18138 3108 18144 3120
rect 16546 3080 18144 3108
rect 18138 3068 18144 3080
rect 18196 3068 18202 3120
rect 18322 3108 18328 3120
rect 18283 3080 18328 3108
rect 18322 3068 18328 3080
rect 18380 3068 18386 3120
rect 19334 3068 19340 3120
rect 19392 3108 19398 3120
rect 24118 3108 24124 3120
rect 19392 3080 22600 3108
rect 24079 3080 24124 3108
rect 19392 3068 19398 3080
rect 5813 3043 5871 3049
rect 5813 3009 5825 3043
rect 5859 3009 5871 3043
rect 5813 3003 5871 3009
rect 6917 3043 6975 3049
rect 6917 3009 6929 3043
rect 6963 3040 6975 3043
rect 8205 3043 8263 3049
rect 6963 3012 7696 3040
rect 6963 3009 6975 3012
rect 6917 3003 6975 3009
rect 1673 2975 1731 2981
rect 1673 2941 1685 2975
rect 1719 2972 1731 2975
rect 2133 2975 2191 2981
rect 2133 2972 2145 2975
rect 1719 2944 2145 2972
rect 1719 2941 1731 2944
rect 1673 2935 1731 2941
rect 2133 2941 2145 2944
rect 2179 2941 2191 2975
rect 2314 2972 2320 2984
rect 2275 2944 2320 2972
rect 2133 2935 2191 2941
rect 2314 2932 2320 2944
rect 2372 2932 2378 2984
rect 2590 2972 2596 2984
rect 2551 2944 2596 2972
rect 2590 2932 2596 2944
rect 2648 2932 2654 2984
rect 3878 2932 3884 2984
rect 3936 2972 3942 2984
rect 5534 2972 5540 2984
rect 3936 2944 5540 2972
rect 3936 2932 3942 2944
rect 5534 2932 5540 2944
rect 5592 2932 5598 2984
rect 5828 2972 5856 3003
rect 7466 2972 7472 2984
rect 5828 2944 7472 2972
rect 7466 2932 7472 2944
rect 7524 2932 7530 2984
rect 4614 2864 4620 2916
rect 4672 2904 4678 2916
rect 6730 2904 6736 2916
rect 4672 2876 6736 2904
rect 4672 2864 4678 2876
rect 6730 2864 6736 2876
rect 6788 2864 6794 2916
rect 7668 2904 7696 3012
rect 8205 3009 8217 3043
rect 8251 3009 8263 3043
rect 11698 3040 11704 3052
rect 11659 3012 11704 3040
rect 8205 3003 8263 3009
rect 11698 3000 11704 3012
rect 11756 3000 11762 3052
rect 12621 3043 12679 3049
rect 12621 3009 12633 3043
rect 12667 3040 12679 3043
rect 12667 3012 14136 3040
rect 12667 3009 12679 3012
rect 12621 3003 12679 3009
rect 7745 2975 7803 2981
rect 7745 2941 7757 2975
rect 7791 2972 7803 2975
rect 8849 2975 8907 2981
rect 8849 2972 8861 2975
rect 7791 2944 8861 2972
rect 7791 2941 7803 2944
rect 7745 2935 7803 2941
rect 8849 2941 8861 2944
rect 8895 2941 8907 2975
rect 9306 2972 9312 2984
rect 9267 2944 9312 2972
rect 8849 2935 8907 2941
rect 9306 2932 9312 2944
rect 9364 2932 9370 2984
rect 13814 2972 13820 2984
rect 13775 2944 13820 2972
rect 13814 2932 13820 2944
rect 13872 2932 13878 2984
rect 14108 2972 14136 3012
rect 15470 3000 15476 3052
rect 15528 3040 15534 3052
rect 15933 3043 15991 3049
rect 15528 3012 15573 3040
rect 15528 3000 15534 3012
rect 15933 3009 15945 3043
rect 15979 3040 15991 3043
rect 20438 3040 20444 3052
rect 15979 3012 16574 3040
rect 20399 3012 20444 3040
rect 15979 3009 15991 3012
rect 15933 3003 15991 3009
rect 15562 2972 15568 2984
rect 14108 2944 15568 2972
rect 15562 2932 15568 2944
rect 15620 2932 15626 2984
rect 12434 2904 12440 2916
rect 7668 2876 12440 2904
rect 12434 2864 12440 2876
rect 12492 2864 12498 2916
rect 16546 2904 16574 3012
rect 20438 3000 20444 3012
rect 20496 3000 20502 3052
rect 22572 3049 22600 3080
rect 24118 3068 24124 3080
rect 24176 3068 24182 3120
rect 25792 3117 25820 3148
rect 27062 3136 27068 3148
rect 27120 3136 27126 3188
rect 39850 3176 39856 3188
rect 31036 3148 39856 3176
rect 25777 3111 25835 3117
rect 25777 3077 25789 3111
rect 25823 3077 25835 3111
rect 25777 3071 25835 3077
rect 28261 3111 28319 3117
rect 28261 3077 28273 3111
rect 28307 3108 28319 3111
rect 28997 3111 29055 3117
rect 28997 3108 29009 3111
rect 28307 3080 29009 3108
rect 28307 3077 28319 3080
rect 28261 3071 28319 3077
rect 28997 3077 29009 3080
rect 29043 3077 29055 3111
rect 28997 3071 29055 3077
rect 22557 3043 22615 3049
rect 22557 3009 22569 3043
rect 22603 3040 22615 3043
rect 23750 3040 23756 3052
rect 22603 3012 23756 3040
rect 22603 3009 22615 3012
rect 22557 3003 22615 3009
rect 23750 3000 23756 3012
rect 23808 3000 23814 3052
rect 23934 3040 23940 3052
rect 23895 3012 23940 3040
rect 23934 3000 23940 3012
rect 23992 3000 23998 3052
rect 26970 3040 26976 3052
rect 26931 3012 26976 3040
rect 26970 3000 26976 3012
rect 27028 3000 27034 3052
rect 28169 3043 28227 3049
rect 28169 3009 28181 3043
rect 28215 3009 28227 3043
rect 28810 3040 28816 3052
rect 28771 3012 28816 3040
rect 28169 3003 28227 3009
rect 17681 2975 17739 2981
rect 17681 2941 17693 2975
rect 17727 2972 17739 2975
rect 18141 2975 18199 2981
rect 18141 2972 18153 2975
rect 17727 2944 18153 2972
rect 17727 2941 17739 2944
rect 17681 2935 17739 2941
rect 18141 2941 18153 2944
rect 18187 2941 18199 2975
rect 19334 2972 19340 2984
rect 19295 2944 19340 2972
rect 18141 2935 18199 2941
rect 19334 2932 19340 2944
rect 19392 2932 19398 2984
rect 28184 2972 28212 3003
rect 28810 3000 28816 3012
rect 28868 3000 28874 3052
rect 29086 2972 29092 2984
rect 21376 2944 29092 2972
rect 21376 2904 21404 2944
rect 29086 2932 29092 2944
rect 29144 2932 29150 2984
rect 29638 2972 29644 2984
rect 29599 2944 29644 2972
rect 29638 2932 29644 2944
rect 29696 2932 29702 2984
rect 16546 2876 21404 2904
rect 22465 2907 22523 2913
rect 22465 2873 22477 2907
rect 22511 2904 22523 2907
rect 23658 2904 23664 2916
rect 22511 2876 23664 2904
rect 22511 2873 22523 2876
rect 22465 2867 22523 2873
rect 23658 2864 23664 2876
rect 23716 2864 23722 2916
rect 23750 2864 23756 2916
rect 23808 2904 23814 2916
rect 31036 2904 31064 3148
rect 39850 3136 39856 3148
rect 39908 3136 39914 3188
rect 41690 3176 41696 3188
rect 41651 3148 41696 3176
rect 41690 3136 41696 3148
rect 41748 3136 41754 3188
rect 46658 3176 46664 3188
rect 42536 3148 45554 3176
rect 46619 3148 46664 3176
rect 31481 3111 31539 3117
rect 31481 3077 31493 3111
rect 31527 3108 31539 3111
rect 32309 3111 32367 3117
rect 32309 3108 32321 3111
rect 31527 3080 32321 3108
rect 31527 3077 31539 3080
rect 31481 3071 31539 3077
rect 32309 3077 32321 3080
rect 32355 3077 32367 3111
rect 35066 3108 35072 3120
rect 35027 3080 35072 3108
rect 32309 3071 32367 3077
rect 35066 3068 35072 3080
rect 35124 3068 35130 3120
rect 35158 3068 35164 3120
rect 35216 3108 35222 3120
rect 42536 3108 42564 3148
rect 35216 3080 42564 3108
rect 35216 3068 35222 3080
rect 31386 3040 31392 3052
rect 31347 3012 31392 3040
rect 31386 3000 31392 3012
rect 31444 3000 31450 3052
rect 31570 3000 31576 3052
rect 31628 3040 31634 3052
rect 32125 3043 32183 3049
rect 32125 3040 32137 3043
rect 31628 3012 32137 3040
rect 31628 3000 31634 3012
rect 32125 3009 32137 3012
rect 32171 3009 32183 3043
rect 34882 3040 34888 3052
rect 34843 3012 34888 3040
rect 32125 3003 32183 3009
rect 34882 3000 34888 3012
rect 34940 3000 34946 3052
rect 37277 3043 37335 3049
rect 37277 3009 37289 3043
rect 37323 3040 37335 3043
rect 37366 3040 37372 3052
rect 37323 3012 37372 3040
rect 37323 3009 37335 3012
rect 37277 3003 37335 3009
rect 37366 3000 37372 3012
rect 37424 3040 37430 3052
rect 38473 3043 38531 3049
rect 38473 3040 38485 3043
rect 37424 3012 38485 3040
rect 37424 3000 37430 3012
rect 38473 3009 38485 3012
rect 38519 3009 38531 3043
rect 39114 3040 39120 3052
rect 39075 3012 39120 3040
rect 38473 3003 38531 3009
rect 39114 3000 39120 3012
rect 39172 3000 39178 3052
rect 41874 3040 41880 3052
rect 41835 3012 41880 3040
rect 41874 3000 41880 3012
rect 41932 3000 41938 3052
rect 42536 3049 42564 3080
rect 42613 3111 42671 3117
rect 42613 3077 42625 3111
rect 42659 3108 42671 3111
rect 43349 3111 43407 3117
rect 43349 3108 43361 3111
rect 42659 3080 43361 3108
rect 42659 3077 42671 3080
rect 42613 3071 42671 3077
rect 43349 3077 43361 3080
rect 43395 3077 43407 3111
rect 45526 3108 45554 3148
rect 46658 3136 46664 3148
rect 46716 3136 46722 3188
rect 45526 3080 47440 3108
rect 43349 3071 43407 3077
rect 47412 3052 47440 3080
rect 42521 3043 42579 3049
rect 42521 3009 42533 3043
rect 42567 3009 42579 3043
rect 45462 3040 45468 3052
rect 45423 3012 45468 3040
rect 42521 3003 42579 3009
rect 45462 3000 45468 3012
rect 45520 3000 45526 3052
rect 46750 3040 46756 3052
rect 46711 3012 46756 3040
rect 46750 3000 46756 3012
rect 46808 3000 46814 3052
rect 47394 3000 47400 3052
rect 47452 3040 47458 3052
rect 47581 3043 47639 3049
rect 47581 3040 47593 3043
rect 47452 3012 47593 3040
rect 47452 3000 47458 3012
rect 47581 3009 47593 3012
rect 47627 3009 47639 3043
rect 47581 3003 47639 3009
rect 33962 2972 33968 2984
rect 33923 2944 33968 2972
rect 33962 2932 33968 2944
rect 34020 2932 34026 2984
rect 36078 2972 36084 2984
rect 36039 2944 36084 2972
rect 36078 2932 36084 2944
rect 36136 2932 36142 2984
rect 38565 2975 38623 2981
rect 38565 2941 38577 2975
rect 38611 2972 38623 2975
rect 39301 2975 39359 2981
rect 39301 2972 39313 2975
rect 38611 2944 39313 2972
rect 38611 2941 38623 2944
rect 38565 2935 38623 2941
rect 39301 2941 39313 2944
rect 39347 2941 39359 2975
rect 39301 2935 39359 2941
rect 40957 2975 41015 2981
rect 40957 2941 40969 2975
rect 41003 2941 41015 2975
rect 40957 2935 41015 2941
rect 43165 2975 43223 2981
rect 43165 2941 43177 2975
rect 43211 2972 43223 2975
rect 43714 2972 43720 2984
rect 43211 2944 43720 2972
rect 43211 2941 43223 2944
rect 43165 2935 43223 2941
rect 23808 2876 31064 2904
rect 40972 2904 41000 2935
rect 43714 2932 43720 2944
rect 43772 2932 43778 2984
rect 43898 2972 43904 2984
rect 43859 2944 43904 2972
rect 43898 2932 43904 2944
rect 43956 2932 43962 2984
rect 44358 2904 44364 2916
rect 40972 2876 44364 2904
rect 23808 2864 23814 2876
rect 44358 2864 44364 2876
rect 44416 2864 44422 2916
rect 46566 2864 46572 2916
rect 46624 2904 46630 2916
rect 49602 2904 49608 2916
rect 46624 2876 49608 2904
rect 46624 2864 46630 2876
rect 49602 2864 49608 2876
rect 49660 2864 49666 2916
rect 4522 2836 4528 2848
rect 4483 2808 4528 2836
rect 4522 2796 4528 2808
rect 4580 2796 4586 2848
rect 6546 2796 6552 2848
rect 6604 2836 6610 2848
rect 6825 2839 6883 2845
rect 6825 2836 6837 2839
rect 6604 2808 6837 2836
rect 6604 2796 6610 2808
rect 6825 2805 6837 2808
rect 6871 2805 6883 2839
rect 6825 2799 6883 2805
rect 12529 2839 12587 2845
rect 12529 2805 12541 2839
rect 12575 2836 12587 2839
rect 13354 2836 13360 2848
rect 12575 2808 13360 2836
rect 12575 2805 12587 2808
rect 12529 2799 12587 2805
rect 13354 2796 13360 2808
rect 13412 2796 13418 2848
rect 16022 2836 16028 2848
rect 15983 2808 16028 2836
rect 16022 2796 16028 2808
rect 16080 2796 16086 2848
rect 16666 2836 16672 2848
rect 16627 2808 16672 2836
rect 16666 2796 16672 2808
rect 16724 2796 16730 2848
rect 20533 2839 20591 2845
rect 20533 2805 20545 2839
rect 20579 2836 20591 2839
rect 21082 2836 21088 2848
rect 20579 2808 21088 2836
rect 20579 2805 20591 2808
rect 20533 2799 20591 2805
rect 21082 2796 21088 2808
rect 21140 2796 21146 2848
rect 21266 2836 21272 2848
rect 21227 2808 21272 2836
rect 21266 2796 21272 2808
rect 21324 2796 21330 2848
rect 23201 2839 23259 2845
rect 23201 2805 23213 2839
rect 23247 2836 23259 2839
rect 23842 2836 23848 2848
rect 23247 2808 23848 2836
rect 23247 2805 23259 2808
rect 23201 2799 23259 2805
rect 23842 2796 23848 2808
rect 23900 2796 23906 2848
rect 26418 2836 26424 2848
rect 26379 2808 26424 2836
rect 26418 2796 26424 2808
rect 26476 2796 26482 2848
rect 37369 2839 37427 2845
rect 37369 2805 37381 2839
rect 37415 2836 37427 2839
rect 37458 2836 37464 2848
rect 37415 2808 37464 2836
rect 37415 2805 37427 2808
rect 37369 2799 37427 2805
rect 37458 2796 37464 2808
rect 37516 2796 37522 2848
rect 45554 2796 45560 2848
rect 45612 2836 45618 2848
rect 47670 2836 47676 2848
rect 45612 2808 45657 2836
rect 47631 2808 47676 2836
rect 45612 2796 45618 2808
rect 47670 2796 47676 2808
rect 47728 2796 47734 2848
rect 1104 2746 48852 2768
rect 1104 2694 8915 2746
rect 8967 2694 8979 2746
rect 9031 2694 9043 2746
rect 9095 2694 9107 2746
rect 9159 2694 9171 2746
rect 9223 2694 24846 2746
rect 24898 2694 24910 2746
rect 24962 2694 24974 2746
rect 25026 2694 25038 2746
rect 25090 2694 25102 2746
rect 25154 2694 40776 2746
rect 40828 2694 40840 2746
rect 40892 2694 40904 2746
rect 40956 2694 40968 2746
rect 41020 2694 41032 2746
rect 41084 2694 48852 2746
rect 1104 2672 48852 2694
rect 2314 2592 2320 2644
rect 2372 2632 2378 2644
rect 2501 2635 2559 2641
rect 2501 2632 2513 2635
rect 2372 2604 2513 2632
rect 2372 2592 2378 2604
rect 2501 2601 2513 2604
rect 2547 2601 2559 2635
rect 2501 2595 2559 2601
rect 5534 2592 5540 2644
rect 5592 2632 5598 2644
rect 37366 2632 37372 2644
rect 5592 2604 11744 2632
rect 5592 2592 5598 2604
rect 3234 2524 3240 2576
rect 3292 2564 3298 2576
rect 3292 2536 4660 2564
rect 3292 2524 3298 2536
rect 3973 2499 4031 2505
rect 3973 2465 3985 2499
rect 4019 2496 4031 2499
rect 4522 2496 4528 2508
rect 4019 2468 4528 2496
rect 4019 2465 4031 2468
rect 3973 2459 4031 2465
rect 4522 2456 4528 2468
rect 4580 2456 4586 2508
rect 4632 2505 4660 2536
rect 7742 2524 7748 2576
rect 7800 2564 7806 2576
rect 7800 2536 9444 2564
rect 7800 2524 7806 2536
rect 4617 2499 4675 2505
rect 4617 2465 4629 2499
rect 4663 2465 4675 2499
rect 4617 2459 4675 2465
rect 5810 2456 5816 2508
rect 5868 2496 5874 2508
rect 6365 2499 6423 2505
rect 6365 2496 6377 2499
rect 5868 2468 6377 2496
rect 5868 2456 5874 2468
rect 6365 2465 6377 2468
rect 6411 2465 6423 2499
rect 6546 2496 6552 2508
rect 6507 2468 6552 2496
rect 6365 2459 6423 2465
rect 6546 2456 6552 2468
rect 6604 2456 6610 2508
rect 6730 2456 6736 2508
rect 6788 2496 6794 2508
rect 6825 2499 6883 2505
rect 6825 2496 6837 2499
rect 6788 2468 6837 2496
rect 6788 2456 6794 2468
rect 6825 2465 6837 2468
rect 6871 2465 6883 2499
rect 6825 2459 6883 2465
rect 8754 2456 8760 2508
rect 8812 2496 8818 2508
rect 9416 2505 9444 2536
rect 11716 2505 11744 2604
rect 31128 2604 37372 2632
rect 12526 2524 12532 2576
rect 12584 2564 12590 2576
rect 12584 2536 13584 2564
rect 12584 2524 12590 2536
rect 8941 2499 8999 2505
rect 8941 2496 8953 2499
rect 8812 2468 8953 2496
rect 8812 2456 8818 2468
rect 8941 2465 8953 2468
rect 8987 2465 8999 2499
rect 8941 2459 8999 2465
rect 9401 2499 9459 2505
rect 9401 2465 9413 2499
rect 9447 2465 9459 2499
rect 9401 2459 9459 2465
rect 11701 2499 11759 2505
rect 11701 2465 11713 2499
rect 11747 2465 11759 2499
rect 13354 2496 13360 2508
rect 13315 2468 13360 2496
rect 11701 2459 11759 2465
rect 13354 2456 13360 2468
rect 13412 2456 13418 2508
rect 13556 2505 13584 2536
rect 13648 2536 17172 2564
rect 13541 2499 13599 2505
rect 13541 2465 13553 2499
rect 13587 2465 13599 2499
rect 13541 2459 13599 2465
rect 2593 2431 2651 2437
rect 2593 2397 2605 2431
rect 2639 2428 2651 2431
rect 2682 2428 2688 2440
rect 2639 2400 2688 2428
rect 2639 2397 2651 2400
rect 2593 2391 2651 2397
rect 2682 2388 2688 2400
rect 2740 2388 2746 2440
rect 3237 2431 3295 2437
rect 3237 2397 3249 2431
rect 3283 2428 3295 2431
rect 3789 2431 3847 2437
rect 3789 2428 3801 2431
rect 3283 2400 3801 2428
rect 3283 2397 3295 2400
rect 3237 2391 3295 2397
rect 3789 2397 3801 2400
rect 3835 2397 3847 2431
rect 3789 2391 3847 2397
rect 3510 2320 3516 2372
rect 3568 2360 3574 2372
rect 8202 2360 8208 2372
rect 3568 2332 8208 2360
rect 3568 2320 3574 2332
rect 8202 2320 8208 2332
rect 8260 2320 8266 2372
rect 8294 2320 8300 2372
rect 8352 2360 8358 2372
rect 9125 2363 9183 2369
rect 9125 2360 9137 2363
rect 8352 2332 9137 2360
rect 8352 2320 8358 2332
rect 9125 2329 9137 2332
rect 9171 2329 9183 2363
rect 9125 2323 9183 2329
rect 3418 2252 3424 2304
rect 3476 2292 3482 2304
rect 13648 2292 13676 2536
rect 14182 2496 14188 2508
rect 14143 2468 14188 2496
rect 14182 2456 14188 2468
rect 14240 2456 14246 2508
rect 14366 2496 14372 2508
rect 14327 2468 14372 2496
rect 14366 2456 14372 2468
rect 14424 2456 14430 2508
rect 14826 2496 14832 2508
rect 14787 2468 14832 2496
rect 14826 2456 14832 2468
rect 14884 2456 14890 2508
rect 16666 2496 16672 2508
rect 16627 2468 16672 2496
rect 16666 2456 16672 2468
rect 16724 2456 16730 2508
rect 17144 2505 17172 2536
rect 25866 2524 25872 2576
rect 25924 2564 25930 2576
rect 31128 2564 31156 2604
rect 37366 2592 37372 2604
rect 37424 2592 37430 2644
rect 25924 2536 31156 2564
rect 25924 2524 25930 2536
rect 17129 2499 17187 2505
rect 17129 2465 17141 2499
rect 17175 2465 17187 2499
rect 20806 2496 20812 2508
rect 20767 2468 20812 2496
rect 17129 2459 17187 2465
rect 20806 2456 20812 2468
rect 20864 2456 20870 2508
rect 21082 2496 21088 2508
rect 21043 2468 21088 2496
rect 21082 2456 21088 2468
rect 21140 2456 21146 2508
rect 21266 2496 21272 2508
rect 21227 2468 21272 2496
rect 21266 2456 21272 2468
rect 21324 2456 21330 2508
rect 22462 2496 22468 2508
rect 22423 2468 22468 2496
rect 22462 2456 22468 2468
rect 22520 2456 22526 2508
rect 23658 2496 23664 2508
rect 23619 2468 23664 2496
rect 23658 2456 23664 2468
rect 23716 2456 23722 2508
rect 23842 2496 23848 2508
rect 23803 2468 23848 2496
rect 23842 2456 23848 2468
rect 23900 2456 23906 2508
rect 26234 2456 26240 2508
rect 26292 2496 26298 2508
rect 26418 2496 26424 2508
rect 26292 2468 26337 2496
rect 26379 2468 26424 2496
rect 26292 2456 26298 2468
rect 26418 2456 26424 2468
rect 26476 2456 26482 2508
rect 28537 2499 28595 2505
rect 28537 2465 28549 2499
rect 28583 2496 28595 2499
rect 28810 2496 28816 2508
rect 28583 2468 28816 2496
rect 28583 2465 28595 2468
rect 28537 2459 28595 2465
rect 28810 2456 28816 2468
rect 28868 2456 28874 2508
rect 28994 2496 29000 2508
rect 28955 2468 29000 2496
rect 28994 2456 29000 2468
rect 29052 2456 29058 2508
rect 29086 2388 29092 2440
rect 29144 2428 29150 2440
rect 31128 2437 31156 2536
rect 31570 2524 31576 2576
rect 31628 2564 31634 2576
rect 31628 2536 32628 2564
rect 31628 2524 31634 2536
rect 31938 2456 31944 2508
rect 31996 2496 32002 2508
rect 32600 2505 32628 2536
rect 34790 2524 34796 2576
rect 34848 2564 34854 2576
rect 45738 2564 45744 2576
rect 34848 2536 34928 2564
rect 34848 2524 34854 2536
rect 32125 2499 32183 2505
rect 32125 2496 32137 2499
rect 31996 2468 32137 2496
rect 31996 2456 32002 2468
rect 32125 2465 32137 2468
rect 32171 2465 32183 2499
rect 32125 2459 32183 2465
rect 32585 2499 32643 2505
rect 32585 2465 32597 2499
rect 32631 2465 32643 2499
rect 32585 2459 32643 2465
rect 34514 2456 34520 2508
rect 34572 2496 34578 2508
rect 34900 2505 34928 2536
rect 43732 2536 45744 2564
rect 34701 2499 34759 2505
rect 34701 2496 34713 2499
rect 34572 2468 34713 2496
rect 34572 2456 34578 2468
rect 34701 2465 34713 2468
rect 34747 2465 34759 2499
rect 34701 2459 34759 2465
rect 34885 2499 34943 2505
rect 34885 2465 34897 2499
rect 34931 2465 34943 2499
rect 37274 2496 37280 2508
rect 37235 2468 37280 2496
rect 34885 2459 34943 2465
rect 37274 2456 37280 2468
rect 37332 2456 37338 2508
rect 37458 2496 37464 2508
rect 37419 2468 37464 2496
rect 37458 2456 37464 2468
rect 37516 2456 37522 2508
rect 39942 2496 39948 2508
rect 39903 2468 39948 2496
rect 39942 2456 39948 2468
rect 40000 2456 40006 2508
rect 40126 2496 40132 2508
rect 40087 2468 40132 2496
rect 40126 2456 40132 2468
rect 40184 2456 40190 2508
rect 43732 2505 43760 2536
rect 45738 2524 45744 2536
rect 45796 2524 45802 2576
rect 43717 2499 43775 2505
rect 43717 2465 43729 2499
rect 43763 2465 43775 2499
rect 43717 2459 43775 2465
rect 43806 2456 43812 2508
rect 43864 2496 43870 2508
rect 46566 2496 46572 2508
rect 43864 2468 45554 2496
rect 46527 2468 46572 2496
rect 43864 2456 43870 2468
rect 29549 2431 29607 2437
rect 29549 2428 29561 2431
rect 29144 2400 29561 2428
rect 29144 2388 29150 2400
rect 29549 2397 29561 2400
rect 29595 2397 29607 2431
rect 29549 2391 29607 2397
rect 31113 2431 31171 2437
rect 31113 2397 31125 2431
rect 31159 2397 31171 2431
rect 31113 2391 31171 2397
rect 44450 2388 44456 2440
rect 44508 2428 44514 2440
rect 45526 2428 45554 2468
rect 46566 2456 46572 2468
rect 46624 2456 46630 2508
rect 46845 2499 46903 2505
rect 46845 2465 46857 2499
rect 46891 2496 46903 2499
rect 47670 2496 47676 2508
rect 46891 2468 47676 2496
rect 46891 2465 46903 2468
rect 46845 2459 46903 2465
rect 47670 2456 47676 2468
rect 47728 2456 47734 2508
rect 45646 2428 45652 2440
rect 44508 2400 44553 2428
rect 45526 2400 45652 2428
rect 44508 2388 44514 2400
rect 45646 2388 45652 2400
rect 45704 2388 45710 2440
rect 47029 2431 47087 2437
rect 47029 2397 47041 2431
rect 47075 2428 47087 2431
rect 47581 2431 47639 2437
rect 47581 2428 47593 2431
rect 47075 2400 47593 2428
rect 47075 2397 47087 2400
rect 47029 2391 47087 2397
rect 47581 2397 47593 2400
rect 47627 2397 47639 2431
rect 47581 2391 47639 2397
rect 16022 2320 16028 2372
rect 16080 2360 16086 2372
rect 16853 2363 16911 2369
rect 16853 2360 16865 2363
rect 16080 2332 16865 2360
rect 16080 2320 16086 2332
rect 16853 2329 16865 2332
rect 16899 2329 16911 2363
rect 24578 2360 24584 2372
rect 24539 2332 24584 2360
rect 16853 2323 16911 2329
rect 24578 2320 24584 2332
rect 24636 2320 24642 2372
rect 28813 2363 28871 2369
rect 28813 2329 28825 2363
rect 28859 2360 28871 2363
rect 29641 2363 29699 2369
rect 29641 2360 29653 2363
rect 28859 2332 29653 2360
rect 28859 2329 28871 2332
rect 28813 2323 28871 2329
rect 29641 2329 29653 2332
rect 29687 2329 29699 2363
rect 29641 2323 29699 2329
rect 31205 2363 31263 2369
rect 31205 2329 31217 2363
rect 31251 2360 31263 2363
rect 32309 2363 32367 2369
rect 32309 2360 32321 2363
rect 31251 2332 32321 2360
rect 31251 2329 31263 2332
rect 31205 2323 31263 2329
rect 32309 2329 32321 2332
rect 32355 2329 32367 2363
rect 32309 2323 32367 2329
rect 36541 2363 36599 2369
rect 36541 2329 36553 2363
rect 36587 2329 36599 2363
rect 36541 2323 36599 2329
rect 39117 2363 39175 2369
rect 39117 2329 39129 2363
rect 39163 2360 39175 2363
rect 39298 2360 39304 2372
rect 39163 2332 39304 2360
rect 39163 2329 39175 2332
rect 39117 2323 39175 2329
rect 3476 2264 13676 2292
rect 36556 2292 36584 2323
rect 39298 2320 39304 2332
rect 39356 2320 39362 2372
rect 41785 2363 41843 2369
rect 41785 2329 41797 2363
rect 41831 2360 41843 2363
rect 44174 2360 44180 2372
rect 41831 2332 44180 2360
rect 41831 2329 41843 2332
rect 41785 2323 41843 2329
rect 44174 2320 44180 2332
rect 44232 2320 44238 2372
rect 44269 2363 44327 2369
rect 44269 2329 44281 2363
rect 44315 2360 44327 2363
rect 45554 2360 45560 2372
rect 44315 2332 45560 2360
rect 44315 2329 44327 2332
rect 44269 2323 44327 2329
rect 45554 2320 45560 2332
rect 45612 2320 45618 2372
rect 47670 2292 47676 2304
rect 36556 2264 47676 2292
rect 3476 2252 3482 2264
rect 47670 2252 47676 2264
rect 47728 2252 47734 2304
rect 1104 2202 48852 2224
rect 1104 2150 16880 2202
rect 16932 2150 16944 2202
rect 16996 2150 17008 2202
rect 17060 2150 17072 2202
rect 17124 2150 17136 2202
rect 17188 2150 32811 2202
rect 32863 2150 32875 2202
rect 32927 2150 32939 2202
rect 32991 2150 33003 2202
rect 33055 2150 33067 2202
rect 33119 2150 48852 2202
rect 1104 2128 48852 2150
rect 8202 2048 8208 2100
rect 8260 2088 8266 2100
rect 13814 2088 13820 2100
rect 8260 2060 13820 2088
rect 8260 2048 8266 2060
rect 13814 2048 13820 2060
rect 13872 2048 13878 2100
rect 658 1980 664 2032
rect 716 2020 722 2032
rect 24578 2020 24584 2032
rect 716 1992 24584 2020
rect 716 1980 722 1992
rect 24578 1980 24584 1992
rect 24636 1980 24642 2032
rect 20806 1912 20812 1964
rect 20864 1952 20870 1964
rect 32214 1952 32220 1964
rect 20864 1924 32220 1952
rect 20864 1912 20870 1924
rect 32214 1912 32220 1924
rect 32272 1912 32278 1964
rect 33962 1300 33968 1352
rect 34020 1340 34026 1352
rect 46658 1340 46664 1352
rect 34020 1312 46664 1340
rect 34020 1300 34026 1312
rect 46658 1300 46664 1312
rect 46716 1300 46722 1352
rect 44174 1028 44180 1080
rect 44232 1068 44238 1080
rect 46842 1068 46848 1080
rect 44232 1040 46848 1068
rect 44232 1028 44238 1040
rect 46842 1028 46848 1040
rect 46900 1028 46906 1080
<< via1 >>
rect 4620 17484 4672 17536
rect 12348 17484 12400 17536
rect 16880 17382 16932 17434
rect 16944 17382 16996 17434
rect 17008 17382 17060 17434
rect 17072 17382 17124 17434
rect 17136 17382 17188 17434
rect 32811 17382 32863 17434
rect 32875 17382 32927 17434
rect 32939 17382 32991 17434
rect 33003 17382 33055 17434
rect 33067 17382 33119 17434
rect 4068 17280 4120 17332
rect 1400 17255 1452 17264
rect 1400 17221 1409 17255
rect 1409 17221 1443 17255
rect 1443 17221 1452 17255
rect 1400 17212 1452 17221
rect 2596 17212 2648 17264
rect 8300 17212 8352 17264
rect 11612 17212 11664 17264
rect 3056 17119 3108 17128
rect 3056 17085 3065 17119
rect 3065 17085 3099 17119
rect 3099 17085 3108 17119
rect 3056 17076 3108 17085
rect 3240 17119 3292 17128
rect 3240 17085 3249 17119
rect 3249 17085 3283 17119
rect 3283 17085 3292 17119
rect 3240 17076 3292 17085
rect 5632 17119 5684 17128
rect 5632 17085 5641 17119
rect 5641 17085 5675 17119
rect 5675 17085 5684 17119
rect 5632 17076 5684 17085
rect 5816 17119 5868 17128
rect 5816 17085 5825 17119
rect 5825 17085 5859 17119
rect 5859 17085 5868 17119
rect 5816 17076 5868 17085
rect 6552 17119 6604 17128
rect 6552 17085 6561 17119
rect 6561 17085 6595 17119
rect 6595 17085 6604 17119
rect 6552 17076 6604 17085
rect 7564 17076 7616 17128
rect 7748 17119 7800 17128
rect 7748 17085 7757 17119
rect 7757 17085 7791 17119
rect 7791 17085 7800 17119
rect 7748 17076 7800 17085
rect 7932 17076 7984 17128
rect 14280 17119 14332 17128
rect 8392 17008 8444 17060
rect 14280 17085 14289 17119
rect 14289 17085 14323 17119
rect 14323 17085 14332 17119
rect 14280 17076 14332 17085
rect 18144 17280 18196 17332
rect 24492 17280 24544 17332
rect 15568 17212 15620 17264
rect 23848 17255 23900 17264
rect 23848 17221 23857 17255
rect 23857 17221 23891 17255
rect 23891 17221 23900 17255
rect 23848 17212 23900 17221
rect 18052 17076 18104 17128
rect 18512 17119 18564 17128
rect 18512 17085 18521 17119
rect 18521 17085 18555 17119
rect 18555 17085 18564 17119
rect 18512 17076 18564 17085
rect 12164 17051 12216 17060
rect 12164 17017 12173 17051
rect 12173 17017 12207 17051
rect 12207 17017 12216 17051
rect 12164 17008 12216 17017
rect 12348 17008 12400 17060
rect 19892 17008 19944 17060
rect 22192 17119 22244 17128
rect 22192 17085 22201 17119
rect 22201 17085 22235 17119
rect 22235 17085 22244 17119
rect 22192 17076 22244 17085
rect 24400 17119 24452 17128
rect 24400 17085 24409 17119
rect 24409 17085 24443 17119
rect 24443 17085 24452 17119
rect 24400 17076 24452 17085
rect 24584 17119 24636 17128
rect 24584 17085 24593 17119
rect 24593 17085 24627 17119
rect 24627 17085 24636 17119
rect 24584 17076 24636 17085
rect 24860 17119 24912 17128
rect 24860 17085 24869 17119
rect 24869 17085 24903 17119
rect 24903 17085 24912 17119
rect 24860 17076 24912 17085
rect 27160 17119 27212 17128
rect 27160 17085 27169 17119
rect 27169 17085 27203 17119
rect 27203 17085 27212 17119
rect 27160 17076 27212 17085
rect 27620 17076 27672 17128
rect 31392 17212 31444 17264
rect 39948 17212 40000 17264
rect 47032 17255 47084 17264
rect 47032 17221 47041 17255
rect 47041 17221 47075 17255
rect 47075 17221 47084 17255
rect 47032 17212 47084 17221
rect 29920 17119 29972 17128
rect 7748 16940 7800 16992
rect 15660 16940 15712 16992
rect 17132 16940 17184 16992
rect 19708 16940 19760 16992
rect 20168 16940 20220 16992
rect 29920 17085 29929 17119
rect 29929 17085 29963 17119
rect 29963 17085 29972 17119
rect 29920 17076 29972 17085
rect 30932 17119 30984 17128
rect 30932 17085 30941 17119
rect 30941 17085 30975 17119
rect 30975 17085 30984 17119
rect 30932 17076 30984 17085
rect 32128 17119 32180 17128
rect 32128 17085 32137 17119
rect 32137 17085 32171 17119
rect 32171 17085 32180 17119
rect 32128 17076 32180 17085
rect 32312 17119 32364 17128
rect 32312 17085 32321 17119
rect 32321 17085 32355 17119
rect 32355 17085 32364 17119
rect 32312 17076 32364 17085
rect 32404 17076 32456 17128
rect 34704 17119 34756 17128
rect 34704 17085 34713 17119
rect 34713 17085 34747 17119
rect 34747 17085 34756 17119
rect 34704 17076 34756 17085
rect 34888 17119 34940 17128
rect 34888 17085 34897 17119
rect 34897 17085 34931 17119
rect 34931 17085 34940 17119
rect 34888 17076 34940 17085
rect 37280 17119 37332 17128
rect 30564 17008 30616 17060
rect 33508 17008 33560 17060
rect 37280 17085 37289 17119
rect 37289 17085 37323 17119
rect 37323 17085 37332 17119
rect 37280 17076 37332 17085
rect 37464 17119 37516 17128
rect 37464 17085 37473 17119
rect 37473 17085 37507 17119
rect 37507 17085 37516 17119
rect 37464 17076 37516 17085
rect 39948 17119 40000 17128
rect 39948 17085 39957 17119
rect 39957 17085 39991 17119
rect 39991 17085 40000 17119
rect 39948 17076 40000 17085
rect 40132 17119 40184 17128
rect 40132 17085 40141 17119
rect 40141 17085 40175 17119
rect 40175 17085 40184 17119
rect 40132 17076 40184 17085
rect 40592 17119 40644 17128
rect 40592 17085 40601 17119
rect 40601 17085 40635 17119
rect 40635 17085 40644 17119
rect 40592 17076 40644 17085
rect 42156 17076 42208 17128
rect 42708 17119 42760 17128
rect 42708 17085 42717 17119
rect 42717 17085 42751 17119
rect 42751 17085 42760 17119
rect 42708 17076 42760 17085
rect 43168 17119 43220 17128
rect 43168 17085 43177 17119
rect 43177 17085 43211 17119
rect 43211 17085 43220 17119
rect 43168 17076 43220 17085
rect 44732 17076 44784 17128
rect 45376 17119 45428 17128
rect 45376 17085 45385 17119
rect 45385 17085 45419 17119
rect 45419 17085 45428 17119
rect 45376 17076 45428 17085
rect 38016 16940 38068 16992
rect 40684 16940 40736 16992
rect 47492 16940 47544 16992
rect 47768 16983 47820 16992
rect 47768 16949 47777 16983
rect 47777 16949 47811 16983
rect 47811 16949 47820 16983
rect 47768 16940 47820 16949
rect 8915 16838 8967 16890
rect 8979 16838 9031 16890
rect 9043 16838 9095 16890
rect 9107 16838 9159 16890
rect 9171 16838 9223 16890
rect 24846 16838 24898 16890
rect 24910 16838 24962 16890
rect 24974 16838 25026 16890
rect 25038 16838 25090 16890
rect 25102 16838 25154 16890
rect 40776 16838 40828 16890
rect 40840 16838 40892 16890
rect 40904 16838 40956 16890
rect 40968 16838 41020 16890
rect 41032 16838 41084 16890
rect 3240 16736 3292 16788
rect 5816 16736 5868 16788
rect 6552 16779 6604 16788
rect 6552 16745 6561 16779
rect 6561 16745 6595 16779
rect 6595 16745 6604 16779
rect 6552 16736 6604 16745
rect 7932 16736 7984 16788
rect 15568 16736 15620 16788
rect 15660 16736 15712 16788
rect 4620 16600 4672 16652
rect 7748 16600 7800 16652
rect 2412 16575 2464 16584
rect 2412 16541 2421 16575
rect 2421 16541 2455 16575
rect 2455 16541 2464 16575
rect 2412 16532 2464 16541
rect 10600 16643 10652 16652
rect 10600 16609 10609 16643
rect 10609 16609 10643 16643
rect 10643 16609 10652 16643
rect 10600 16600 10652 16609
rect 8300 16532 8352 16584
rect 12440 16575 12492 16584
rect 12440 16541 12449 16575
rect 12449 16541 12483 16575
rect 12483 16541 12492 16575
rect 12440 16532 12492 16541
rect 17132 16668 17184 16720
rect 18512 16736 18564 16788
rect 22192 16736 22244 16788
rect 24584 16736 24636 16788
rect 24676 16736 24728 16788
rect 26792 16736 26844 16788
rect 27160 16736 27212 16788
rect 29920 16736 29972 16788
rect 30564 16779 30616 16788
rect 30564 16745 30573 16779
rect 30573 16745 30607 16779
rect 30607 16745 30616 16779
rect 30564 16736 30616 16745
rect 32312 16736 32364 16788
rect 37464 16779 37516 16788
rect 37464 16745 37473 16779
rect 37473 16745 37507 16779
rect 37507 16745 37516 16779
rect 37464 16736 37516 16745
rect 39948 16736 40000 16788
rect 42156 16779 42208 16788
rect 42156 16745 42165 16779
rect 42165 16745 42199 16779
rect 42199 16745 42208 16779
rect 42156 16736 42208 16745
rect 45376 16736 45428 16788
rect 19892 16668 19944 16720
rect 16120 16643 16172 16652
rect 16120 16609 16129 16643
rect 16129 16609 16163 16643
rect 16163 16609 16172 16643
rect 16120 16600 16172 16609
rect 17960 16600 18012 16652
rect 20168 16643 20220 16652
rect 20168 16609 20177 16643
rect 20177 16609 20211 16643
rect 20211 16609 20220 16643
rect 20168 16600 20220 16609
rect 27896 16668 27948 16720
rect 18144 16532 18196 16584
rect 18236 16532 18288 16584
rect 25136 16600 25188 16652
rect 30012 16600 30064 16652
rect 40684 16668 40736 16720
rect 42432 16668 42484 16720
rect 46572 16668 46624 16720
rect 24676 16532 24728 16584
rect 25228 16575 25280 16584
rect 25228 16541 25237 16575
rect 25237 16541 25271 16575
rect 25271 16541 25280 16575
rect 25228 16532 25280 16541
rect 27068 16575 27120 16584
rect 27068 16541 27077 16575
rect 27077 16541 27111 16575
rect 27111 16541 27120 16575
rect 27528 16575 27580 16584
rect 27068 16532 27120 16541
rect 27528 16541 27537 16575
rect 27537 16541 27571 16575
rect 27571 16541 27580 16575
rect 27528 16532 27580 16541
rect 27620 16575 27672 16584
rect 27620 16541 27629 16575
rect 27629 16541 27663 16575
rect 27663 16541 27672 16575
rect 28816 16575 28868 16584
rect 27620 16532 27672 16541
rect 28816 16541 28825 16575
rect 28825 16541 28859 16575
rect 28859 16541 28868 16575
rect 28816 16532 28868 16541
rect 31300 16600 31352 16652
rect 32680 16643 32732 16652
rect 32680 16609 32689 16643
rect 32689 16609 32723 16643
rect 32723 16609 32732 16643
rect 32680 16600 32732 16609
rect 35440 16643 35492 16652
rect 35440 16609 35449 16643
rect 35449 16609 35483 16643
rect 35483 16609 35492 16643
rect 35440 16600 35492 16609
rect 43260 16600 43312 16652
rect 43812 16643 43864 16652
rect 43812 16609 43821 16643
rect 43821 16609 43855 16643
rect 43855 16609 43864 16643
rect 43812 16600 43864 16609
rect 32220 16575 32272 16584
rect 32220 16541 32229 16575
rect 32229 16541 32263 16575
rect 32263 16541 32272 16575
rect 32220 16532 32272 16541
rect 36912 16575 36964 16584
rect 36912 16541 36921 16575
rect 36921 16541 36955 16575
rect 36955 16541 36964 16575
rect 37372 16575 37424 16584
rect 36912 16532 36964 16541
rect 37372 16541 37381 16575
rect 37381 16541 37415 16575
rect 37415 16541 37424 16575
rect 37372 16532 37424 16541
rect 3056 16464 3108 16516
rect 5632 16464 5684 16516
rect 10324 16507 10376 16516
rect 10324 16473 10333 16507
rect 10333 16473 10367 16507
rect 10367 16473 10376 16507
rect 10324 16464 10376 16473
rect 14280 16464 14332 16516
rect 15752 16507 15804 16516
rect 15752 16473 15761 16507
rect 15761 16473 15795 16507
rect 15795 16473 15804 16507
rect 15752 16464 15804 16473
rect 22560 16464 22612 16516
rect 24584 16464 24636 16516
rect 32404 16507 32456 16516
rect 32404 16473 32413 16507
rect 32413 16473 32447 16507
rect 32447 16473 32456 16507
rect 32404 16464 32456 16473
rect 35256 16464 35308 16516
rect 9680 16396 9732 16448
rect 10600 16396 10652 16448
rect 33784 16396 33836 16448
rect 38936 16532 38988 16584
rect 39856 16575 39908 16584
rect 39856 16541 39865 16575
rect 39865 16541 39899 16575
rect 39899 16541 39908 16575
rect 39856 16532 39908 16541
rect 40132 16532 40184 16584
rect 43444 16464 43496 16516
rect 39120 16396 39172 16448
rect 43168 16396 43220 16448
rect 48320 16532 48372 16584
rect 47676 16464 47728 16516
rect 16880 16294 16932 16346
rect 16944 16294 16996 16346
rect 17008 16294 17060 16346
rect 17072 16294 17124 16346
rect 17136 16294 17188 16346
rect 32811 16294 32863 16346
rect 32875 16294 32927 16346
rect 32939 16294 32991 16346
rect 33003 16294 33055 16346
rect 33067 16294 33119 16346
rect 7564 16192 7616 16244
rect 10324 16235 10376 16244
rect 10324 16201 10333 16235
rect 10333 16201 10367 16235
rect 10367 16201 10376 16235
rect 10324 16192 10376 16201
rect 10232 16099 10284 16108
rect 10232 16065 10241 16099
rect 10241 16065 10275 16099
rect 10275 16065 10284 16099
rect 10232 16056 10284 16065
rect 12440 16192 12492 16244
rect 15752 16235 15804 16244
rect 15752 16201 15761 16235
rect 15761 16201 15795 16235
rect 15795 16201 15804 16235
rect 15752 16192 15804 16201
rect 24584 16235 24636 16244
rect 24584 16201 24593 16235
rect 24593 16201 24627 16235
rect 24627 16201 24636 16235
rect 24584 16192 24636 16201
rect 32404 16235 32456 16244
rect 32404 16201 32413 16235
rect 32413 16201 32447 16235
rect 32447 16201 32456 16235
rect 32404 16192 32456 16201
rect 34888 16192 34940 16244
rect 35256 16235 35308 16244
rect 35256 16201 35265 16235
rect 35265 16201 35299 16235
rect 35299 16201 35308 16235
rect 35256 16192 35308 16201
rect 42708 16192 42760 16244
rect 43444 16235 43496 16244
rect 43444 16201 43453 16235
rect 43453 16201 43487 16235
rect 43487 16201 43496 16235
rect 43444 16192 43496 16201
rect 47676 16235 47728 16244
rect 47676 16201 47685 16235
rect 47685 16201 47719 16235
rect 47719 16201 47728 16235
rect 47676 16192 47728 16201
rect 22100 16124 22152 16176
rect 15568 16056 15620 16108
rect 18236 16099 18288 16108
rect 18236 16065 18245 16099
rect 18245 16065 18279 16099
rect 18279 16065 18288 16099
rect 18236 16056 18288 16065
rect 24400 16056 24452 16108
rect 29000 16124 29052 16176
rect 45560 16124 45612 16176
rect 24676 16056 24728 16108
rect 12532 16031 12584 16040
rect 12532 15997 12541 16031
rect 12541 15997 12575 16031
rect 12575 15997 12584 16031
rect 12532 15988 12584 15997
rect 12900 16031 12952 16040
rect 12900 15997 12909 16031
rect 12909 15997 12943 16031
rect 12943 15997 12952 16031
rect 12900 15988 12952 15997
rect 18512 15988 18564 16040
rect 18696 16031 18748 16040
rect 18696 15997 18705 16031
rect 18705 15997 18739 16031
rect 18739 15997 18748 16031
rect 18696 15988 18748 15997
rect 19248 15988 19300 16040
rect 25320 16031 25372 16040
rect 25320 15997 25329 16031
rect 25329 15997 25363 16031
rect 25363 15997 25372 16031
rect 25320 15988 25372 15997
rect 19616 15920 19668 15972
rect 27068 16056 27120 16108
rect 28816 16099 28868 16108
rect 28816 16065 28825 16099
rect 28825 16065 28859 16099
rect 28859 16065 28868 16099
rect 28816 16056 28868 16065
rect 32128 16056 32180 16108
rect 32680 16056 32732 16108
rect 28448 15988 28500 16040
rect 32220 15988 32272 16040
rect 33784 16099 33836 16108
rect 33784 16065 33793 16099
rect 33793 16065 33827 16099
rect 33827 16065 33836 16099
rect 33784 16056 33836 16065
rect 34704 16056 34756 16108
rect 36912 16056 36964 16108
rect 37280 16099 37332 16108
rect 37280 16065 37289 16099
rect 37289 16065 37323 16099
rect 37323 16065 37332 16099
rect 37280 16056 37332 16065
rect 38936 16099 38988 16108
rect 38936 16065 38945 16099
rect 38945 16065 38979 16099
rect 38979 16065 38988 16099
rect 38936 16056 38988 16065
rect 42432 16056 42484 16108
rect 43168 16056 43220 16108
rect 44732 16099 44784 16108
rect 39120 16031 39172 16040
rect 39120 15997 39129 16031
rect 39129 15997 39163 16031
rect 39163 15997 39172 16031
rect 39120 15988 39172 15997
rect 42800 15988 42852 16040
rect 44732 16065 44741 16099
rect 44741 16065 44775 16099
rect 44775 16065 44784 16099
rect 44732 16056 44784 16065
rect 47308 16056 47360 16108
rect 45376 16031 45428 16040
rect 26976 15920 27028 15972
rect 28540 15920 28592 15972
rect 45376 15997 45385 16031
rect 45385 15997 45419 16031
rect 45419 15997 45428 16031
rect 45376 15988 45428 15997
rect 46848 16031 46900 16040
rect 46848 15997 46857 16031
rect 46857 15997 46891 16031
rect 46891 15997 46900 16031
rect 46848 15988 46900 15997
rect 45560 15920 45612 15972
rect 2044 15895 2096 15904
rect 2044 15861 2053 15895
rect 2053 15861 2087 15895
rect 2087 15861 2096 15895
rect 2044 15852 2096 15861
rect 11704 15895 11756 15904
rect 11704 15861 11713 15895
rect 11713 15861 11747 15895
rect 11747 15861 11756 15895
rect 11704 15852 11756 15861
rect 16120 15852 16172 15904
rect 25412 15852 25464 15904
rect 35624 15852 35676 15904
rect 41236 15895 41288 15904
rect 41236 15861 41245 15895
rect 41245 15861 41279 15895
rect 41279 15861 41288 15895
rect 41236 15852 41288 15861
rect 8915 15750 8967 15802
rect 8979 15750 9031 15802
rect 9043 15750 9095 15802
rect 9107 15750 9159 15802
rect 9171 15750 9223 15802
rect 24846 15750 24898 15802
rect 24910 15750 24962 15802
rect 24974 15750 25026 15802
rect 25038 15750 25090 15802
rect 25102 15750 25154 15802
rect 40776 15750 40828 15802
rect 40840 15750 40892 15802
rect 40904 15750 40956 15802
rect 40968 15750 41020 15802
rect 41032 15750 41084 15802
rect 18512 15691 18564 15700
rect 18512 15657 18521 15691
rect 18521 15657 18555 15691
rect 18555 15657 18564 15691
rect 18512 15648 18564 15657
rect 28448 15691 28500 15700
rect 28448 15657 28457 15691
rect 28457 15657 28491 15691
rect 28491 15657 28500 15691
rect 28448 15648 28500 15657
rect 28540 15648 28592 15700
rect 42800 15648 42852 15700
rect 43260 15691 43312 15700
rect 43260 15657 43269 15691
rect 43269 15657 43303 15691
rect 43303 15657 43312 15691
rect 43260 15648 43312 15657
rect 45376 15648 45428 15700
rect 15568 15580 15620 15632
rect 22100 15580 22152 15632
rect 11704 15555 11756 15564
rect 11704 15521 11713 15555
rect 11713 15521 11747 15555
rect 11747 15521 11756 15555
rect 11704 15512 11756 15521
rect 12256 15512 12308 15564
rect 16120 15555 16172 15564
rect 16120 15521 16129 15555
rect 16129 15521 16163 15555
rect 16163 15521 16172 15555
rect 16120 15512 16172 15521
rect 16764 15555 16816 15564
rect 16764 15521 16773 15555
rect 16773 15521 16807 15555
rect 16807 15521 16816 15555
rect 16764 15512 16816 15521
rect 25228 15555 25280 15564
rect 2412 15444 2464 15496
rect 15660 15487 15712 15496
rect 15660 15453 15669 15487
rect 15669 15453 15703 15487
rect 15703 15453 15712 15487
rect 15660 15444 15712 15453
rect 18420 15444 18472 15496
rect 19248 15444 19300 15496
rect 19892 15487 19944 15496
rect 19892 15453 19901 15487
rect 19901 15453 19935 15487
rect 19935 15453 19944 15487
rect 19892 15444 19944 15453
rect 11888 15419 11940 15428
rect 11888 15385 11897 15419
rect 11897 15385 11931 15419
rect 11931 15385 11940 15419
rect 11888 15376 11940 15385
rect 19432 15419 19484 15428
rect 19432 15385 19441 15419
rect 19441 15385 19475 15419
rect 19475 15385 19484 15419
rect 25228 15521 25237 15555
rect 25237 15521 25271 15555
rect 25271 15521 25280 15555
rect 25228 15512 25280 15521
rect 25412 15555 25464 15564
rect 25412 15521 25421 15555
rect 25421 15521 25455 15555
rect 25455 15521 25464 15555
rect 25412 15512 25464 15521
rect 25780 15555 25832 15564
rect 25780 15521 25789 15555
rect 25789 15521 25823 15555
rect 25823 15521 25832 15555
rect 25780 15512 25832 15521
rect 35624 15555 35676 15564
rect 35624 15521 35633 15555
rect 35633 15521 35667 15555
rect 35667 15521 35676 15555
rect 35624 15512 35676 15521
rect 36084 15555 36136 15564
rect 36084 15521 36093 15555
rect 36093 15521 36127 15555
rect 36127 15521 36136 15555
rect 36084 15512 36136 15521
rect 41236 15512 41288 15564
rect 41880 15555 41932 15564
rect 41880 15521 41889 15555
rect 41889 15521 41923 15555
rect 41923 15521 41932 15555
rect 41880 15512 41932 15521
rect 27712 15444 27764 15496
rect 40132 15444 40184 15496
rect 46756 15555 46808 15564
rect 46756 15521 46765 15555
rect 46765 15521 46799 15555
rect 46799 15521 46808 15555
rect 46756 15512 46808 15521
rect 47768 15512 47820 15564
rect 24584 15419 24636 15428
rect 19432 15376 19484 15385
rect 24584 15385 24593 15419
rect 24593 15385 24627 15419
rect 24627 15385 24636 15419
rect 24584 15376 24636 15385
rect 35900 15376 35952 15428
rect 47952 15419 48004 15428
rect 47952 15385 47961 15419
rect 47961 15385 47995 15419
rect 47995 15385 48004 15419
rect 47952 15376 48004 15385
rect 2228 15308 2280 15360
rect 24676 15351 24728 15360
rect 24676 15317 24685 15351
rect 24685 15317 24719 15351
rect 24719 15317 24728 15351
rect 24676 15308 24728 15317
rect 16880 15206 16932 15258
rect 16944 15206 16996 15258
rect 17008 15206 17060 15258
rect 17072 15206 17124 15258
rect 17136 15206 17188 15258
rect 32811 15206 32863 15258
rect 32875 15206 32927 15258
rect 32939 15206 32991 15258
rect 33003 15206 33055 15258
rect 33067 15206 33119 15258
rect 11888 15147 11940 15156
rect 11888 15113 11897 15147
rect 11897 15113 11931 15147
rect 11931 15113 11940 15147
rect 11888 15104 11940 15113
rect 12532 15147 12584 15156
rect 12532 15113 12541 15147
rect 12541 15113 12575 15147
rect 12575 15113 12584 15147
rect 12532 15104 12584 15113
rect 17960 15104 18012 15156
rect 18328 15104 18380 15156
rect 27528 15104 27580 15156
rect 27620 15104 27672 15156
rect 33784 15104 33836 15156
rect 35900 15147 35952 15156
rect 35900 15113 35909 15147
rect 35909 15113 35943 15147
rect 35943 15113 35952 15147
rect 35900 15104 35952 15113
rect 47952 15104 48004 15156
rect 2228 15079 2280 15088
rect 2228 15045 2237 15079
rect 2237 15045 2271 15079
rect 2271 15045 2280 15079
rect 2228 15036 2280 15045
rect 18052 15036 18104 15088
rect 25872 15079 25924 15088
rect 25872 15045 25881 15079
rect 25881 15045 25915 15079
rect 25915 15045 25924 15079
rect 25872 15036 25924 15045
rect 2044 15011 2096 15020
rect 2044 14977 2053 15011
rect 2053 14977 2087 15011
rect 2087 14977 2096 15011
rect 2044 14968 2096 14977
rect 11796 15011 11848 15020
rect 11796 14977 11805 15011
rect 11805 14977 11839 15011
rect 11839 14977 11848 15011
rect 11796 14968 11848 14977
rect 12440 15011 12492 15020
rect 12440 14977 12449 15011
rect 12449 14977 12483 15011
rect 12483 14977 12492 15011
rect 12440 14968 12492 14977
rect 18512 15011 18564 15020
rect 18512 14977 18521 15011
rect 18521 14977 18555 15011
rect 18555 14977 18564 15011
rect 18512 14968 18564 14977
rect 19892 14968 19944 15020
rect 24676 15011 24728 15020
rect 24676 14977 24685 15011
rect 24685 14977 24719 15011
rect 24719 14977 24728 15011
rect 24676 14968 24728 14977
rect 25228 14968 25280 15020
rect 2780 14943 2832 14952
rect 2780 14909 2789 14943
rect 2789 14909 2823 14943
rect 2823 14909 2832 14943
rect 2780 14900 2832 14909
rect 15660 14900 15712 14952
rect 11796 14832 11848 14884
rect 18328 14943 18380 14952
rect 18328 14909 18337 14943
rect 18337 14909 18371 14943
rect 18371 14909 18380 14943
rect 19708 14943 19760 14952
rect 18328 14900 18380 14909
rect 19708 14909 19717 14943
rect 19717 14909 19751 14943
rect 19751 14909 19760 14943
rect 19708 14900 19760 14909
rect 20628 14943 20680 14952
rect 20628 14909 20637 14943
rect 20637 14909 20671 14943
rect 20671 14909 20680 14943
rect 20628 14900 20680 14909
rect 24492 14943 24544 14952
rect 24492 14909 24501 14943
rect 24501 14909 24535 14943
rect 24535 14909 24544 14943
rect 24492 14900 24544 14909
rect 24584 14900 24636 14952
rect 31668 14968 31720 15020
rect 35992 15011 36044 15020
rect 35992 14977 36001 15011
rect 36001 14977 36035 15011
rect 36035 14977 36044 15011
rect 35992 14968 36044 14977
rect 45560 15011 45612 15020
rect 45560 14977 45569 15011
rect 45569 14977 45603 15011
rect 45603 14977 45612 15011
rect 45560 14968 45612 14977
rect 46756 14968 46808 15020
rect 27804 14900 27856 14952
rect 12440 14764 12492 14816
rect 18052 14764 18104 14816
rect 29092 14832 29144 14884
rect 20628 14764 20680 14816
rect 24492 14764 24544 14816
rect 27620 14764 27672 14816
rect 27712 14764 27764 14816
rect 32680 14900 32732 14952
rect 46940 14900 46992 14952
rect 31484 14764 31536 14816
rect 46296 14764 46348 14816
rect 46480 14764 46532 14816
rect 8915 14662 8967 14714
rect 8979 14662 9031 14714
rect 9043 14662 9095 14714
rect 9107 14662 9159 14714
rect 9171 14662 9223 14714
rect 24846 14662 24898 14714
rect 24910 14662 24962 14714
rect 24974 14662 25026 14714
rect 25038 14662 25090 14714
rect 25102 14662 25154 14714
rect 40776 14662 40828 14714
rect 40840 14662 40892 14714
rect 40904 14662 40956 14714
rect 40968 14662 41020 14714
rect 41032 14662 41084 14714
rect 18512 14603 18564 14612
rect 18512 14569 18521 14603
rect 18521 14569 18555 14603
rect 18555 14569 18564 14603
rect 18512 14560 18564 14569
rect 2044 14356 2096 14408
rect 2688 14356 2740 14408
rect 7748 14356 7800 14408
rect 19616 14467 19668 14476
rect 19616 14433 19625 14467
rect 19625 14433 19659 14467
rect 19659 14433 19668 14467
rect 19616 14424 19668 14433
rect 39856 14424 39908 14476
rect 46296 14467 46348 14476
rect 46296 14433 46305 14467
rect 46305 14433 46339 14467
rect 46339 14433 46348 14467
rect 46296 14424 46348 14433
rect 46480 14467 46532 14476
rect 46480 14433 46489 14467
rect 46489 14433 46523 14467
rect 46523 14433 46532 14467
rect 46480 14424 46532 14433
rect 48136 14467 48188 14476
rect 48136 14433 48145 14467
rect 48145 14433 48179 14467
rect 48179 14433 48188 14467
rect 48136 14424 48188 14433
rect 25228 14399 25280 14408
rect 25228 14365 25237 14399
rect 25237 14365 25271 14399
rect 25271 14365 25280 14399
rect 25228 14356 25280 14365
rect 25780 14356 25832 14408
rect 26976 14399 27028 14408
rect 12164 14288 12216 14340
rect 2228 14220 2280 14272
rect 24584 14220 24636 14272
rect 26976 14365 26985 14399
rect 26985 14365 27019 14399
rect 27019 14365 27028 14399
rect 26976 14356 27028 14365
rect 31392 14399 31444 14408
rect 31392 14365 31401 14399
rect 31401 14365 31435 14399
rect 31435 14365 31444 14399
rect 31392 14356 31444 14365
rect 31668 14399 31720 14408
rect 31668 14365 31677 14399
rect 31677 14365 31711 14399
rect 31711 14365 31720 14399
rect 31668 14356 31720 14365
rect 45192 14356 45244 14408
rect 27804 14331 27856 14340
rect 27804 14297 27813 14331
rect 27813 14297 27847 14331
rect 27847 14297 27856 14331
rect 27804 14288 27856 14297
rect 27988 14331 28040 14340
rect 27988 14297 27997 14331
rect 27997 14297 28031 14331
rect 28031 14297 28040 14331
rect 27988 14288 28040 14297
rect 33232 14288 33284 14340
rect 35992 14220 36044 14272
rect 16880 14118 16932 14170
rect 16944 14118 16996 14170
rect 17008 14118 17060 14170
rect 17072 14118 17124 14170
rect 17136 14118 17188 14170
rect 32811 14118 32863 14170
rect 32875 14118 32927 14170
rect 32939 14118 32991 14170
rect 33003 14118 33055 14170
rect 33067 14118 33119 14170
rect 2228 13991 2280 14000
rect 2228 13957 2237 13991
rect 2237 13957 2271 13991
rect 2271 13957 2280 13991
rect 2228 13948 2280 13957
rect 27896 13948 27948 14000
rect 2044 13923 2096 13932
rect 2044 13889 2053 13923
rect 2053 13889 2087 13923
rect 2087 13889 2096 13923
rect 2044 13880 2096 13889
rect 25228 13923 25280 13932
rect 25228 13889 25237 13923
rect 25237 13889 25271 13923
rect 25271 13889 25280 13923
rect 25228 13880 25280 13889
rect 27988 13880 28040 13932
rect 2780 13855 2832 13864
rect 2780 13821 2789 13855
rect 2789 13821 2823 13855
rect 2823 13821 2832 13855
rect 2780 13812 2832 13821
rect 10232 13812 10284 13864
rect 30012 13880 30064 13932
rect 34704 13880 34756 13932
rect 45192 13923 45244 13932
rect 45192 13889 45201 13923
rect 45201 13889 45235 13923
rect 45235 13889 45244 13923
rect 45192 13880 45244 13889
rect 47032 13880 47084 13932
rect 29000 13855 29052 13864
rect 29000 13821 29009 13855
rect 29009 13821 29043 13855
rect 29043 13821 29052 13855
rect 29000 13812 29052 13821
rect 31392 13812 31444 13864
rect 46848 13855 46900 13864
rect 46848 13821 46857 13855
rect 46857 13821 46891 13855
rect 46891 13821 46900 13855
rect 46848 13812 46900 13821
rect 8915 13574 8967 13626
rect 8979 13574 9031 13626
rect 9043 13574 9095 13626
rect 9107 13574 9159 13626
rect 9171 13574 9223 13626
rect 24846 13574 24898 13626
rect 24910 13574 24962 13626
rect 24974 13574 25026 13626
rect 25038 13574 25090 13626
rect 25102 13574 25154 13626
rect 40776 13574 40828 13626
rect 40840 13574 40892 13626
rect 40904 13574 40956 13626
rect 40968 13574 41020 13626
rect 41032 13574 41084 13626
rect 26792 13336 26844 13388
rect 27436 13336 27488 13388
rect 2044 13268 2096 13320
rect 3792 13311 3844 13320
rect 3792 13277 3801 13311
rect 3801 13277 3835 13311
rect 3835 13277 3844 13311
rect 3792 13268 3844 13277
rect 27620 13268 27672 13320
rect 27988 13268 28040 13320
rect 27436 13200 27488 13252
rect 36544 13132 36596 13184
rect 37372 13132 37424 13184
rect 48136 13243 48188 13252
rect 48136 13209 48145 13243
rect 48145 13209 48179 13243
rect 48179 13209 48188 13243
rect 48136 13200 48188 13209
rect 46940 13132 46992 13184
rect 16880 13030 16932 13082
rect 16944 13030 16996 13082
rect 17008 13030 17060 13082
rect 17072 13030 17124 13082
rect 17136 13030 17188 13082
rect 32811 13030 32863 13082
rect 32875 13030 32927 13082
rect 32939 13030 32991 13082
rect 33003 13030 33055 13082
rect 33067 13030 33119 13082
rect 2044 12835 2096 12844
rect 2044 12801 2053 12835
rect 2053 12801 2087 12835
rect 2087 12801 2096 12835
rect 2044 12792 2096 12801
rect 27620 12835 27672 12844
rect 27620 12801 27629 12835
rect 27629 12801 27663 12835
rect 27663 12801 27672 12835
rect 27620 12792 27672 12801
rect 47492 12792 47544 12844
rect 2228 12767 2280 12776
rect 2228 12733 2237 12767
rect 2237 12733 2271 12767
rect 2271 12733 2280 12767
rect 2228 12724 2280 12733
rect 2780 12767 2832 12776
rect 2780 12733 2789 12767
rect 2789 12733 2823 12767
rect 2823 12733 2832 12767
rect 27344 12767 27396 12776
rect 2780 12724 2832 12733
rect 27344 12733 27353 12767
rect 27353 12733 27387 12767
rect 27387 12733 27396 12767
rect 27344 12724 27396 12733
rect 42340 12724 42392 12776
rect 45192 12767 45244 12776
rect 45192 12733 45201 12767
rect 45201 12733 45235 12767
rect 45235 12733 45244 12767
rect 45192 12724 45244 12733
rect 46848 12767 46900 12776
rect 46848 12733 46857 12767
rect 46857 12733 46891 12767
rect 46891 12733 46900 12767
rect 46848 12724 46900 12733
rect 32680 12656 32732 12708
rect 47492 12656 47544 12708
rect 8915 12486 8967 12538
rect 8979 12486 9031 12538
rect 9043 12486 9095 12538
rect 9107 12486 9159 12538
rect 9171 12486 9223 12538
rect 24846 12486 24898 12538
rect 24910 12486 24962 12538
rect 24974 12486 25026 12538
rect 25038 12486 25090 12538
rect 25102 12486 25154 12538
rect 40776 12486 40828 12538
rect 40840 12486 40892 12538
rect 40904 12486 40956 12538
rect 40968 12486 41020 12538
rect 41032 12486 41084 12538
rect 2228 12384 2280 12436
rect 45192 12384 45244 12436
rect 3792 12291 3844 12300
rect 3792 12257 3801 12291
rect 3801 12257 3835 12291
rect 3835 12257 3844 12291
rect 3792 12248 3844 12257
rect 4068 12248 4120 12300
rect 47584 12291 47636 12300
rect 47584 12257 47593 12291
rect 47593 12257 47627 12291
rect 47627 12257 47636 12291
rect 47584 12248 47636 12257
rect 2596 12223 2648 12232
rect 2596 12189 2605 12223
rect 2605 12189 2639 12223
rect 2639 12189 2648 12223
rect 2596 12180 2648 12189
rect 3976 12155 4028 12164
rect 3976 12121 3985 12155
rect 3985 12121 4019 12155
rect 4019 12121 4028 12155
rect 3976 12112 4028 12121
rect 47676 12112 47728 12164
rect 16880 11942 16932 11994
rect 16944 11942 16996 11994
rect 17008 11942 17060 11994
rect 17072 11942 17124 11994
rect 17136 11942 17188 11994
rect 32811 11942 32863 11994
rect 32875 11942 32927 11994
rect 32939 11942 32991 11994
rect 33003 11942 33055 11994
rect 33067 11942 33119 11994
rect 3976 11840 4028 11892
rect 47676 11883 47728 11892
rect 47676 11849 47685 11883
rect 47685 11849 47719 11883
rect 47719 11849 47728 11883
rect 47676 11840 47728 11849
rect 8208 11704 8260 11756
rect 27344 11704 27396 11756
rect 47400 11704 47452 11756
rect 46572 11636 46624 11688
rect 46848 11679 46900 11688
rect 46848 11645 46857 11679
rect 46857 11645 46891 11679
rect 46891 11645 46900 11679
rect 46848 11636 46900 11645
rect 8915 11398 8967 11450
rect 8979 11398 9031 11450
rect 9043 11398 9095 11450
rect 9107 11398 9159 11450
rect 9171 11398 9223 11450
rect 24846 11398 24898 11450
rect 24910 11398 24962 11450
rect 24974 11398 25026 11450
rect 25038 11398 25090 11450
rect 25102 11398 25154 11450
rect 40776 11398 40828 11450
rect 40840 11398 40892 11450
rect 40904 11398 40956 11450
rect 40968 11398 41020 11450
rect 41032 11398 41084 11450
rect 2044 11092 2096 11144
rect 47676 11024 47728 11076
rect 48136 11067 48188 11076
rect 48136 11033 48145 11067
rect 48145 11033 48179 11067
rect 48179 11033 48188 11067
rect 48136 11024 48188 11033
rect 16880 10854 16932 10906
rect 16944 10854 16996 10906
rect 17008 10854 17060 10906
rect 17072 10854 17124 10906
rect 17136 10854 17188 10906
rect 32811 10854 32863 10906
rect 32875 10854 32927 10906
rect 32939 10854 32991 10906
rect 33003 10854 33055 10906
rect 33067 10854 33119 10906
rect 46572 10795 46624 10804
rect 46572 10761 46581 10795
rect 46581 10761 46615 10795
rect 46615 10761 46624 10795
rect 46572 10752 46624 10761
rect 47676 10795 47728 10804
rect 47676 10761 47685 10795
rect 47685 10761 47719 10795
rect 47719 10761 47728 10795
rect 47676 10752 47728 10761
rect 2044 10659 2096 10668
rect 2044 10625 2053 10659
rect 2053 10625 2087 10659
rect 2087 10625 2096 10659
rect 2044 10616 2096 10625
rect 46664 10659 46716 10668
rect 46664 10625 46673 10659
rect 46673 10625 46707 10659
rect 46707 10625 46716 10659
rect 46664 10616 46716 10625
rect 47032 10616 47084 10668
rect 47400 10616 47452 10668
rect 2504 10548 2556 10600
rect 2780 10591 2832 10600
rect 2780 10557 2789 10591
rect 2789 10557 2823 10591
rect 2823 10557 2832 10591
rect 2780 10548 2832 10557
rect 11060 10412 11112 10464
rect 12992 10455 13044 10464
rect 12992 10421 13001 10455
rect 13001 10421 13035 10455
rect 13035 10421 13044 10455
rect 12992 10412 13044 10421
rect 46296 10412 46348 10464
rect 8915 10310 8967 10362
rect 8979 10310 9031 10362
rect 9043 10310 9095 10362
rect 9107 10310 9159 10362
rect 9171 10310 9223 10362
rect 24846 10310 24898 10362
rect 24910 10310 24962 10362
rect 24974 10310 25026 10362
rect 25038 10310 25090 10362
rect 25102 10310 25154 10362
rect 40776 10310 40828 10362
rect 40840 10310 40892 10362
rect 40904 10310 40956 10362
rect 40968 10310 41020 10362
rect 41032 10310 41084 10362
rect 2504 10251 2556 10260
rect 2504 10217 2513 10251
rect 2513 10217 2547 10251
rect 2547 10217 2556 10251
rect 2504 10208 2556 10217
rect 2688 10004 2740 10056
rect 3424 9936 3476 9988
rect 11060 10115 11112 10124
rect 11060 10081 11069 10115
rect 11069 10081 11103 10115
rect 11103 10081 11112 10115
rect 11060 10072 11112 10081
rect 46296 10115 46348 10124
rect 46296 10081 46305 10115
rect 46305 10081 46339 10115
rect 46339 10081 46348 10115
rect 46296 10072 46348 10081
rect 48136 10115 48188 10124
rect 48136 10081 48145 10115
rect 48145 10081 48179 10115
rect 48179 10081 48188 10115
rect 48136 10072 48188 10081
rect 18328 10004 18380 10056
rect 40040 10047 40092 10056
rect 40040 10013 40049 10047
rect 40049 10013 40083 10047
rect 40083 10013 40092 10047
rect 40040 10004 40092 10013
rect 11244 9979 11296 9988
rect 11244 9945 11253 9979
rect 11253 9945 11287 9979
rect 11287 9945 11296 9979
rect 11244 9936 11296 9945
rect 47676 9936 47728 9988
rect 13176 9868 13228 9920
rect 16880 9766 16932 9818
rect 16944 9766 16996 9818
rect 17008 9766 17060 9818
rect 17072 9766 17124 9818
rect 17136 9766 17188 9818
rect 32811 9766 32863 9818
rect 32875 9766 32927 9818
rect 32939 9766 32991 9818
rect 33003 9766 33055 9818
rect 33067 9766 33119 9818
rect 11244 9664 11296 9716
rect 13176 9639 13228 9648
rect 13176 9605 13185 9639
rect 13185 9605 13219 9639
rect 13219 9605 13228 9639
rect 13176 9596 13228 9605
rect 25320 9596 25372 9648
rect 47676 9639 47728 9648
rect 11796 9528 11848 9580
rect 12992 9571 13044 9580
rect 12992 9537 13001 9571
rect 13001 9537 13035 9571
rect 13035 9537 13044 9571
rect 12992 9528 13044 9537
rect 40040 9571 40092 9580
rect 40040 9537 40049 9571
rect 40049 9537 40083 9571
rect 40083 9537 40092 9571
rect 40040 9528 40092 9537
rect 47676 9605 47685 9639
rect 47685 9605 47719 9639
rect 47719 9605 47728 9639
rect 47676 9596 47728 9605
rect 47584 9571 47636 9580
rect 47584 9537 47593 9571
rect 47593 9537 47627 9571
rect 47627 9537 47636 9571
rect 47584 9528 47636 9537
rect 13544 9503 13596 9512
rect 13544 9469 13553 9503
rect 13553 9469 13587 9503
rect 13587 9469 13596 9503
rect 13544 9460 13596 9469
rect 40224 9503 40276 9512
rect 40224 9469 40233 9503
rect 40233 9469 40267 9503
rect 40267 9469 40276 9503
rect 40224 9460 40276 9469
rect 40592 9503 40644 9512
rect 40592 9469 40601 9503
rect 40601 9469 40635 9503
rect 40635 9469 40644 9503
rect 40592 9460 40644 9469
rect 8915 9222 8967 9274
rect 8979 9222 9031 9274
rect 9043 9222 9095 9274
rect 9107 9222 9159 9274
rect 9171 9222 9223 9274
rect 24846 9222 24898 9274
rect 24910 9222 24962 9274
rect 24974 9222 25026 9274
rect 25038 9222 25090 9274
rect 25102 9222 25154 9274
rect 40776 9222 40828 9274
rect 40840 9222 40892 9274
rect 40904 9222 40956 9274
rect 40968 9222 41020 9274
rect 41032 9222 41084 9274
rect 40224 9120 40276 9172
rect 2044 8959 2096 8968
rect 2044 8925 2053 8959
rect 2053 8925 2087 8959
rect 2087 8925 2096 8959
rect 2044 8916 2096 8925
rect 20628 8916 20680 8968
rect 46664 8916 46716 8968
rect 16880 8678 16932 8730
rect 16944 8678 16996 8730
rect 17008 8678 17060 8730
rect 17072 8678 17124 8730
rect 17136 8678 17188 8730
rect 32811 8678 32863 8730
rect 32875 8678 32927 8730
rect 32939 8678 32991 8730
rect 33003 8678 33055 8730
rect 33067 8678 33119 8730
rect 2044 8483 2096 8492
rect 2044 8449 2053 8483
rect 2053 8449 2087 8483
rect 2087 8449 2096 8483
rect 2044 8440 2096 8449
rect 2228 8415 2280 8424
rect 2228 8381 2237 8415
rect 2237 8381 2271 8415
rect 2271 8381 2280 8415
rect 2228 8372 2280 8381
rect 2780 8415 2832 8424
rect 2780 8381 2789 8415
rect 2789 8381 2823 8415
rect 2823 8381 2832 8415
rect 2780 8372 2832 8381
rect 10324 8236 10376 8288
rect 8915 8134 8967 8186
rect 8979 8134 9031 8186
rect 9043 8134 9095 8186
rect 9107 8134 9159 8186
rect 9171 8134 9223 8186
rect 24846 8134 24898 8186
rect 24910 8134 24962 8186
rect 24974 8134 25026 8186
rect 25038 8134 25090 8186
rect 25102 8134 25154 8186
rect 40776 8134 40828 8186
rect 40840 8134 40892 8186
rect 40904 8134 40956 8186
rect 40968 8134 41020 8186
rect 41032 8134 41084 8186
rect 2228 8032 2280 8084
rect 10324 7939 10376 7948
rect 10324 7905 10333 7939
rect 10333 7905 10367 7939
rect 10367 7905 10376 7939
rect 10324 7896 10376 7905
rect 10968 7939 11020 7948
rect 10968 7905 10977 7939
rect 10977 7905 11011 7939
rect 11011 7905 11020 7939
rect 10968 7896 11020 7905
rect 2412 7871 2464 7880
rect 2412 7837 2421 7871
rect 2421 7837 2455 7871
rect 2455 7837 2464 7871
rect 2412 7828 2464 7837
rect 17684 7871 17736 7880
rect 17684 7837 17693 7871
rect 17693 7837 17727 7871
rect 17727 7837 17736 7871
rect 17684 7828 17736 7837
rect 29736 7828 29788 7880
rect 33232 7871 33284 7880
rect 33232 7837 33241 7871
rect 33241 7837 33275 7871
rect 33275 7837 33284 7871
rect 33232 7828 33284 7837
rect 10508 7803 10560 7812
rect 10508 7769 10517 7803
rect 10517 7769 10551 7803
rect 10551 7769 10560 7803
rect 10508 7760 10560 7769
rect 33876 7692 33928 7744
rect 16880 7590 16932 7642
rect 16944 7590 16996 7642
rect 17008 7590 17060 7642
rect 17072 7590 17124 7642
rect 17136 7590 17188 7642
rect 32811 7590 32863 7642
rect 32875 7590 32927 7642
rect 32939 7590 32991 7642
rect 33003 7590 33055 7642
rect 33067 7590 33119 7642
rect 10508 7531 10560 7540
rect 10508 7497 10517 7531
rect 10517 7497 10551 7531
rect 10551 7497 10560 7531
rect 10508 7488 10560 7497
rect 33876 7463 33928 7472
rect 33876 7429 33885 7463
rect 33885 7429 33919 7463
rect 33919 7429 33928 7463
rect 33876 7420 33928 7429
rect 10416 7395 10468 7404
rect 10416 7361 10425 7395
rect 10425 7361 10459 7395
rect 10459 7361 10468 7395
rect 10416 7352 10468 7361
rect 17684 7395 17736 7404
rect 17684 7361 17693 7395
rect 17693 7361 17727 7395
rect 17727 7361 17736 7395
rect 17684 7352 17736 7361
rect 29092 7395 29144 7404
rect 29092 7361 29101 7395
rect 29101 7361 29135 7395
rect 29135 7361 29144 7395
rect 29092 7352 29144 7361
rect 29736 7395 29788 7404
rect 29736 7361 29745 7395
rect 29745 7361 29779 7395
rect 29779 7361 29788 7395
rect 29736 7352 29788 7361
rect 18052 7284 18104 7336
rect 33692 7327 33744 7336
rect 3424 7216 3476 7268
rect 33692 7293 33701 7327
rect 33701 7293 33735 7327
rect 33735 7293 33744 7327
rect 33692 7284 33744 7293
rect 34612 7327 34664 7336
rect 34612 7293 34621 7327
rect 34621 7293 34655 7327
rect 34655 7293 34664 7327
rect 34612 7284 34664 7293
rect 46756 7284 46808 7336
rect 2136 7148 2188 7200
rect 8915 7046 8967 7098
rect 8979 7046 9031 7098
rect 9043 7046 9095 7098
rect 9107 7046 9159 7098
rect 9171 7046 9223 7098
rect 24846 7046 24898 7098
rect 24910 7046 24962 7098
rect 24974 7046 25026 7098
rect 25038 7046 25090 7098
rect 25102 7046 25154 7098
rect 40776 7046 40828 7098
rect 40840 7046 40892 7098
rect 40904 7046 40956 7098
rect 40968 7046 41020 7098
rect 41032 7046 41084 7098
rect 33692 6987 33744 6996
rect 33692 6953 33701 6987
rect 33701 6953 33735 6987
rect 33735 6953 33744 6987
rect 33692 6944 33744 6953
rect 18052 6808 18104 6860
rect 2688 6783 2740 6792
rect 2688 6749 2697 6783
rect 2697 6749 2731 6783
rect 2731 6749 2740 6783
rect 2688 6740 2740 6749
rect 18420 6740 18472 6792
rect 46296 6740 46348 6792
rect 48136 6740 48188 6792
rect 2320 6604 2372 6656
rect 16880 6502 16932 6554
rect 16944 6502 16996 6554
rect 17008 6502 17060 6554
rect 17072 6502 17124 6554
rect 17136 6502 17188 6554
rect 32811 6502 32863 6554
rect 32875 6502 32927 6554
rect 32939 6502 32991 6554
rect 33003 6502 33055 6554
rect 33067 6502 33119 6554
rect 2320 6375 2372 6384
rect 2320 6341 2329 6375
rect 2329 6341 2363 6375
rect 2363 6341 2372 6375
rect 2320 6332 2372 6341
rect 2136 6307 2188 6316
rect 2136 6273 2145 6307
rect 2145 6273 2179 6307
rect 2179 6273 2188 6307
rect 2136 6264 2188 6273
rect 47492 6264 47544 6316
rect 2780 6239 2832 6248
rect 2780 6205 2789 6239
rect 2789 6205 2823 6239
rect 2823 6205 2832 6239
rect 2780 6196 2832 6205
rect 45192 6239 45244 6248
rect 45192 6205 45201 6239
rect 45201 6205 45235 6239
rect 45235 6205 45244 6239
rect 45192 6196 45244 6205
rect 45376 6239 45428 6248
rect 45376 6205 45385 6239
rect 45385 6205 45419 6239
rect 45419 6205 45428 6239
rect 45376 6196 45428 6205
rect 46572 6239 46624 6248
rect 46572 6205 46581 6239
rect 46581 6205 46615 6239
rect 46615 6205 46624 6239
rect 46572 6196 46624 6205
rect 46388 6060 46440 6112
rect 8915 5958 8967 6010
rect 8979 5958 9031 6010
rect 9043 5958 9095 6010
rect 9107 5958 9159 6010
rect 9171 5958 9223 6010
rect 24846 5958 24898 6010
rect 24910 5958 24962 6010
rect 24974 5958 25026 6010
rect 25038 5958 25090 6010
rect 25102 5958 25154 6010
rect 40776 5958 40828 6010
rect 40840 5958 40892 6010
rect 40904 5958 40956 6010
rect 40968 5958 41020 6010
rect 41032 5958 41084 6010
rect 45192 5899 45244 5908
rect 45192 5865 45201 5899
rect 45201 5865 45235 5899
rect 45235 5865 45244 5899
rect 45192 5856 45244 5865
rect 46664 5763 46716 5772
rect 46664 5729 46673 5763
rect 46673 5729 46707 5763
rect 46707 5729 46716 5763
rect 46664 5720 46716 5729
rect 48136 5763 48188 5772
rect 48136 5729 48145 5763
rect 48145 5729 48179 5763
rect 48179 5729 48188 5763
rect 48136 5720 48188 5729
rect 1952 5695 2004 5704
rect 1952 5661 1961 5695
rect 1961 5661 1995 5695
rect 1995 5661 2004 5695
rect 1952 5652 2004 5661
rect 2504 5652 2556 5704
rect 3240 5695 3292 5704
rect 3240 5661 3249 5695
rect 3249 5661 3283 5695
rect 3283 5661 3292 5695
rect 3240 5652 3292 5661
rect 5724 5695 5776 5704
rect 5724 5661 5733 5695
rect 5733 5661 5767 5695
rect 5767 5661 5776 5695
rect 5724 5652 5776 5661
rect 45652 5695 45704 5704
rect 45652 5661 45661 5695
rect 45661 5661 45695 5695
rect 45695 5661 45704 5695
rect 45652 5652 45704 5661
rect 27988 5584 28040 5636
rect 47952 5627 48004 5636
rect 47952 5593 47961 5627
rect 47961 5593 47995 5627
rect 47995 5593 48004 5627
rect 47952 5584 48004 5593
rect 2320 5516 2372 5568
rect 16880 5414 16932 5466
rect 16944 5414 16996 5466
rect 17008 5414 17060 5466
rect 17072 5414 17124 5466
rect 17136 5414 17188 5466
rect 32811 5414 32863 5466
rect 32875 5414 32927 5466
rect 32939 5414 32991 5466
rect 33003 5414 33055 5466
rect 33067 5414 33119 5466
rect 47952 5312 48004 5364
rect 2320 5287 2372 5296
rect 2320 5253 2329 5287
rect 2329 5253 2363 5287
rect 2363 5253 2372 5287
rect 2320 5244 2372 5253
rect 1952 5176 2004 5228
rect 10232 5244 10284 5296
rect 8300 5176 8352 5228
rect 27988 5219 28040 5228
rect 27988 5185 27997 5219
rect 27997 5185 28031 5219
rect 28031 5185 28040 5219
rect 27988 5176 28040 5185
rect 31484 5176 31536 5228
rect 45652 5244 45704 5296
rect 47308 5176 47360 5228
rect 2780 5151 2832 5160
rect 2780 5117 2789 5151
rect 2789 5117 2823 5151
rect 2823 5117 2832 5151
rect 2780 5108 2832 5117
rect 46388 5108 46440 5160
rect 46848 5151 46900 5160
rect 46848 5117 46857 5151
rect 46857 5117 46891 5151
rect 46891 5117 46900 5151
rect 46848 5108 46900 5117
rect 1492 5015 1544 5024
rect 1492 4981 1501 5015
rect 1501 4981 1535 5015
rect 1535 4981 1544 5015
rect 1492 4972 1544 4981
rect 5172 4972 5224 5024
rect 6552 4972 6604 5024
rect 28080 5015 28132 5024
rect 28080 4981 28089 5015
rect 28089 4981 28123 5015
rect 28123 4981 28132 5015
rect 28080 4972 28132 4981
rect 32680 4972 32732 5024
rect 44456 4972 44508 5024
rect 44732 5015 44784 5024
rect 44732 4981 44741 5015
rect 44741 4981 44775 5015
rect 44775 4981 44784 5015
rect 44732 4972 44784 4981
rect 8915 4870 8967 4922
rect 8979 4870 9031 4922
rect 9043 4870 9095 4922
rect 9107 4870 9159 4922
rect 9171 4870 9223 4922
rect 24846 4870 24898 4922
rect 24910 4870 24962 4922
rect 24974 4870 25026 4922
rect 25038 4870 25090 4922
rect 25102 4870 25154 4922
rect 40776 4870 40828 4922
rect 40840 4870 40892 4922
rect 40904 4870 40956 4922
rect 40968 4870 41020 4922
rect 41032 4870 41084 4922
rect 45376 4768 45428 4820
rect 1400 4675 1452 4684
rect 1400 4641 1409 4675
rect 1409 4641 1443 4675
rect 1443 4641 1452 4675
rect 1400 4632 1452 4641
rect 3240 4675 3292 4684
rect 3240 4641 3249 4675
rect 3249 4641 3283 4675
rect 3283 4641 3292 4675
rect 3240 4632 3292 4641
rect 5172 4675 5224 4684
rect 5172 4641 5181 4675
rect 5181 4641 5215 4675
rect 5215 4641 5224 4675
rect 5172 4632 5224 4641
rect 5540 4675 5592 4684
rect 5540 4641 5549 4675
rect 5549 4641 5583 4675
rect 5583 4641 5592 4675
rect 5540 4632 5592 4641
rect 46296 4675 46348 4684
rect 4068 4564 4120 4616
rect 4988 4607 5040 4616
rect 4988 4573 4997 4607
rect 4997 4573 5031 4607
rect 5031 4573 5040 4607
rect 4988 4564 5040 4573
rect 8760 4564 8812 4616
rect 15752 4607 15804 4616
rect 15752 4573 15761 4607
rect 15761 4573 15795 4607
rect 15795 4573 15804 4607
rect 15752 4564 15804 4573
rect 27896 4607 27948 4616
rect 27896 4573 27905 4607
rect 27905 4573 27939 4607
rect 27939 4573 27948 4607
rect 27896 4564 27948 4573
rect 29000 4564 29052 4616
rect 32036 4607 32088 4616
rect 32036 4573 32045 4607
rect 32045 4573 32079 4607
rect 32079 4573 32088 4607
rect 32036 4564 32088 4573
rect 32772 4564 32824 4616
rect 34520 4564 34572 4616
rect 34704 4607 34756 4616
rect 34704 4573 34713 4607
rect 34713 4573 34747 4607
rect 34747 4573 34756 4607
rect 34704 4564 34756 4573
rect 35900 4607 35952 4616
rect 35900 4573 35909 4607
rect 35909 4573 35943 4607
rect 35943 4573 35952 4607
rect 35900 4564 35952 4573
rect 37280 4564 37332 4616
rect 42340 4607 42392 4616
rect 42340 4573 42349 4607
rect 42349 4573 42383 4607
rect 42383 4573 42392 4607
rect 42340 4564 42392 4573
rect 43260 4607 43312 4616
rect 43260 4573 43269 4607
rect 43269 4573 43303 4607
rect 43303 4573 43312 4607
rect 43260 4564 43312 4573
rect 43720 4607 43772 4616
rect 43720 4573 43729 4607
rect 43729 4573 43763 4607
rect 43763 4573 43772 4607
rect 43720 4564 43772 4573
rect 46296 4641 46305 4675
rect 46305 4641 46339 4675
rect 46339 4641 46348 4675
rect 46296 4632 46348 4641
rect 45468 4564 45520 4616
rect 7840 4539 7892 4548
rect 7840 4505 7849 4539
rect 7849 4505 7883 4539
rect 7883 4505 7892 4539
rect 7840 4496 7892 4505
rect 2688 4428 2740 4480
rect 9956 4496 10008 4548
rect 10416 4496 10468 4548
rect 46664 4496 46716 4548
rect 48320 4496 48372 4548
rect 33140 4471 33192 4480
rect 33140 4437 33149 4471
rect 33149 4437 33183 4471
rect 33183 4437 33192 4471
rect 33140 4428 33192 4437
rect 34796 4471 34848 4480
rect 34796 4437 34805 4471
rect 34805 4437 34839 4471
rect 34839 4437 34848 4471
rect 34796 4428 34848 4437
rect 42616 4428 42668 4480
rect 43168 4471 43220 4480
rect 43168 4437 43177 4471
rect 43177 4437 43211 4471
rect 43211 4437 43220 4471
rect 43168 4428 43220 4437
rect 16880 4326 16932 4378
rect 16944 4326 16996 4378
rect 17008 4326 17060 4378
rect 17072 4326 17124 4378
rect 17136 4326 17188 4378
rect 32811 4326 32863 4378
rect 32875 4326 32927 4378
rect 32939 4326 32991 4378
rect 33003 4326 33055 4378
rect 33067 4326 33119 4378
rect 4068 4156 4120 4208
rect 6552 4199 6604 4208
rect 6552 4165 6561 4199
rect 6561 4165 6595 4199
rect 6595 4165 6604 4199
rect 6552 4156 6604 4165
rect 28080 4199 28132 4208
rect 28080 4165 28089 4199
rect 28089 4165 28123 4199
rect 28123 4165 28132 4199
rect 28080 4156 28132 4165
rect 33140 4199 33192 4208
rect 33140 4165 33149 4199
rect 33149 4165 33183 4199
rect 33183 4165 33192 4199
rect 33140 4156 33192 4165
rect 4988 4131 5040 4140
rect 4988 4097 4997 4131
rect 4997 4097 5031 4131
rect 5031 4097 5040 4131
rect 4988 4088 5040 4097
rect 8300 4088 8352 4140
rect 2872 4063 2924 4072
rect 2872 4029 2881 4063
rect 2881 4029 2915 4063
rect 2915 4029 2924 4063
rect 2872 4020 2924 4029
rect 3884 4020 3936 4072
rect 4528 4063 4580 4072
rect 4528 4029 4537 4063
rect 4537 4029 4571 4063
rect 4571 4029 4580 4063
rect 4528 4020 4580 4029
rect 5264 4020 5316 4072
rect 15108 4088 15160 4140
rect 17960 4088 18012 4140
rect 20168 4088 20220 4140
rect 27712 4088 27764 4140
rect 27896 4131 27948 4140
rect 27896 4097 27905 4131
rect 27905 4097 27939 4131
rect 27939 4097 27948 4131
rect 27896 4088 27948 4097
rect 32128 4131 32180 4140
rect 32128 4097 32137 4131
rect 32137 4097 32171 4131
rect 32171 4097 32180 4131
rect 32128 4088 32180 4097
rect 32680 4088 32732 4140
rect 36544 4131 36596 4140
rect 18696 4063 18748 4072
rect 3976 3952 4028 4004
rect 7472 3952 7524 4004
rect 7840 3952 7892 4004
rect 13176 3952 13228 4004
rect 15476 3952 15528 4004
rect 18696 4029 18705 4063
rect 18705 4029 18739 4063
rect 18739 4029 18748 4063
rect 18696 4020 18748 4029
rect 19340 4020 19392 4072
rect 20076 4063 20128 4072
rect 20076 4029 20085 4063
rect 20085 4029 20119 4063
rect 20119 4029 20128 4063
rect 20076 4020 20128 4029
rect 25504 4020 25556 4072
rect 27252 4063 27304 4072
rect 27252 4029 27261 4063
rect 27261 4029 27295 4063
rect 27295 4029 27304 4063
rect 27252 4020 27304 4029
rect 28356 4063 28408 4072
rect 28356 4029 28365 4063
rect 28365 4029 28399 4063
rect 28399 4029 28408 4063
rect 28356 4020 28408 4029
rect 33508 4063 33560 4072
rect 33508 4029 33517 4063
rect 33517 4029 33551 4063
rect 33551 4029 33560 4063
rect 33508 4020 33560 4029
rect 36544 4097 36553 4131
rect 36553 4097 36587 4131
rect 36587 4097 36596 4131
rect 36544 4088 36596 4097
rect 37280 4131 37332 4140
rect 37280 4097 37289 4131
rect 37289 4097 37323 4131
rect 37323 4097 37332 4131
rect 37280 4088 37332 4097
rect 27436 3952 27488 4004
rect 32128 3952 32180 4004
rect 37556 4020 37608 4072
rect 40132 4088 40184 4140
rect 44732 4131 44784 4140
rect 44732 4097 44741 4131
rect 44741 4097 44775 4131
rect 44775 4097 44784 4131
rect 44732 4088 44784 4097
rect 47584 4131 47636 4140
rect 47584 4097 47593 4131
rect 47593 4097 47627 4131
rect 47627 4097 47636 4131
rect 47584 4088 47636 4097
rect 1584 3884 1636 3936
rect 5816 3927 5868 3936
rect 5816 3893 5825 3927
rect 5825 3893 5859 3927
rect 5859 3893 5868 3927
rect 5816 3884 5868 3893
rect 9312 3927 9364 3936
rect 9312 3893 9321 3927
rect 9321 3893 9355 3927
rect 9355 3893 9364 3927
rect 9312 3884 9364 3893
rect 9864 3927 9916 3936
rect 9864 3893 9873 3927
rect 9873 3893 9907 3927
rect 9907 3893 9916 3927
rect 9864 3884 9916 3893
rect 11612 3884 11664 3936
rect 12532 3927 12584 3936
rect 12532 3893 12541 3927
rect 12541 3893 12575 3927
rect 12575 3893 12584 3927
rect 12532 3884 12584 3893
rect 14188 3884 14240 3936
rect 15936 3927 15988 3936
rect 15936 3893 15945 3927
rect 15945 3893 15979 3927
rect 15979 3893 15988 3927
rect 15936 3884 15988 3893
rect 18144 3884 18196 3936
rect 25780 3884 25832 3936
rect 31576 3927 31628 3936
rect 31576 3893 31585 3927
rect 31585 3893 31619 3927
rect 31619 3893 31628 3927
rect 31576 3884 31628 3893
rect 32220 3927 32272 3936
rect 32220 3893 32229 3927
rect 32229 3893 32263 3927
rect 32263 3893 32272 3927
rect 32220 3884 32272 3893
rect 34888 3884 34940 3936
rect 36084 3884 36136 3936
rect 41880 4020 41932 4072
rect 43168 4020 43220 4072
rect 43260 3952 43312 4004
rect 45100 4020 45152 4072
rect 47032 4020 47084 4072
rect 46848 3952 46900 4004
rect 39948 3927 40000 3936
rect 39948 3893 39957 3927
rect 39957 3893 39991 3927
rect 39991 3893 40000 3927
rect 39948 3884 40000 3893
rect 42432 3884 42484 3936
rect 46480 3884 46532 3936
rect 8915 3782 8967 3834
rect 8979 3782 9031 3834
rect 9043 3782 9095 3834
rect 9107 3782 9159 3834
rect 9171 3782 9223 3834
rect 24846 3782 24898 3834
rect 24910 3782 24962 3834
rect 24974 3782 25026 3834
rect 25038 3782 25090 3834
rect 25102 3782 25154 3834
rect 40776 3782 40828 3834
rect 40840 3782 40892 3834
rect 40904 3782 40956 3834
rect 40968 3782 41020 3834
rect 41032 3782 41084 3834
rect 3884 3723 3936 3732
rect 3884 3689 3893 3723
rect 3893 3689 3927 3723
rect 3927 3689 3936 3723
rect 3884 3680 3936 3689
rect 4528 3680 4580 3732
rect 5264 3723 5316 3732
rect 5264 3689 5273 3723
rect 5273 3689 5307 3723
rect 5307 3689 5316 3723
rect 5264 3680 5316 3689
rect 1492 3612 1544 3664
rect 4068 3612 4120 3664
rect 11704 3680 11756 3732
rect 19340 3723 19392 3732
rect 1584 3587 1636 3596
rect 1584 3553 1593 3587
rect 1593 3553 1627 3587
rect 1627 3553 1636 3587
rect 1584 3544 1636 3553
rect 2780 3587 2832 3596
rect 2780 3553 2789 3587
rect 2789 3553 2823 3587
rect 2823 3553 2832 3587
rect 2780 3544 2832 3553
rect 5724 3587 5776 3596
rect 5724 3553 5733 3587
rect 5733 3553 5767 3587
rect 5767 3553 5776 3587
rect 5724 3544 5776 3553
rect 5908 3544 5960 3596
rect 9864 3612 9916 3664
rect 9956 3612 10008 3664
rect 9312 3587 9364 3596
rect 9312 3553 9321 3587
rect 9321 3553 9355 3587
rect 9355 3553 9364 3587
rect 9312 3544 9364 3553
rect 9680 3587 9732 3596
rect 9680 3553 9689 3587
rect 9689 3553 9723 3587
rect 9723 3553 9732 3587
rect 9680 3544 9732 3553
rect 11612 3587 11664 3596
rect 11612 3553 11621 3587
rect 11621 3553 11655 3587
rect 11655 3553 11664 3587
rect 11612 3544 11664 3553
rect 12256 3587 12308 3596
rect 12256 3553 12265 3587
rect 12265 3553 12299 3587
rect 12299 3553 12308 3587
rect 12256 3544 12308 3553
rect 8208 3519 8260 3528
rect 8208 3485 8217 3519
rect 8217 3485 8251 3519
rect 8251 3485 8260 3519
rect 8208 3476 8260 3485
rect 13176 3612 13228 3664
rect 19340 3689 19349 3723
rect 19349 3689 19383 3723
rect 19383 3689 19392 3723
rect 19340 3680 19392 3689
rect 20076 3723 20128 3732
rect 20076 3689 20085 3723
rect 20085 3689 20119 3723
rect 20119 3689 20128 3723
rect 20076 3680 20128 3689
rect 15752 3587 15804 3596
rect 15752 3553 15761 3587
rect 15761 3553 15795 3587
rect 15795 3553 15804 3587
rect 15752 3544 15804 3553
rect 15936 3587 15988 3596
rect 15936 3553 15945 3587
rect 15945 3553 15979 3587
rect 15979 3553 15988 3587
rect 15936 3544 15988 3553
rect 16120 3544 16172 3596
rect 19432 3612 19484 3664
rect 19708 3612 19760 3664
rect 32128 3680 32180 3732
rect 45100 3723 45152 3732
rect 45100 3689 45109 3723
rect 45109 3689 45143 3723
rect 45143 3689 45152 3723
rect 45100 3680 45152 3689
rect 26976 3612 27028 3664
rect 27712 3587 27764 3596
rect 15108 3519 15160 3528
rect 5724 3408 5776 3460
rect 11796 3451 11848 3460
rect 11796 3417 11805 3451
rect 11805 3417 11839 3451
rect 11839 3417 11848 3451
rect 11796 3408 11848 3417
rect 15108 3485 15117 3519
rect 15117 3485 15151 3519
rect 15151 3485 15160 3519
rect 15108 3476 15160 3485
rect 19156 3476 19208 3528
rect 20168 3476 20220 3528
rect 23940 3476 23992 3528
rect 27712 3553 27721 3587
rect 27721 3553 27755 3587
rect 27755 3553 27764 3587
rect 27712 3544 27764 3553
rect 32036 3587 32088 3596
rect 32036 3553 32045 3587
rect 32045 3553 32079 3587
rect 32079 3553 32088 3587
rect 32036 3544 32088 3553
rect 32220 3587 32272 3596
rect 32220 3553 32229 3587
rect 32229 3553 32263 3587
rect 32263 3553 32272 3587
rect 32220 3544 32272 3553
rect 32680 3587 32732 3596
rect 32680 3553 32689 3587
rect 32689 3553 32723 3587
rect 32723 3553 32732 3587
rect 32680 3544 32732 3553
rect 35900 3587 35952 3596
rect 35900 3553 35909 3587
rect 35909 3553 35943 3587
rect 35943 3553 35952 3587
rect 36084 3587 36136 3596
rect 35900 3544 35952 3553
rect 36084 3553 36093 3587
rect 36093 3553 36127 3587
rect 36127 3553 36136 3587
rect 36084 3544 36136 3553
rect 36728 3587 36780 3596
rect 36728 3553 36737 3587
rect 36737 3553 36771 3587
rect 36771 3553 36780 3587
rect 36728 3544 36780 3553
rect 43812 3544 43864 3596
rect 25504 3519 25556 3528
rect 25504 3485 25513 3519
rect 25513 3485 25547 3519
rect 25547 3485 25556 3519
rect 25504 3476 25556 3485
rect 28816 3476 28868 3528
rect 31944 3476 31996 3528
rect 34704 3519 34756 3528
rect 34704 3485 34713 3519
rect 34713 3485 34747 3519
rect 34747 3485 34756 3519
rect 34704 3476 34756 3485
rect 37280 3476 37332 3528
rect 39120 3519 39172 3528
rect 39120 3485 39129 3519
rect 39129 3485 39163 3519
rect 39163 3485 39172 3519
rect 39120 3476 39172 3485
rect 39856 3519 39908 3528
rect 39856 3485 39865 3519
rect 39865 3485 39899 3519
rect 39899 3485 39908 3519
rect 39856 3476 39908 3485
rect 42432 3519 42484 3528
rect 42432 3485 42441 3519
rect 42441 3485 42475 3519
rect 42475 3485 42484 3519
rect 42432 3476 42484 3485
rect 47584 3612 47636 3664
rect 46480 3587 46532 3596
rect 46480 3553 46489 3587
rect 46489 3553 46523 3587
rect 46523 3553 46532 3587
rect 46480 3544 46532 3553
rect 20444 3408 20496 3460
rect 27068 3451 27120 3460
rect 27068 3417 27077 3451
rect 27077 3417 27111 3451
rect 27111 3417 27120 3451
rect 27068 3408 27120 3417
rect 27252 3408 27304 3460
rect 35164 3408 35216 3460
rect 41696 3451 41748 3460
rect 41696 3417 41714 3451
rect 41714 3417 41748 3451
rect 42616 3451 42668 3460
rect 41696 3408 41748 3417
rect 42616 3417 42625 3451
rect 42625 3417 42659 3451
rect 42659 3417 42668 3451
rect 42616 3408 42668 3417
rect 45100 3408 45152 3460
rect 48136 3451 48188 3460
rect 48136 3417 48145 3451
rect 48145 3417 48179 3451
rect 48179 3417 48188 3451
rect 48136 3408 48188 3417
rect 8116 3340 8168 3392
rect 8300 3383 8352 3392
rect 8300 3349 8309 3383
rect 8309 3349 8343 3383
rect 8343 3349 8352 3383
rect 8300 3340 8352 3349
rect 14372 3383 14424 3392
rect 14372 3349 14381 3383
rect 14381 3349 14415 3383
rect 14415 3349 14424 3383
rect 14372 3340 14424 3349
rect 15292 3340 15344 3392
rect 18328 3340 18380 3392
rect 24124 3340 24176 3392
rect 26240 3340 26292 3392
rect 35072 3340 35124 3392
rect 40132 3340 40184 3392
rect 41880 3340 41932 3392
rect 16880 3238 16932 3290
rect 16944 3238 16996 3290
rect 17008 3238 17060 3290
rect 17072 3238 17124 3290
rect 17136 3238 17188 3290
rect 32811 3238 32863 3290
rect 32875 3238 32927 3290
rect 32939 3238 32991 3290
rect 33003 3238 33055 3290
rect 33067 3238 33119 3290
rect 5724 3179 5776 3188
rect 5724 3145 5733 3179
rect 5733 3145 5767 3179
rect 5767 3145 5776 3179
rect 5724 3136 5776 3145
rect 8116 3136 8168 3188
rect 11796 3179 11848 3188
rect 4620 3043 4672 3052
rect 4620 3009 4629 3043
rect 4629 3009 4663 3043
rect 4663 3009 4672 3043
rect 4620 3000 4672 3009
rect 11796 3145 11805 3179
rect 11805 3145 11839 3179
rect 11839 3145 11848 3179
rect 11796 3136 11848 3145
rect 15292 3111 15344 3120
rect 15292 3077 15301 3111
rect 15301 3077 15335 3111
rect 15335 3077 15344 3111
rect 15292 3068 15344 3077
rect 18052 3136 18104 3188
rect 27068 3179 27120 3188
rect 18144 3068 18196 3120
rect 18328 3111 18380 3120
rect 18328 3077 18337 3111
rect 18337 3077 18371 3111
rect 18371 3077 18380 3111
rect 18328 3068 18380 3077
rect 19340 3068 19392 3120
rect 24124 3111 24176 3120
rect 2320 2975 2372 2984
rect 2320 2941 2329 2975
rect 2329 2941 2363 2975
rect 2363 2941 2372 2975
rect 2320 2932 2372 2941
rect 2596 2975 2648 2984
rect 2596 2941 2605 2975
rect 2605 2941 2639 2975
rect 2639 2941 2648 2975
rect 2596 2932 2648 2941
rect 3884 2932 3936 2984
rect 5540 2932 5592 2984
rect 7472 2932 7524 2984
rect 4620 2864 4672 2916
rect 6736 2864 6788 2916
rect 11704 3043 11756 3052
rect 11704 3009 11713 3043
rect 11713 3009 11747 3043
rect 11747 3009 11756 3043
rect 11704 3000 11756 3009
rect 9312 2975 9364 2984
rect 9312 2941 9321 2975
rect 9321 2941 9355 2975
rect 9355 2941 9364 2975
rect 9312 2932 9364 2941
rect 13820 2975 13872 2984
rect 13820 2941 13829 2975
rect 13829 2941 13863 2975
rect 13863 2941 13872 2975
rect 13820 2932 13872 2941
rect 15476 3043 15528 3052
rect 15476 3009 15485 3043
rect 15485 3009 15519 3043
rect 15519 3009 15528 3043
rect 15476 3000 15528 3009
rect 20444 3043 20496 3052
rect 15568 2932 15620 2984
rect 12440 2864 12492 2916
rect 20444 3009 20453 3043
rect 20453 3009 20487 3043
rect 20487 3009 20496 3043
rect 20444 3000 20496 3009
rect 24124 3077 24133 3111
rect 24133 3077 24167 3111
rect 24167 3077 24176 3111
rect 24124 3068 24176 3077
rect 27068 3145 27077 3179
rect 27077 3145 27111 3179
rect 27111 3145 27120 3179
rect 27068 3136 27120 3145
rect 23756 3000 23808 3052
rect 23940 3043 23992 3052
rect 23940 3009 23949 3043
rect 23949 3009 23983 3043
rect 23983 3009 23992 3043
rect 23940 3000 23992 3009
rect 26976 3043 27028 3052
rect 26976 3009 26985 3043
rect 26985 3009 27019 3043
rect 27019 3009 27028 3043
rect 26976 3000 27028 3009
rect 28816 3043 28868 3052
rect 19340 2975 19392 2984
rect 19340 2941 19349 2975
rect 19349 2941 19383 2975
rect 19383 2941 19392 2975
rect 19340 2932 19392 2941
rect 28816 3009 28825 3043
rect 28825 3009 28859 3043
rect 28859 3009 28868 3043
rect 28816 3000 28868 3009
rect 29092 2932 29144 2984
rect 29644 2975 29696 2984
rect 29644 2941 29653 2975
rect 29653 2941 29687 2975
rect 29687 2941 29696 2975
rect 29644 2932 29696 2941
rect 23664 2864 23716 2916
rect 23756 2864 23808 2916
rect 39856 3136 39908 3188
rect 41696 3179 41748 3188
rect 41696 3145 41705 3179
rect 41705 3145 41739 3179
rect 41739 3145 41748 3179
rect 41696 3136 41748 3145
rect 46664 3179 46716 3188
rect 35072 3111 35124 3120
rect 35072 3077 35081 3111
rect 35081 3077 35115 3111
rect 35115 3077 35124 3111
rect 35072 3068 35124 3077
rect 35164 3068 35216 3120
rect 31392 3043 31444 3052
rect 31392 3009 31401 3043
rect 31401 3009 31435 3043
rect 31435 3009 31444 3043
rect 31392 3000 31444 3009
rect 31576 3000 31628 3052
rect 34888 3043 34940 3052
rect 34888 3009 34897 3043
rect 34897 3009 34931 3043
rect 34931 3009 34940 3043
rect 34888 3000 34940 3009
rect 37372 3000 37424 3052
rect 39120 3043 39172 3052
rect 39120 3009 39129 3043
rect 39129 3009 39163 3043
rect 39163 3009 39172 3043
rect 39120 3000 39172 3009
rect 41880 3043 41932 3052
rect 41880 3009 41889 3043
rect 41889 3009 41923 3043
rect 41923 3009 41932 3043
rect 41880 3000 41932 3009
rect 46664 3145 46673 3179
rect 46673 3145 46707 3179
rect 46707 3145 46716 3179
rect 46664 3136 46716 3145
rect 45468 3043 45520 3052
rect 45468 3009 45477 3043
rect 45477 3009 45511 3043
rect 45511 3009 45520 3043
rect 45468 3000 45520 3009
rect 46756 3043 46808 3052
rect 46756 3009 46765 3043
rect 46765 3009 46799 3043
rect 46799 3009 46808 3043
rect 46756 3000 46808 3009
rect 47400 3000 47452 3052
rect 33968 2975 34020 2984
rect 33968 2941 33977 2975
rect 33977 2941 34011 2975
rect 34011 2941 34020 2975
rect 33968 2932 34020 2941
rect 36084 2975 36136 2984
rect 36084 2941 36093 2975
rect 36093 2941 36127 2975
rect 36127 2941 36136 2975
rect 36084 2932 36136 2941
rect 43720 2932 43772 2984
rect 43904 2975 43956 2984
rect 43904 2941 43913 2975
rect 43913 2941 43947 2975
rect 43947 2941 43956 2975
rect 43904 2932 43956 2941
rect 44364 2864 44416 2916
rect 46572 2864 46624 2916
rect 49608 2864 49660 2916
rect 4528 2839 4580 2848
rect 4528 2805 4537 2839
rect 4537 2805 4571 2839
rect 4571 2805 4580 2839
rect 4528 2796 4580 2805
rect 6552 2796 6604 2848
rect 13360 2796 13412 2848
rect 16028 2839 16080 2848
rect 16028 2805 16037 2839
rect 16037 2805 16071 2839
rect 16071 2805 16080 2839
rect 16028 2796 16080 2805
rect 16672 2839 16724 2848
rect 16672 2805 16681 2839
rect 16681 2805 16715 2839
rect 16715 2805 16724 2839
rect 16672 2796 16724 2805
rect 21088 2796 21140 2848
rect 21272 2839 21324 2848
rect 21272 2805 21281 2839
rect 21281 2805 21315 2839
rect 21315 2805 21324 2839
rect 21272 2796 21324 2805
rect 23848 2796 23900 2848
rect 26424 2839 26476 2848
rect 26424 2805 26433 2839
rect 26433 2805 26467 2839
rect 26467 2805 26476 2839
rect 26424 2796 26476 2805
rect 37464 2796 37516 2848
rect 45560 2839 45612 2848
rect 45560 2805 45569 2839
rect 45569 2805 45603 2839
rect 45603 2805 45612 2839
rect 47676 2839 47728 2848
rect 45560 2796 45612 2805
rect 47676 2805 47685 2839
rect 47685 2805 47719 2839
rect 47719 2805 47728 2839
rect 47676 2796 47728 2805
rect 8915 2694 8967 2746
rect 8979 2694 9031 2746
rect 9043 2694 9095 2746
rect 9107 2694 9159 2746
rect 9171 2694 9223 2746
rect 24846 2694 24898 2746
rect 24910 2694 24962 2746
rect 24974 2694 25026 2746
rect 25038 2694 25090 2746
rect 25102 2694 25154 2746
rect 40776 2694 40828 2746
rect 40840 2694 40892 2746
rect 40904 2694 40956 2746
rect 40968 2694 41020 2746
rect 41032 2694 41084 2746
rect 2320 2592 2372 2644
rect 5540 2592 5592 2644
rect 3240 2524 3292 2576
rect 4528 2456 4580 2508
rect 7748 2524 7800 2576
rect 5816 2456 5868 2508
rect 6552 2499 6604 2508
rect 6552 2465 6561 2499
rect 6561 2465 6595 2499
rect 6595 2465 6604 2499
rect 6552 2456 6604 2465
rect 6736 2456 6788 2508
rect 8760 2456 8812 2508
rect 12532 2524 12584 2576
rect 13360 2499 13412 2508
rect 13360 2465 13369 2499
rect 13369 2465 13403 2499
rect 13403 2465 13412 2499
rect 13360 2456 13412 2465
rect 2688 2388 2740 2440
rect 3516 2320 3568 2372
rect 8208 2320 8260 2372
rect 8300 2320 8352 2372
rect 3424 2252 3476 2304
rect 14188 2499 14240 2508
rect 14188 2465 14197 2499
rect 14197 2465 14231 2499
rect 14231 2465 14240 2499
rect 14188 2456 14240 2465
rect 14372 2499 14424 2508
rect 14372 2465 14381 2499
rect 14381 2465 14415 2499
rect 14415 2465 14424 2499
rect 14372 2456 14424 2465
rect 14832 2499 14884 2508
rect 14832 2465 14841 2499
rect 14841 2465 14875 2499
rect 14875 2465 14884 2499
rect 14832 2456 14884 2465
rect 16672 2499 16724 2508
rect 16672 2465 16681 2499
rect 16681 2465 16715 2499
rect 16715 2465 16724 2499
rect 16672 2456 16724 2465
rect 25872 2524 25924 2576
rect 37372 2592 37424 2644
rect 20812 2499 20864 2508
rect 20812 2465 20821 2499
rect 20821 2465 20855 2499
rect 20855 2465 20864 2499
rect 20812 2456 20864 2465
rect 21088 2499 21140 2508
rect 21088 2465 21097 2499
rect 21097 2465 21131 2499
rect 21131 2465 21140 2499
rect 21088 2456 21140 2465
rect 21272 2499 21324 2508
rect 21272 2465 21281 2499
rect 21281 2465 21315 2499
rect 21315 2465 21324 2499
rect 21272 2456 21324 2465
rect 22468 2499 22520 2508
rect 22468 2465 22477 2499
rect 22477 2465 22511 2499
rect 22511 2465 22520 2499
rect 22468 2456 22520 2465
rect 23664 2499 23716 2508
rect 23664 2465 23673 2499
rect 23673 2465 23707 2499
rect 23707 2465 23716 2499
rect 23664 2456 23716 2465
rect 23848 2499 23900 2508
rect 23848 2465 23857 2499
rect 23857 2465 23891 2499
rect 23891 2465 23900 2499
rect 23848 2456 23900 2465
rect 26240 2499 26292 2508
rect 26240 2465 26249 2499
rect 26249 2465 26283 2499
rect 26283 2465 26292 2499
rect 26424 2499 26476 2508
rect 26240 2456 26292 2465
rect 26424 2465 26433 2499
rect 26433 2465 26467 2499
rect 26467 2465 26476 2499
rect 26424 2456 26476 2465
rect 28816 2456 28868 2508
rect 29000 2499 29052 2508
rect 29000 2465 29009 2499
rect 29009 2465 29043 2499
rect 29043 2465 29052 2499
rect 29000 2456 29052 2465
rect 29092 2388 29144 2440
rect 31576 2524 31628 2576
rect 31944 2456 31996 2508
rect 34796 2524 34848 2576
rect 34520 2456 34572 2508
rect 37280 2499 37332 2508
rect 37280 2465 37289 2499
rect 37289 2465 37323 2499
rect 37323 2465 37332 2499
rect 37280 2456 37332 2465
rect 37464 2499 37516 2508
rect 37464 2465 37473 2499
rect 37473 2465 37507 2499
rect 37507 2465 37516 2499
rect 37464 2456 37516 2465
rect 39948 2499 40000 2508
rect 39948 2465 39957 2499
rect 39957 2465 39991 2499
rect 39991 2465 40000 2499
rect 39948 2456 40000 2465
rect 40132 2499 40184 2508
rect 40132 2465 40141 2499
rect 40141 2465 40175 2499
rect 40175 2465 40184 2499
rect 40132 2456 40184 2465
rect 45744 2524 45796 2576
rect 43812 2456 43864 2508
rect 46572 2499 46624 2508
rect 44456 2431 44508 2440
rect 44456 2397 44465 2431
rect 44465 2397 44499 2431
rect 44499 2397 44508 2431
rect 46572 2465 46581 2499
rect 46581 2465 46615 2499
rect 46615 2465 46624 2499
rect 46572 2456 46624 2465
rect 47676 2456 47728 2508
rect 44456 2388 44508 2397
rect 45652 2388 45704 2440
rect 16028 2320 16080 2372
rect 24584 2363 24636 2372
rect 24584 2329 24593 2363
rect 24593 2329 24627 2363
rect 24627 2329 24636 2363
rect 24584 2320 24636 2329
rect 39304 2320 39356 2372
rect 44180 2320 44232 2372
rect 45560 2320 45612 2372
rect 47676 2252 47728 2304
rect 16880 2150 16932 2202
rect 16944 2150 16996 2202
rect 17008 2150 17060 2202
rect 17072 2150 17124 2202
rect 17136 2150 17188 2202
rect 32811 2150 32863 2202
rect 32875 2150 32927 2202
rect 32939 2150 32991 2202
rect 33003 2150 33055 2202
rect 33067 2150 33119 2202
rect 8208 2048 8260 2100
rect 13820 2048 13872 2100
rect 664 1980 716 2032
rect 24584 1980 24636 2032
rect 20812 1912 20864 1964
rect 32220 1912 32272 1964
rect 33968 1300 34020 1352
rect 46664 1300 46716 1352
rect 44180 1028 44232 1080
rect 46848 1028 46900 1080
<< metal2 >>
rect -10 19200 102 20000
rect 634 19200 746 20000
rect 1278 19200 1390 20000
rect 1922 19200 2034 20000
rect 2566 19200 2678 20000
rect 3210 19200 3322 20000
rect 3854 19200 3966 20000
rect 4498 19200 4610 20000
rect 5142 19200 5254 20000
rect 5786 19200 5898 20000
rect 6430 19200 6542 20000
rect 7074 19200 7186 20000
rect 7718 19200 7830 20000
rect 8362 19200 8474 20000
rect 9006 19200 9118 20000
rect 9650 19200 9762 20000
rect 10294 19200 10406 20000
rect 10938 19200 11050 20000
rect 11582 19200 11694 20000
rect 12226 19200 12338 20000
rect 12870 19200 12982 20000
rect 13514 19200 13626 20000
rect 14158 19200 14270 20000
rect 14802 19200 14914 20000
rect 16090 19200 16202 20000
rect 16734 19200 16846 20000
rect 17378 19200 17490 20000
rect 18022 19200 18134 20000
rect 18666 19200 18778 20000
rect 19310 19200 19422 20000
rect 19954 19200 20066 20000
rect 20598 19200 20710 20000
rect 21242 19200 21354 20000
rect 21886 19200 21998 20000
rect 22530 19200 22642 20000
rect 23174 19200 23286 20000
rect 23818 19200 23930 20000
rect 24462 19200 24574 20000
rect 25106 19200 25218 20000
rect 25750 19200 25862 20000
rect 26394 19200 26506 20000
rect 27038 19200 27150 20000
rect 27682 19200 27794 20000
rect 28326 19200 28438 20000
rect 28970 19200 29082 20000
rect 29614 19200 29726 20000
rect 30258 19200 30370 20000
rect 30902 19200 31014 20000
rect 31546 19200 31658 20000
rect 32190 19200 32302 20000
rect 32834 19200 32946 20000
rect 33478 19200 33590 20000
rect 34122 19200 34234 20000
rect 34766 19200 34878 20000
rect 35410 19200 35522 20000
rect 36054 19200 36166 20000
rect 36698 19200 36810 20000
rect 37342 19200 37454 20000
rect 37986 19200 38098 20000
rect 38630 19200 38742 20000
rect 39274 19200 39386 20000
rect 39918 19200 40030 20000
rect 40562 19200 40674 20000
rect 41206 19200 41318 20000
rect 41850 19200 41962 20000
rect 42494 19200 42606 20000
rect 43138 19200 43250 20000
rect 43782 19200 43894 20000
rect 44426 19200 44538 20000
rect 45070 19200 45182 20000
rect 45714 19200 45826 20000
rect 46358 19200 46470 20000
rect 47002 19200 47114 20000
rect 47646 19200 47758 20000
rect 48290 19200 48402 20000
rect 48934 19200 49046 20000
rect 49578 19200 49690 20000
rect 1398 17776 1454 17785
rect 1398 17711 1454 17720
rect 1412 17270 1440 17711
rect 2608 17270 2636 19200
rect 4620 17536 4672 17542
rect 4620 17478 4672 17484
rect 4068 17332 4120 17338
rect 4068 17274 4120 17280
rect 1400 17264 1452 17270
rect 1400 17206 1452 17212
rect 2596 17264 2648 17270
rect 2596 17206 2648 17212
rect 3056 17128 3108 17134
rect 3056 17070 3108 17076
rect 3240 17128 3292 17134
rect 4080 17105 4108 17274
rect 3240 17070 3292 17076
rect 4066 17096 4122 17105
rect 2412 16584 2464 16590
rect 2412 16526 2464 16532
rect 2044 15904 2096 15910
rect 2044 15846 2096 15852
rect 2056 15026 2084 15846
rect 2424 15502 2452 16526
rect 3068 16522 3096 17070
rect 3252 16794 3280 17070
rect 4066 17031 4122 17040
rect 3240 16788 3292 16794
rect 3240 16730 3292 16736
rect 4632 16658 4660 17478
rect 7760 17134 7788 19200
rect 8300 17264 8352 17270
rect 8300 17206 8352 17212
rect 5632 17128 5684 17134
rect 5632 17070 5684 17076
rect 5816 17128 5868 17134
rect 5816 17070 5868 17076
rect 6552 17128 6604 17134
rect 6552 17070 6604 17076
rect 7564 17128 7616 17134
rect 7564 17070 7616 17076
rect 7748 17128 7800 17134
rect 7748 17070 7800 17076
rect 7932 17128 7984 17134
rect 7932 17070 7984 17076
rect 4620 16652 4672 16658
rect 4620 16594 4672 16600
rect 3056 16516 3108 16522
rect 3056 16458 3108 16464
rect 2778 15736 2834 15745
rect 2778 15671 2834 15680
rect 2412 15496 2464 15502
rect 2412 15438 2464 15444
rect 2228 15360 2280 15366
rect 2228 15302 2280 15308
rect 2240 15094 2268 15302
rect 2228 15088 2280 15094
rect 2228 15030 2280 15036
rect 2044 15020 2096 15026
rect 2044 14962 2096 14968
rect 2044 14408 2096 14414
rect 2044 14350 2096 14356
rect 2056 13938 2084 14350
rect 2228 14272 2280 14278
rect 2228 14214 2280 14220
rect 2240 14006 2268 14214
rect 2228 14000 2280 14006
rect 2228 13942 2280 13948
rect 2044 13932 2096 13938
rect 2044 13874 2096 13880
rect 2044 13320 2096 13326
rect 2044 13262 2096 13268
rect 2056 12850 2084 13262
rect 2044 12844 2096 12850
rect 2044 12786 2096 12792
rect 2228 12776 2280 12782
rect 2228 12718 2280 12724
rect 2240 12442 2268 12718
rect 2228 12436 2280 12442
rect 2228 12378 2280 12384
rect 2044 11144 2096 11150
rect 2044 11086 2096 11092
rect 2056 10674 2084 11086
rect 2044 10668 2096 10674
rect 2044 10610 2096 10616
rect 2044 8968 2096 8974
rect 2044 8910 2096 8916
rect 2056 8498 2084 8910
rect 2044 8492 2096 8498
rect 2044 8434 2096 8440
rect 2228 8424 2280 8430
rect 2228 8366 2280 8372
rect 2240 8090 2268 8366
rect 2228 8084 2280 8090
rect 2228 8026 2280 8032
rect 2424 7886 2452 15438
rect 2792 14958 2820 15671
rect 2780 14952 2832 14958
rect 2780 14894 2832 14900
rect 2688 14408 2740 14414
rect 2688 14350 2740 14356
rect 2778 14376 2834 14385
rect 2596 12232 2648 12238
rect 2596 12174 2648 12180
rect 2504 10600 2556 10606
rect 2504 10542 2556 10548
rect 2516 10266 2544 10542
rect 2504 10260 2556 10266
rect 2504 10202 2556 10208
rect 2412 7880 2464 7886
rect 2412 7822 2464 7828
rect 2136 7200 2188 7206
rect 2136 7142 2188 7148
rect 2148 6322 2176 7142
rect 2608 6914 2636 12174
rect 2700 10062 2728 14350
rect 2778 14311 2834 14320
rect 2792 13870 2820 14311
rect 2780 13864 2832 13870
rect 2780 13806 2832 13812
rect 3792 13320 3844 13326
rect 3792 13262 3844 13268
rect 2778 13016 2834 13025
rect 2778 12951 2834 12960
rect 2792 12782 2820 12951
rect 2780 12776 2832 12782
rect 2780 12718 2832 12724
rect 3804 12306 3832 13262
rect 4066 12336 4122 12345
rect 3792 12300 3844 12306
rect 4066 12271 4068 12280
rect 3792 12242 3844 12248
rect 4120 12271 4122 12280
rect 4068 12242 4120 12248
rect 3976 12164 4028 12170
rect 3976 12106 4028 12112
rect 3988 11898 4016 12106
rect 3976 11892 4028 11898
rect 3976 11834 4028 11840
rect 2778 10976 2834 10985
rect 2778 10911 2834 10920
rect 2792 10606 2820 10911
rect 2780 10600 2832 10606
rect 2780 10542 2832 10548
rect 3422 10296 3478 10305
rect 3422 10231 3478 10240
rect 2688 10056 2740 10062
rect 2688 9998 2740 10004
rect 3436 9994 3464 10231
rect 3424 9988 3476 9994
rect 3424 9930 3476 9936
rect 2780 8424 2832 8430
rect 2780 8366 2832 8372
rect 2792 8265 2820 8366
rect 2778 8256 2834 8265
rect 2778 8191 2834 8200
rect 3422 7576 3478 7585
rect 3422 7511 3478 7520
rect 3436 7274 3464 7511
rect 3424 7268 3476 7274
rect 3424 7210 3476 7216
rect 2516 6886 2636 6914
rect 2778 6896 2834 6905
rect 2320 6656 2372 6662
rect 2320 6598 2372 6604
rect 2332 6390 2360 6598
rect 2320 6384 2372 6390
rect 2320 6326 2372 6332
rect 2136 6316 2188 6322
rect 2136 6258 2188 6264
rect 2516 5710 2544 6886
rect 2778 6831 2834 6840
rect 2688 6792 2740 6798
rect 2688 6734 2740 6740
rect 1952 5704 2004 5710
rect 1952 5646 2004 5652
rect 2504 5704 2556 5710
rect 2504 5646 2556 5652
rect 1964 5234 1992 5646
rect 2320 5568 2372 5574
rect 2320 5510 2372 5516
rect 2332 5302 2360 5510
rect 2320 5296 2372 5302
rect 2320 5238 2372 5244
rect 1952 5228 2004 5234
rect 1952 5170 2004 5176
rect 1492 5024 1544 5030
rect 1492 4966 1544 4972
rect 1398 4856 1454 4865
rect 1398 4791 1454 4800
rect 1412 4690 1440 4791
rect 1400 4684 1452 4690
rect 1400 4626 1452 4632
rect 1504 3670 1532 4966
rect 2700 4486 2728 6734
rect 2792 6254 2820 6831
rect 2780 6248 2832 6254
rect 2780 6190 2832 6196
rect 3240 5704 3292 5710
rect 3240 5646 3292 5652
rect 2778 5536 2834 5545
rect 2778 5471 2834 5480
rect 2792 5166 2820 5471
rect 2780 5160 2832 5166
rect 2780 5102 2832 5108
rect 3252 4690 3280 5646
rect 3240 4684 3292 4690
rect 3240 4626 3292 4632
rect 4068 4616 4120 4622
rect 4068 4558 4120 4564
rect 2688 4480 2740 4486
rect 2688 4422 2740 4428
rect 1584 3936 1636 3942
rect 1584 3878 1636 3884
rect 1492 3664 1544 3670
rect 1492 3606 1544 3612
rect 1596 3602 1624 3878
rect 1584 3596 1636 3602
rect 1584 3538 1636 3544
rect 2320 2984 2372 2990
rect 2320 2926 2372 2932
rect 2596 2984 2648 2990
rect 2596 2926 2648 2932
rect 2332 2650 2360 2926
rect 2320 2644 2372 2650
rect 2320 2586 2372 2592
rect 664 2032 716 2038
rect 664 1974 716 1980
rect 676 800 704 1974
rect 2608 800 2636 2926
rect 2700 2446 2728 4422
rect 4080 4214 4108 4558
rect 4068 4208 4120 4214
rect 2778 4176 2834 4185
rect 4068 4150 4120 4156
rect 2778 4111 2834 4120
rect 2792 3602 2820 4111
rect 2872 4072 2924 4078
rect 2872 4014 2924 4020
rect 3884 4072 3936 4078
rect 3884 4014 3936 4020
rect 2780 3596 2832 3602
rect 2780 3538 2832 3544
rect 2884 2825 2912 4014
rect 3896 3738 3924 4014
rect 3976 4004 4028 4010
rect 3976 3946 4028 3952
rect 3884 3732 3936 3738
rect 3884 3674 3936 3680
rect 3988 3505 4016 3946
rect 4080 3670 4108 4150
rect 4528 4072 4580 4078
rect 4528 4014 4580 4020
rect 4540 3738 4568 4014
rect 4528 3732 4580 3738
rect 4528 3674 4580 3680
rect 4068 3664 4120 3670
rect 4068 3606 4120 3612
rect 3974 3496 4030 3505
rect 3974 3431 4030 3440
rect 4632 3058 4660 16594
rect 5644 16522 5672 17070
rect 5828 16794 5856 17070
rect 6564 16794 6592 17070
rect 5816 16788 5868 16794
rect 5816 16730 5868 16736
rect 6552 16788 6604 16794
rect 6552 16730 6604 16736
rect 5632 16516 5684 16522
rect 5632 16458 5684 16464
rect 7576 16250 7604 17070
rect 7748 16992 7800 16998
rect 7748 16934 7800 16940
rect 7760 16658 7788 16934
rect 7944 16794 7972 17070
rect 7932 16788 7984 16794
rect 7932 16730 7984 16736
rect 7748 16652 7800 16658
rect 7748 16594 7800 16600
rect 7564 16244 7616 16250
rect 7564 16186 7616 16192
rect 7760 14414 7788 16594
rect 8312 16590 8340 17206
rect 8404 17066 8432 19200
rect 8392 17060 8444 17066
rect 8392 17002 8444 17008
rect 8915 16892 9223 16912
rect 8915 16890 8921 16892
rect 8977 16890 9001 16892
rect 9057 16890 9081 16892
rect 9137 16890 9161 16892
rect 9217 16890 9223 16892
rect 8977 16838 8979 16890
rect 9159 16838 9161 16890
rect 8915 16836 8921 16838
rect 8977 16836 9001 16838
rect 9057 16836 9081 16838
rect 9137 16836 9161 16838
rect 9217 16836 9223 16838
rect 8915 16816 9223 16836
rect 8300 16584 8352 16590
rect 8300 16526 8352 16532
rect 9692 16454 9720 19200
rect 10600 16652 10652 16658
rect 10600 16594 10652 16600
rect 10324 16516 10376 16522
rect 10324 16458 10376 16464
rect 9680 16448 9732 16454
rect 9680 16390 9732 16396
rect 10336 16250 10364 16458
rect 10612 16454 10640 16594
rect 10600 16448 10652 16454
rect 10600 16390 10652 16396
rect 10324 16244 10376 16250
rect 10324 16186 10376 16192
rect 10232 16108 10284 16114
rect 10232 16050 10284 16056
rect 8915 15804 9223 15824
rect 8915 15802 8921 15804
rect 8977 15802 9001 15804
rect 9057 15802 9081 15804
rect 9137 15802 9161 15804
rect 9217 15802 9223 15804
rect 8977 15750 8979 15802
rect 9159 15750 9161 15802
rect 8915 15748 8921 15750
rect 8977 15748 9001 15750
rect 9057 15748 9081 15750
rect 9137 15748 9161 15750
rect 9217 15748 9223 15750
rect 8915 15728 9223 15748
rect 8915 14716 9223 14736
rect 8915 14714 8921 14716
rect 8977 14714 9001 14716
rect 9057 14714 9081 14716
rect 9137 14714 9161 14716
rect 9217 14714 9223 14716
rect 8977 14662 8979 14714
rect 9159 14662 9161 14714
rect 8915 14660 8921 14662
rect 8977 14660 9001 14662
rect 9057 14660 9081 14662
rect 9137 14660 9161 14662
rect 9217 14660 9223 14662
rect 8915 14640 9223 14660
rect 7748 14408 7800 14414
rect 7748 14350 7800 14356
rect 10244 13870 10272 16050
rect 10232 13864 10284 13870
rect 10232 13806 10284 13812
rect 8915 13628 9223 13648
rect 8915 13626 8921 13628
rect 8977 13626 9001 13628
rect 9057 13626 9081 13628
rect 9137 13626 9161 13628
rect 9217 13626 9223 13628
rect 8977 13574 8979 13626
rect 9159 13574 9161 13626
rect 8915 13572 8921 13574
rect 8977 13572 9001 13574
rect 9057 13572 9081 13574
rect 9137 13572 9161 13574
rect 9217 13572 9223 13574
rect 8915 13552 9223 13572
rect 8915 12540 9223 12560
rect 8915 12538 8921 12540
rect 8977 12538 9001 12540
rect 9057 12538 9081 12540
rect 9137 12538 9161 12540
rect 9217 12538 9223 12540
rect 8977 12486 8979 12538
rect 9159 12486 9161 12538
rect 8915 12484 8921 12486
rect 8977 12484 9001 12486
rect 9057 12484 9081 12486
rect 9137 12484 9161 12486
rect 9217 12484 9223 12486
rect 8915 12464 9223 12484
rect 8208 11756 8260 11762
rect 8208 11698 8260 11704
rect 5724 5704 5776 5710
rect 5724 5646 5776 5652
rect 5172 5024 5224 5030
rect 5172 4966 5224 4972
rect 5184 4690 5212 4966
rect 5172 4684 5224 4690
rect 5172 4626 5224 4632
rect 5540 4684 5592 4690
rect 5540 4626 5592 4632
rect 4988 4616 5040 4622
rect 4988 4558 5040 4564
rect 5000 4146 5028 4558
rect 4988 4140 5040 4146
rect 4988 4082 5040 4088
rect 5264 4072 5316 4078
rect 5264 4014 5316 4020
rect 5276 3738 5304 4014
rect 5264 3732 5316 3738
rect 5264 3674 5316 3680
rect 5552 3074 5580 4626
rect 5736 3602 5764 5646
rect 6552 5024 6604 5030
rect 6552 4966 6604 4972
rect 6564 4214 6592 4966
rect 7840 4548 7892 4554
rect 7840 4490 7892 4496
rect 6552 4208 6604 4214
rect 6552 4150 6604 4156
rect 7852 4010 7880 4490
rect 7472 4004 7524 4010
rect 7472 3946 7524 3952
rect 7840 4004 7892 4010
rect 7840 3946 7892 3952
rect 5816 3936 5868 3942
rect 5816 3878 5868 3884
rect 5724 3596 5776 3602
rect 5724 3538 5776 3544
rect 5724 3460 5776 3466
rect 5724 3402 5776 3408
rect 5736 3194 5764 3402
rect 5724 3188 5776 3194
rect 5724 3130 5776 3136
rect 4620 3052 4672 3058
rect 4620 2994 4672 3000
rect 5184 3046 5580 3074
rect 3884 2984 3936 2990
rect 3884 2926 3936 2932
rect 2870 2816 2926 2825
rect 2870 2751 2926 2760
rect 3240 2576 3292 2582
rect 3240 2518 3292 2524
rect 2688 2440 2740 2446
rect 2688 2382 2740 2388
rect 3252 800 3280 2518
rect 3516 2372 3568 2378
rect 3516 2314 3568 2320
rect 3424 2304 3476 2310
rect 3424 2246 3476 2252
rect 3436 2145 3464 2246
rect 3422 2136 3478 2145
rect 3422 2071 3478 2080
rect 3528 1465 3556 2314
rect 3514 1456 3570 1465
rect 3514 1391 3570 1400
rect 3896 800 3924 2926
rect 4620 2916 4672 2922
rect 4620 2858 4672 2864
rect 4528 2848 4580 2854
rect 4528 2790 4580 2796
rect 4540 2514 4568 2790
rect 4528 2508 4580 2514
rect 4528 2450 4580 2456
rect 4632 2394 4660 2858
rect 4540 2366 4660 2394
rect 4540 800 4568 2366
rect 5184 800 5212 3046
rect 5540 2984 5592 2990
rect 5540 2926 5592 2932
rect 5552 2650 5580 2926
rect 5540 2644 5592 2650
rect 5540 2586 5592 2592
rect 5828 2514 5856 3878
rect 5908 3596 5960 3602
rect 5908 3538 5960 3544
rect 5816 2508 5868 2514
rect 5816 2450 5868 2456
rect 5920 1850 5948 3538
rect 7484 2990 7512 3946
rect 8220 3534 8248 11698
rect 8915 11452 9223 11472
rect 8915 11450 8921 11452
rect 8977 11450 9001 11452
rect 9057 11450 9081 11452
rect 9137 11450 9161 11452
rect 9217 11450 9223 11452
rect 8977 11398 8979 11450
rect 9159 11398 9161 11450
rect 8915 11396 8921 11398
rect 8977 11396 9001 11398
rect 9057 11396 9081 11398
rect 9137 11396 9161 11398
rect 9217 11396 9223 11398
rect 8915 11376 9223 11396
rect 8915 10364 9223 10384
rect 8915 10362 8921 10364
rect 8977 10362 9001 10364
rect 9057 10362 9081 10364
rect 9137 10362 9161 10364
rect 9217 10362 9223 10364
rect 8977 10310 8979 10362
rect 9159 10310 9161 10362
rect 8915 10308 8921 10310
rect 8977 10308 9001 10310
rect 9057 10308 9081 10310
rect 9137 10308 9161 10310
rect 9217 10308 9223 10310
rect 8915 10288 9223 10308
rect 8915 9276 9223 9296
rect 8915 9274 8921 9276
rect 8977 9274 9001 9276
rect 9057 9274 9081 9276
rect 9137 9274 9161 9276
rect 9217 9274 9223 9276
rect 8977 9222 8979 9274
rect 9159 9222 9161 9274
rect 8915 9220 8921 9222
rect 8977 9220 9001 9222
rect 9057 9220 9081 9222
rect 9137 9220 9161 9222
rect 9217 9220 9223 9222
rect 8915 9200 9223 9220
rect 8915 8188 9223 8208
rect 8915 8186 8921 8188
rect 8977 8186 9001 8188
rect 9057 8186 9081 8188
rect 9137 8186 9161 8188
rect 9217 8186 9223 8188
rect 8977 8134 8979 8186
rect 9159 8134 9161 8186
rect 8915 8132 8921 8134
rect 8977 8132 9001 8134
rect 9057 8132 9081 8134
rect 9137 8132 9161 8134
rect 9217 8132 9223 8134
rect 8915 8112 9223 8132
rect 8915 7100 9223 7120
rect 8915 7098 8921 7100
rect 8977 7098 9001 7100
rect 9057 7098 9081 7100
rect 9137 7098 9161 7100
rect 9217 7098 9223 7100
rect 8977 7046 8979 7098
rect 9159 7046 9161 7098
rect 8915 7044 8921 7046
rect 8977 7044 9001 7046
rect 9057 7044 9081 7046
rect 9137 7044 9161 7046
rect 9217 7044 9223 7046
rect 8915 7024 9223 7044
rect 8915 6012 9223 6032
rect 8915 6010 8921 6012
rect 8977 6010 9001 6012
rect 9057 6010 9081 6012
rect 9137 6010 9161 6012
rect 9217 6010 9223 6012
rect 8977 5958 8979 6010
rect 9159 5958 9161 6010
rect 8915 5956 8921 5958
rect 8977 5956 9001 5958
rect 9057 5956 9081 5958
rect 9137 5956 9161 5958
rect 9217 5956 9223 5958
rect 8915 5936 9223 5956
rect 10244 5302 10272 13806
rect 10324 8288 10376 8294
rect 10324 8230 10376 8236
rect 10336 7954 10364 8230
rect 10980 7954 11008 19200
rect 11624 17270 11652 19200
rect 11612 17264 11664 17270
rect 11612 17206 11664 17212
rect 12164 17060 12216 17066
rect 12164 17002 12216 17008
rect 11704 15904 11756 15910
rect 11704 15846 11756 15852
rect 11716 15570 11744 15846
rect 11704 15564 11756 15570
rect 11704 15506 11756 15512
rect 11888 15428 11940 15434
rect 11888 15370 11940 15376
rect 11900 15162 11928 15370
rect 11888 15156 11940 15162
rect 11888 15098 11940 15104
rect 11796 15020 11848 15026
rect 11796 14962 11848 14968
rect 11808 14890 11836 14962
rect 11796 14884 11848 14890
rect 11796 14826 11848 14832
rect 11060 10464 11112 10470
rect 11060 10406 11112 10412
rect 11072 10130 11100 10406
rect 11060 10124 11112 10130
rect 11060 10066 11112 10072
rect 11244 9988 11296 9994
rect 11244 9930 11296 9936
rect 11256 9722 11284 9930
rect 11244 9716 11296 9722
rect 11244 9658 11296 9664
rect 11808 9586 11836 14826
rect 12176 14346 12204 17002
rect 12268 15570 12296 19200
rect 12348 17536 12400 17542
rect 12348 17478 12400 17484
rect 12360 17066 12388 17478
rect 12348 17060 12400 17066
rect 12348 17002 12400 17008
rect 12440 16584 12492 16590
rect 12440 16526 12492 16532
rect 12452 16250 12480 16526
rect 12440 16244 12492 16250
rect 12440 16186 12492 16192
rect 12912 16046 12940 19200
rect 15568 17264 15620 17270
rect 15568 17206 15620 17212
rect 14280 17128 14332 17134
rect 14280 17070 14332 17076
rect 14292 16522 14320 17070
rect 15580 16794 15608 17206
rect 15660 16992 15712 16998
rect 15660 16934 15712 16940
rect 15672 16794 15700 16934
rect 15568 16788 15620 16794
rect 15568 16730 15620 16736
rect 15660 16788 15712 16794
rect 15660 16730 15712 16736
rect 16132 16658 16160 19200
rect 16120 16652 16172 16658
rect 16120 16594 16172 16600
rect 14280 16516 14332 16522
rect 14280 16458 14332 16464
rect 15752 16516 15804 16522
rect 15752 16458 15804 16464
rect 15764 16250 15792 16458
rect 15752 16244 15804 16250
rect 15752 16186 15804 16192
rect 15568 16108 15620 16114
rect 15568 16050 15620 16056
rect 12532 16040 12584 16046
rect 12532 15982 12584 15988
rect 12900 16040 12952 16046
rect 12900 15982 12952 15988
rect 12256 15564 12308 15570
rect 12256 15506 12308 15512
rect 12544 15162 12572 15982
rect 15580 15638 15608 16050
rect 16120 15904 16172 15910
rect 16120 15846 16172 15852
rect 15568 15632 15620 15638
rect 15568 15574 15620 15580
rect 12532 15156 12584 15162
rect 12532 15098 12584 15104
rect 12440 15020 12492 15026
rect 12440 14962 12492 14968
rect 12452 14822 12480 14962
rect 12440 14816 12492 14822
rect 12440 14758 12492 14764
rect 12164 14340 12216 14346
rect 12164 14282 12216 14288
rect 11796 9580 11848 9586
rect 11796 9522 11848 9528
rect 10324 7948 10376 7954
rect 10324 7890 10376 7896
rect 10968 7948 11020 7954
rect 10968 7890 11020 7896
rect 10508 7812 10560 7818
rect 10508 7754 10560 7760
rect 10520 7546 10548 7754
rect 10508 7540 10560 7546
rect 10508 7482 10560 7488
rect 10416 7404 10468 7410
rect 10416 7346 10468 7352
rect 10232 5296 10284 5302
rect 10232 5238 10284 5244
rect 8300 5228 8352 5234
rect 8300 5170 8352 5176
rect 8312 4146 8340 5170
rect 8915 4924 9223 4944
rect 8915 4922 8921 4924
rect 8977 4922 9001 4924
rect 9057 4922 9081 4924
rect 9137 4922 9161 4924
rect 9217 4922 9223 4924
rect 8977 4870 8979 4922
rect 9159 4870 9161 4922
rect 8915 4868 8921 4870
rect 8977 4868 9001 4870
rect 9057 4868 9081 4870
rect 9137 4868 9161 4870
rect 9217 4868 9223 4870
rect 8915 4848 9223 4868
rect 8760 4616 8812 4622
rect 8760 4558 8812 4564
rect 8300 4140 8352 4146
rect 8300 4082 8352 4088
rect 8208 3528 8260 3534
rect 8208 3470 8260 3476
rect 8116 3392 8168 3398
rect 8116 3334 8168 3340
rect 8300 3392 8352 3398
rect 8300 3334 8352 3340
rect 8128 3194 8156 3334
rect 8116 3188 8168 3194
rect 8116 3130 8168 3136
rect 7472 2984 7524 2990
rect 7472 2926 7524 2932
rect 6736 2916 6788 2922
rect 6736 2858 6788 2864
rect 6552 2848 6604 2854
rect 6552 2790 6604 2796
rect 6564 2514 6592 2790
rect 6748 2514 6776 2858
rect 7748 2576 7800 2582
rect 7748 2518 7800 2524
rect 6552 2508 6604 2514
rect 6552 2450 6604 2456
rect 6736 2508 6788 2514
rect 6736 2450 6788 2456
rect 5828 1822 5948 1850
rect 5828 800 5856 1822
rect 7760 800 7788 2518
rect 8312 2378 8340 3334
rect 8772 2514 8800 4558
rect 10428 4554 10456 7346
rect 9956 4548 10008 4554
rect 9956 4490 10008 4496
rect 10416 4548 10468 4554
rect 10416 4490 10468 4496
rect 9312 3936 9364 3942
rect 9312 3878 9364 3884
rect 9864 3936 9916 3942
rect 9864 3878 9916 3884
rect 8915 3836 9223 3856
rect 8915 3834 8921 3836
rect 8977 3834 9001 3836
rect 9057 3834 9081 3836
rect 9137 3834 9161 3836
rect 9217 3834 9223 3836
rect 8977 3782 8979 3834
rect 9159 3782 9161 3834
rect 8915 3780 8921 3782
rect 8977 3780 9001 3782
rect 9057 3780 9081 3782
rect 9137 3780 9161 3782
rect 9217 3780 9223 3782
rect 8915 3760 9223 3780
rect 9324 3602 9352 3878
rect 9876 3670 9904 3878
rect 9968 3670 9996 4490
rect 11612 3936 11664 3942
rect 11612 3878 11664 3884
rect 9864 3664 9916 3670
rect 9864 3606 9916 3612
rect 9956 3664 10008 3670
rect 9956 3606 10008 3612
rect 11624 3602 11652 3878
rect 11704 3732 11756 3738
rect 11704 3674 11756 3680
rect 9312 3596 9364 3602
rect 9312 3538 9364 3544
rect 9680 3596 9732 3602
rect 9680 3538 9732 3544
rect 11612 3596 11664 3602
rect 11612 3538 11664 3544
rect 9312 2984 9364 2990
rect 9312 2926 9364 2932
rect 8915 2748 9223 2768
rect 8915 2746 8921 2748
rect 8977 2746 9001 2748
rect 9057 2746 9081 2748
rect 9137 2746 9161 2748
rect 9217 2746 9223 2748
rect 8977 2694 8979 2746
rect 9159 2694 9161 2746
rect 8915 2692 8921 2694
rect 8977 2692 9001 2694
rect 9057 2692 9081 2694
rect 9137 2692 9161 2694
rect 9217 2692 9223 2694
rect 8915 2672 9223 2692
rect 8760 2508 8812 2514
rect 8760 2450 8812 2456
rect 8208 2372 8260 2378
rect 8208 2314 8260 2320
rect 8300 2372 8352 2378
rect 8300 2314 8352 2320
rect 8220 2106 8248 2314
rect 8208 2100 8260 2106
rect 8208 2042 8260 2048
rect 9324 1578 9352 2926
rect 9048 1550 9352 1578
rect 9048 800 9076 1550
rect 9692 800 9720 3538
rect 11716 3058 11744 3674
rect 12256 3596 12308 3602
rect 12256 3538 12308 3544
rect 11796 3460 11848 3466
rect 11796 3402 11848 3408
rect 11808 3194 11836 3402
rect 11796 3188 11848 3194
rect 11796 3130 11848 3136
rect 11704 3052 11756 3058
rect 11704 2994 11756 3000
rect 12268 800 12296 3538
rect 12452 2922 12480 14758
rect 12992 10464 13044 10470
rect 12992 10406 13044 10412
rect 13004 9586 13032 10406
rect 13176 9920 13228 9926
rect 13176 9862 13228 9868
rect 13188 9654 13216 9862
rect 13176 9648 13228 9654
rect 13176 9590 13228 9596
rect 12992 9580 13044 9586
rect 12992 9522 13044 9528
rect 13544 9512 13596 9518
rect 13544 9454 13596 9460
rect 13176 4004 13228 4010
rect 13176 3946 13228 3952
rect 12532 3936 12584 3942
rect 12532 3878 12584 3884
rect 12440 2916 12492 2922
rect 12440 2858 12492 2864
rect 12544 2582 12572 3878
rect 13188 3670 13216 3946
rect 13176 3664 13228 3670
rect 13176 3606 13228 3612
rect 13360 2848 13412 2854
rect 13360 2790 13412 2796
rect 12532 2576 12584 2582
rect 12532 2518 12584 2524
rect 13372 2514 13400 2790
rect 13360 2508 13412 2514
rect 13360 2450 13412 2456
rect 13556 800 13584 9454
rect 15108 4140 15160 4146
rect 15108 4082 15160 4088
rect 14188 3936 14240 3942
rect 14188 3878 14240 3884
rect 13820 2984 13872 2990
rect 13820 2926 13872 2932
rect 13832 2106 13860 2926
rect 14200 2514 14228 3878
rect 15120 3534 15148 4082
rect 15476 4004 15528 4010
rect 15476 3946 15528 3952
rect 15108 3528 15160 3534
rect 15108 3470 15160 3476
rect 14372 3392 14424 3398
rect 14372 3334 14424 3340
rect 15292 3392 15344 3398
rect 15292 3334 15344 3340
rect 14384 2514 14412 3334
rect 15304 3126 15332 3334
rect 15292 3120 15344 3126
rect 15292 3062 15344 3068
rect 15488 3058 15516 3946
rect 15476 3052 15528 3058
rect 15476 2994 15528 3000
rect 15580 2990 15608 15574
rect 16132 15570 16160 15846
rect 16776 15570 16804 19200
rect 16880 17436 17188 17456
rect 16880 17434 16886 17436
rect 16942 17434 16966 17436
rect 17022 17434 17046 17436
rect 17102 17434 17126 17436
rect 17182 17434 17188 17436
rect 16942 17382 16944 17434
rect 17124 17382 17126 17434
rect 16880 17380 16886 17382
rect 16942 17380 16966 17382
rect 17022 17380 17046 17382
rect 17102 17380 17126 17382
rect 17182 17380 17188 17382
rect 16880 17360 17188 17380
rect 18064 17134 18092 19200
rect 18144 17332 18196 17338
rect 18144 17274 18196 17280
rect 18052 17128 18104 17134
rect 18052 17070 18104 17076
rect 17132 16992 17184 16998
rect 17132 16934 17184 16940
rect 17144 16726 17172 16934
rect 17132 16720 17184 16726
rect 17132 16662 17184 16668
rect 17960 16652 18012 16658
rect 17960 16594 18012 16600
rect 16880 16348 17188 16368
rect 16880 16346 16886 16348
rect 16942 16346 16966 16348
rect 17022 16346 17046 16348
rect 17102 16346 17126 16348
rect 17182 16346 17188 16348
rect 16942 16294 16944 16346
rect 17124 16294 17126 16346
rect 16880 16292 16886 16294
rect 16942 16292 16966 16294
rect 17022 16292 17046 16294
rect 17102 16292 17126 16294
rect 17182 16292 17188 16294
rect 16880 16272 17188 16292
rect 16120 15564 16172 15570
rect 16120 15506 16172 15512
rect 16764 15564 16816 15570
rect 16764 15506 16816 15512
rect 15660 15496 15712 15502
rect 15660 15438 15712 15444
rect 15672 14958 15700 15438
rect 16880 15260 17188 15280
rect 16880 15258 16886 15260
rect 16942 15258 16966 15260
rect 17022 15258 17046 15260
rect 17102 15258 17126 15260
rect 17182 15258 17188 15260
rect 16942 15206 16944 15258
rect 17124 15206 17126 15258
rect 16880 15204 16886 15206
rect 16942 15204 16966 15206
rect 17022 15204 17046 15206
rect 17102 15204 17126 15206
rect 17182 15204 17188 15206
rect 16880 15184 17188 15204
rect 17972 15162 18000 16594
rect 18156 16590 18184 17274
rect 18512 17128 18564 17134
rect 18512 17070 18564 17076
rect 18524 16794 18552 17070
rect 18512 16788 18564 16794
rect 18512 16730 18564 16736
rect 18144 16584 18196 16590
rect 18144 16526 18196 16532
rect 18236 16584 18288 16590
rect 18236 16526 18288 16532
rect 17960 15156 18012 15162
rect 17960 15098 18012 15104
rect 18052 15088 18104 15094
rect 18052 15030 18104 15036
rect 15660 14952 15712 14958
rect 15660 14894 15712 14900
rect 18064 14822 18092 15030
rect 18052 14816 18104 14822
rect 18052 14758 18104 14764
rect 18156 14634 18184 16526
rect 18248 16114 18276 16526
rect 18236 16108 18288 16114
rect 18236 16050 18288 16056
rect 18708 16046 18736 19200
rect 22192 17128 22244 17134
rect 22192 17070 22244 17076
rect 19892 17060 19944 17066
rect 19892 17002 19944 17008
rect 19708 16992 19760 16998
rect 19708 16934 19760 16940
rect 18512 16040 18564 16046
rect 18512 15982 18564 15988
rect 18696 16040 18748 16046
rect 18696 15982 18748 15988
rect 19248 16040 19300 16046
rect 19248 15982 19300 15988
rect 18524 15706 18552 15982
rect 18512 15700 18564 15706
rect 18512 15642 18564 15648
rect 19260 15502 19288 15982
rect 19616 15972 19668 15978
rect 19616 15914 19668 15920
rect 18420 15496 18472 15502
rect 18420 15438 18472 15444
rect 19248 15496 19300 15502
rect 19248 15438 19300 15444
rect 18328 15156 18380 15162
rect 18328 15098 18380 15104
rect 18340 14958 18368 15098
rect 18328 14952 18380 14958
rect 18328 14894 18380 14900
rect 17972 14606 18184 14634
rect 16880 14172 17188 14192
rect 16880 14170 16886 14172
rect 16942 14170 16966 14172
rect 17022 14170 17046 14172
rect 17102 14170 17126 14172
rect 17182 14170 17188 14172
rect 16942 14118 16944 14170
rect 17124 14118 17126 14170
rect 16880 14116 16886 14118
rect 16942 14116 16966 14118
rect 17022 14116 17046 14118
rect 17102 14116 17126 14118
rect 17182 14116 17188 14118
rect 16880 14096 17188 14116
rect 16880 13084 17188 13104
rect 16880 13082 16886 13084
rect 16942 13082 16966 13084
rect 17022 13082 17046 13084
rect 17102 13082 17126 13084
rect 17182 13082 17188 13084
rect 16942 13030 16944 13082
rect 17124 13030 17126 13082
rect 16880 13028 16886 13030
rect 16942 13028 16966 13030
rect 17022 13028 17046 13030
rect 17102 13028 17126 13030
rect 17182 13028 17188 13030
rect 16880 13008 17188 13028
rect 16880 11996 17188 12016
rect 16880 11994 16886 11996
rect 16942 11994 16966 11996
rect 17022 11994 17046 11996
rect 17102 11994 17126 11996
rect 17182 11994 17188 11996
rect 16942 11942 16944 11994
rect 17124 11942 17126 11994
rect 16880 11940 16886 11942
rect 16942 11940 16966 11942
rect 17022 11940 17046 11942
rect 17102 11940 17126 11942
rect 17182 11940 17188 11942
rect 16880 11920 17188 11940
rect 16880 10908 17188 10928
rect 16880 10906 16886 10908
rect 16942 10906 16966 10908
rect 17022 10906 17046 10908
rect 17102 10906 17126 10908
rect 17182 10906 17188 10908
rect 16942 10854 16944 10906
rect 17124 10854 17126 10906
rect 16880 10852 16886 10854
rect 16942 10852 16966 10854
rect 17022 10852 17046 10854
rect 17102 10852 17126 10854
rect 17182 10852 17188 10854
rect 16880 10832 17188 10852
rect 16880 9820 17188 9840
rect 16880 9818 16886 9820
rect 16942 9818 16966 9820
rect 17022 9818 17046 9820
rect 17102 9818 17126 9820
rect 17182 9818 17188 9820
rect 16942 9766 16944 9818
rect 17124 9766 17126 9818
rect 16880 9764 16886 9766
rect 16942 9764 16966 9766
rect 17022 9764 17046 9766
rect 17102 9764 17126 9766
rect 17182 9764 17188 9766
rect 16880 9744 17188 9764
rect 16880 8732 17188 8752
rect 16880 8730 16886 8732
rect 16942 8730 16966 8732
rect 17022 8730 17046 8732
rect 17102 8730 17126 8732
rect 17182 8730 17188 8732
rect 16942 8678 16944 8730
rect 17124 8678 17126 8730
rect 16880 8676 16886 8678
rect 16942 8676 16966 8678
rect 17022 8676 17046 8678
rect 17102 8676 17126 8678
rect 17182 8676 17188 8678
rect 16880 8656 17188 8676
rect 17684 7880 17736 7886
rect 17684 7822 17736 7828
rect 16880 7644 17188 7664
rect 16880 7642 16886 7644
rect 16942 7642 16966 7644
rect 17022 7642 17046 7644
rect 17102 7642 17126 7644
rect 17182 7642 17188 7644
rect 16942 7590 16944 7642
rect 17124 7590 17126 7642
rect 16880 7588 16886 7590
rect 16942 7588 16966 7590
rect 17022 7588 17046 7590
rect 17102 7588 17126 7590
rect 17182 7588 17188 7590
rect 16880 7568 17188 7588
rect 17696 7410 17724 7822
rect 17684 7404 17736 7410
rect 17684 7346 17736 7352
rect 16880 6556 17188 6576
rect 16880 6554 16886 6556
rect 16942 6554 16966 6556
rect 17022 6554 17046 6556
rect 17102 6554 17126 6556
rect 17182 6554 17188 6556
rect 16942 6502 16944 6554
rect 17124 6502 17126 6554
rect 16880 6500 16886 6502
rect 16942 6500 16966 6502
rect 17022 6500 17046 6502
rect 17102 6500 17126 6502
rect 17182 6500 17188 6502
rect 16880 6480 17188 6500
rect 16880 5468 17188 5488
rect 16880 5466 16886 5468
rect 16942 5466 16966 5468
rect 17022 5466 17046 5468
rect 17102 5466 17126 5468
rect 17182 5466 17188 5468
rect 16942 5414 16944 5466
rect 17124 5414 17126 5466
rect 16880 5412 16886 5414
rect 16942 5412 16966 5414
rect 17022 5412 17046 5414
rect 17102 5412 17126 5414
rect 17182 5412 17188 5414
rect 16880 5392 17188 5412
rect 15752 4616 15804 4622
rect 15752 4558 15804 4564
rect 15764 3602 15792 4558
rect 16880 4380 17188 4400
rect 16880 4378 16886 4380
rect 16942 4378 16966 4380
rect 17022 4378 17046 4380
rect 17102 4378 17126 4380
rect 17182 4378 17188 4380
rect 16942 4326 16944 4378
rect 17124 4326 17126 4378
rect 16880 4324 16886 4326
rect 16942 4324 16966 4326
rect 17022 4324 17046 4326
rect 17102 4324 17126 4326
rect 17182 4324 17188 4326
rect 16880 4304 17188 4324
rect 17972 4146 18000 14606
rect 18340 10062 18368 14894
rect 18328 10056 18380 10062
rect 18328 9998 18380 10004
rect 18052 7336 18104 7342
rect 18052 7278 18104 7284
rect 18064 6866 18092 7278
rect 18052 6860 18104 6866
rect 18052 6802 18104 6808
rect 18432 6798 18460 15438
rect 19432 15428 19484 15434
rect 19432 15370 19484 15376
rect 18512 15020 18564 15026
rect 18512 14962 18564 14968
rect 18524 14618 18552 14962
rect 18512 14612 18564 14618
rect 18512 14554 18564 14560
rect 18420 6792 18472 6798
rect 18420 6734 18472 6740
rect 17960 4140 18012 4146
rect 17960 4082 18012 4088
rect 18696 4072 18748 4078
rect 18696 4014 18748 4020
rect 19340 4072 19392 4078
rect 19340 4014 19392 4020
rect 15936 3936 15988 3942
rect 15936 3878 15988 3884
rect 18144 3936 18196 3942
rect 18144 3878 18196 3884
rect 15948 3602 15976 3878
rect 15752 3596 15804 3602
rect 15752 3538 15804 3544
rect 15936 3596 15988 3602
rect 15936 3538 15988 3544
rect 16120 3596 16172 3602
rect 16120 3538 16172 3544
rect 15568 2984 15620 2990
rect 15568 2926 15620 2932
rect 16028 2848 16080 2854
rect 16028 2790 16080 2796
rect 14188 2508 14240 2514
rect 14188 2450 14240 2456
rect 14372 2508 14424 2514
rect 14372 2450 14424 2456
rect 14832 2508 14884 2514
rect 14832 2450 14884 2456
rect 13820 2100 13872 2106
rect 13820 2042 13872 2048
rect 14844 800 14872 2450
rect 16040 2378 16068 2790
rect 16028 2372 16080 2378
rect 16028 2314 16080 2320
rect 16132 800 16160 3538
rect 16880 3292 17188 3312
rect 16880 3290 16886 3292
rect 16942 3290 16966 3292
rect 17022 3290 17046 3292
rect 17102 3290 17126 3292
rect 17182 3290 17188 3292
rect 16942 3238 16944 3290
rect 17124 3238 17126 3290
rect 16880 3236 16886 3238
rect 16942 3236 16966 3238
rect 17022 3236 17046 3238
rect 17102 3236 17126 3238
rect 17182 3236 17188 3238
rect 16880 3216 17188 3236
rect 18052 3188 18104 3194
rect 18052 3130 18104 3136
rect 16672 2848 16724 2854
rect 16672 2790 16724 2796
rect 16684 2514 16712 2790
rect 16672 2508 16724 2514
rect 16672 2450 16724 2456
rect 16880 2204 17188 2224
rect 16880 2202 16886 2204
rect 16942 2202 16966 2204
rect 17022 2202 17046 2204
rect 17102 2202 17126 2204
rect 17182 2202 17188 2204
rect 16942 2150 16944 2202
rect 17124 2150 17126 2202
rect 16880 2148 16886 2150
rect 16942 2148 16966 2150
rect 17022 2148 17046 2150
rect 17102 2148 17126 2150
rect 17182 2148 17188 2150
rect 16880 2128 17188 2148
rect 18064 800 18092 3130
rect 18156 3126 18184 3878
rect 18328 3392 18380 3398
rect 18328 3334 18380 3340
rect 18340 3126 18368 3334
rect 18144 3120 18196 3126
rect 18144 3062 18196 3068
rect 18328 3120 18380 3126
rect 18328 3062 18380 3068
rect 18708 800 18736 4014
rect 19352 3738 19380 4014
rect 19340 3732 19392 3738
rect 19340 3674 19392 3680
rect 19444 3670 19472 15370
rect 19628 14482 19656 15914
rect 19720 14958 19748 16934
rect 19904 16726 19932 17002
rect 20168 16992 20220 16998
rect 20168 16934 20220 16940
rect 19892 16720 19944 16726
rect 19892 16662 19944 16668
rect 20180 16658 20208 16934
rect 22204 16794 22232 17070
rect 22192 16788 22244 16794
rect 22192 16730 22244 16736
rect 20168 16652 20220 16658
rect 20168 16594 20220 16600
rect 22572 16522 22600 19200
rect 23860 17270 23888 19200
rect 24504 17898 24532 19200
rect 25148 17898 25176 19200
rect 24504 17870 24900 17898
rect 25148 17870 25268 17898
rect 24492 17332 24544 17338
rect 24492 17274 24544 17280
rect 23848 17264 23900 17270
rect 23848 17206 23900 17212
rect 24400 17128 24452 17134
rect 24400 17070 24452 17076
rect 22560 16516 22612 16522
rect 22560 16458 22612 16464
rect 22100 16176 22152 16182
rect 22100 16118 22152 16124
rect 22112 15638 22140 16118
rect 24412 16114 24440 17070
rect 24400 16108 24452 16114
rect 24400 16050 24452 16056
rect 22100 15632 22152 15638
rect 22100 15574 22152 15580
rect 19892 15496 19944 15502
rect 19892 15438 19944 15444
rect 19904 15026 19932 15438
rect 19892 15020 19944 15026
rect 19892 14962 19944 14968
rect 24504 14958 24532 17274
rect 24872 17134 24900 17870
rect 24584 17128 24636 17134
rect 24584 17070 24636 17076
rect 24860 17128 24912 17134
rect 24860 17070 24912 17076
rect 24596 16794 24624 17070
rect 24846 16892 25154 16912
rect 24846 16890 24852 16892
rect 24908 16890 24932 16892
rect 24988 16890 25012 16892
rect 25068 16890 25092 16892
rect 25148 16890 25154 16892
rect 24908 16838 24910 16890
rect 25090 16838 25092 16890
rect 24846 16836 24852 16838
rect 24908 16836 24932 16838
rect 24988 16836 25012 16838
rect 25068 16836 25092 16838
rect 25148 16836 25154 16838
rect 24846 16816 25154 16836
rect 24584 16788 24636 16794
rect 24584 16730 24636 16736
rect 24676 16788 24728 16794
rect 24676 16730 24728 16736
rect 24688 16590 24716 16730
rect 25136 16652 25188 16658
rect 25136 16594 25188 16600
rect 24676 16584 24728 16590
rect 24676 16526 24728 16532
rect 24584 16516 24636 16522
rect 24584 16458 24636 16464
rect 24596 16250 24624 16458
rect 24584 16244 24636 16250
rect 24584 16186 24636 16192
rect 24676 16108 24728 16114
rect 24676 16050 24728 16056
rect 24584 15428 24636 15434
rect 24584 15370 24636 15376
rect 24596 14958 24624 15370
rect 24688 15366 24716 16050
rect 25148 15994 25176 16594
rect 25240 16590 25268 17870
rect 25228 16584 25280 16590
rect 25228 16526 25280 16532
rect 25320 16040 25372 16046
rect 25148 15966 25268 15994
rect 25320 15982 25372 15988
rect 24846 15804 25154 15824
rect 24846 15802 24852 15804
rect 24908 15802 24932 15804
rect 24988 15802 25012 15804
rect 25068 15802 25092 15804
rect 25148 15802 25154 15804
rect 24908 15750 24910 15802
rect 25090 15750 25092 15802
rect 24846 15748 24852 15750
rect 24908 15748 24932 15750
rect 24988 15748 25012 15750
rect 25068 15748 25092 15750
rect 25148 15748 25154 15750
rect 24846 15728 25154 15748
rect 25240 15570 25268 15966
rect 25228 15564 25280 15570
rect 25228 15506 25280 15512
rect 24676 15360 24728 15366
rect 24676 15302 24728 15308
rect 24688 15026 24716 15302
rect 24676 15020 24728 15026
rect 24676 14962 24728 14968
rect 25228 15020 25280 15026
rect 25228 14962 25280 14968
rect 19708 14952 19760 14958
rect 19708 14894 19760 14900
rect 20628 14952 20680 14958
rect 20628 14894 20680 14900
rect 24492 14952 24544 14958
rect 24492 14894 24544 14900
rect 24584 14952 24636 14958
rect 24584 14894 24636 14900
rect 19616 14476 19668 14482
rect 19616 14418 19668 14424
rect 19628 6914 19656 14418
rect 19536 6886 19656 6914
rect 19432 3664 19484 3670
rect 19432 3606 19484 3612
rect 19156 3528 19208 3534
rect 19536 3482 19564 6886
rect 19720 3670 19748 14894
rect 20640 14822 20668 14894
rect 24504 14822 24532 14894
rect 20628 14816 20680 14822
rect 20628 14758 20680 14764
rect 24492 14816 24544 14822
rect 24492 14758 24544 14764
rect 20640 8974 20668 14758
rect 24596 14278 24624 14894
rect 24846 14716 25154 14736
rect 24846 14714 24852 14716
rect 24908 14714 24932 14716
rect 24988 14714 25012 14716
rect 25068 14714 25092 14716
rect 25148 14714 25154 14716
rect 24908 14662 24910 14714
rect 25090 14662 25092 14714
rect 24846 14660 24852 14662
rect 24908 14660 24932 14662
rect 24988 14660 25012 14662
rect 25068 14660 25092 14662
rect 25148 14660 25154 14662
rect 24846 14640 25154 14660
rect 25240 14414 25268 14962
rect 25228 14408 25280 14414
rect 25228 14350 25280 14356
rect 24584 14272 24636 14278
rect 24584 14214 24636 14220
rect 25240 13938 25268 14350
rect 25228 13932 25280 13938
rect 25228 13874 25280 13880
rect 24846 13628 25154 13648
rect 24846 13626 24852 13628
rect 24908 13626 24932 13628
rect 24988 13626 25012 13628
rect 25068 13626 25092 13628
rect 25148 13626 25154 13628
rect 24908 13574 24910 13626
rect 25090 13574 25092 13626
rect 24846 13572 24852 13574
rect 24908 13572 24932 13574
rect 24988 13572 25012 13574
rect 25068 13572 25092 13574
rect 25148 13572 25154 13574
rect 24846 13552 25154 13572
rect 24846 12540 25154 12560
rect 24846 12538 24852 12540
rect 24908 12538 24932 12540
rect 24988 12538 25012 12540
rect 25068 12538 25092 12540
rect 25148 12538 25154 12540
rect 24908 12486 24910 12538
rect 25090 12486 25092 12538
rect 24846 12484 24852 12486
rect 24908 12484 24932 12486
rect 24988 12484 25012 12486
rect 25068 12484 25092 12486
rect 25148 12484 25154 12486
rect 24846 12464 25154 12484
rect 24846 11452 25154 11472
rect 24846 11450 24852 11452
rect 24908 11450 24932 11452
rect 24988 11450 25012 11452
rect 25068 11450 25092 11452
rect 25148 11450 25154 11452
rect 24908 11398 24910 11450
rect 25090 11398 25092 11450
rect 24846 11396 24852 11398
rect 24908 11396 24932 11398
rect 24988 11396 25012 11398
rect 25068 11396 25092 11398
rect 25148 11396 25154 11398
rect 24846 11376 25154 11396
rect 24846 10364 25154 10384
rect 24846 10362 24852 10364
rect 24908 10362 24932 10364
rect 24988 10362 25012 10364
rect 25068 10362 25092 10364
rect 25148 10362 25154 10364
rect 24908 10310 24910 10362
rect 25090 10310 25092 10362
rect 24846 10308 24852 10310
rect 24908 10308 24932 10310
rect 24988 10308 25012 10310
rect 25068 10308 25092 10310
rect 25148 10308 25154 10310
rect 24846 10288 25154 10308
rect 25332 9654 25360 15982
rect 25412 15904 25464 15910
rect 25412 15846 25464 15852
rect 25424 15570 25452 15846
rect 25792 15570 25820 19200
rect 30944 17134 30972 19200
rect 32232 17490 32260 19200
rect 32876 17898 32904 19200
rect 32692 17870 32904 17898
rect 32232 17462 32444 17490
rect 31392 17264 31444 17270
rect 31392 17206 31444 17212
rect 27160 17128 27212 17134
rect 27160 17070 27212 17076
rect 27620 17128 27672 17134
rect 27620 17070 27672 17076
rect 29920 17128 29972 17134
rect 29920 17070 29972 17076
rect 30932 17128 30984 17134
rect 30932 17070 30984 17076
rect 27172 16794 27200 17070
rect 26792 16788 26844 16794
rect 26792 16730 26844 16736
rect 27160 16788 27212 16794
rect 27160 16730 27212 16736
rect 25412 15564 25464 15570
rect 25412 15506 25464 15512
rect 25780 15564 25832 15570
rect 25780 15506 25832 15512
rect 25872 15088 25924 15094
rect 25872 15030 25924 15036
rect 25780 14408 25832 14414
rect 25780 14350 25832 14356
rect 25320 9648 25372 9654
rect 25320 9590 25372 9596
rect 24846 9276 25154 9296
rect 24846 9274 24852 9276
rect 24908 9274 24932 9276
rect 24988 9274 25012 9276
rect 25068 9274 25092 9276
rect 25148 9274 25154 9276
rect 24908 9222 24910 9274
rect 25090 9222 25092 9274
rect 24846 9220 24852 9222
rect 24908 9220 24932 9222
rect 24988 9220 25012 9222
rect 25068 9220 25092 9222
rect 25148 9220 25154 9222
rect 24846 9200 25154 9220
rect 20628 8968 20680 8974
rect 20628 8910 20680 8916
rect 24846 8188 25154 8208
rect 24846 8186 24852 8188
rect 24908 8186 24932 8188
rect 24988 8186 25012 8188
rect 25068 8186 25092 8188
rect 25148 8186 25154 8188
rect 24908 8134 24910 8186
rect 25090 8134 25092 8186
rect 24846 8132 24852 8134
rect 24908 8132 24932 8134
rect 24988 8132 25012 8134
rect 25068 8132 25092 8134
rect 25148 8132 25154 8134
rect 24846 8112 25154 8132
rect 24846 7100 25154 7120
rect 24846 7098 24852 7100
rect 24908 7098 24932 7100
rect 24988 7098 25012 7100
rect 25068 7098 25092 7100
rect 25148 7098 25154 7100
rect 24908 7046 24910 7098
rect 25090 7046 25092 7098
rect 24846 7044 24852 7046
rect 24908 7044 24932 7046
rect 24988 7044 25012 7046
rect 25068 7044 25092 7046
rect 25148 7044 25154 7046
rect 24846 7024 25154 7044
rect 24846 6012 25154 6032
rect 24846 6010 24852 6012
rect 24908 6010 24932 6012
rect 24988 6010 25012 6012
rect 25068 6010 25092 6012
rect 25148 6010 25154 6012
rect 24908 5958 24910 6010
rect 25090 5958 25092 6010
rect 24846 5956 24852 5958
rect 24908 5956 24932 5958
rect 24988 5956 25012 5958
rect 25068 5956 25092 5958
rect 25148 5956 25154 5958
rect 24846 5936 25154 5956
rect 24846 4924 25154 4944
rect 24846 4922 24852 4924
rect 24908 4922 24932 4924
rect 24988 4922 25012 4924
rect 25068 4922 25092 4924
rect 25148 4922 25154 4924
rect 24908 4870 24910 4922
rect 25090 4870 25092 4922
rect 24846 4868 24852 4870
rect 24908 4868 24932 4870
rect 24988 4868 25012 4870
rect 25068 4868 25092 4870
rect 25148 4868 25154 4870
rect 24846 4848 25154 4868
rect 20168 4140 20220 4146
rect 20168 4082 20220 4088
rect 20076 4072 20128 4078
rect 20076 4014 20128 4020
rect 20088 3738 20116 4014
rect 20076 3732 20128 3738
rect 20076 3674 20128 3680
rect 19708 3664 19760 3670
rect 19708 3606 19760 3612
rect 20180 3534 20208 4082
rect 25504 4072 25556 4078
rect 25504 4014 25556 4020
rect 24846 3836 25154 3856
rect 24846 3834 24852 3836
rect 24908 3834 24932 3836
rect 24988 3834 25012 3836
rect 25068 3834 25092 3836
rect 25148 3834 25154 3836
rect 24908 3782 24910 3834
rect 25090 3782 25092 3834
rect 24846 3780 24852 3782
rect 24908 3780 24932 3782
rect 24988 3780 25012 3782
rect 25068 3780 25092 3782
rect 25148 3780 25154 3782
rect 24846 3760 25154 3780
rect 25516 3534 25544 4014
rect 25792 3942 25820 14350
rect 25780 3936 25832 3942
rect 25780 3878 25832 3884
rect 19208 3476 19564 3482
rect 19156 3470 19564 3476
rect 20168 3528 20220 3534
rect 20168 3470 20220 3476
rect 23940 3528 23992 3534
rect 23940 3470 23992 3476
rect 25504 3528 25556 3534
rect 25504 3470 25556 3476
rect 19168 3454 19564 3470
rect 20444 3460 20496 3466
rect 19352 3126 19380 3454
rect 20444 3402 20496 3408
rect 19340 3120 19392 3126
rect 19340 3062 19392 3068
rect 20456 3058 20484 3402
rect 23952 3058 23980 3470
rect 24124 3392 24176 3398
rect 24124 3334 24176 3340
rect 24136 3126 24164 3334
rect 24124 3120 24176 3126
rect 24124 3062 24176 3068
rect 20444 3052 20496 3058
rect 20444 2994 20496 3000
rect 23756 3052 23808 3058
rect 23756 2994 23808 3000
rect 23940 3052 23992 3058
rect 23940 2994 23992 3000
rect 19340 2984 19392 2990
rect 19340 2926 19392 2932
rect 19352 800 19380 2926
rect 23768 2922 23796 2994
rect 23664 2916 23716 2922
rect 23664 2858 23716 2864
rect 23756 2916 23808 2922
rect 23756 2858 23808 2864
rect 21088 2848 21140 2854
rect 21088 2790 21140 2796
rect 21272 2848 21324 2854
rect 21272 2790 21324 2796
rect 21100 2514 21128 2790
rect 21284 2514 21312 2790
rect 23676 2514 23704 2858
rect 23848 2848 23900 2854
rect 23848 2790 23900 2796
rect 23860 2514 23888 2790
rect 24846 2748 25154 2768
rect 24846 2746 24852 2748
rect 24908 2746 24932 2748
rect 24988 2746 25012 2748
rect 25068 2746 25092 2748
rect 25148 2746 25154 2748
rect 24908 2694 24910 2746
rect 25090 2694 25092 2746
rect 24846 2692 24852 2694
rect 24908 2692 24932 2694
rect 24988 2692 25012 2694
rect 25068 2692 25092 2694
rect 25148 2692 25154 2694
rect 24846 2672 25154 2692
rect 25884 2582 25912 15030
rect 26804 13394 26832 16730
rect 27632 16590 27660 17070
rect 29932 16794 29960 17070
rect 30564 17060 30616 17066
rect 30564 17002 30616 17008
rect 30576 16794 30604 17002
rect 29920 16788 29972 16794
rect 29920 16730 29972 16736
rect 30564 16788 30616 16794
rect 30564 16730 30616 16736
rect 27896 16720 27948 16726
rect 27896 16662 27948 16668
rect 27068 16584 27120 16590
rect 27068 16526 27120 16532
rect 27528 16584 27580 16590
rect 27528 16526 27580 16532
rect 27620 16584 27672 16590
rect 27620 16526 27672 16532
rect 27080 16114 27108 16526
rect 27068 16108 27120 16114
rect 27068 16050 27120 16056
rect 26976 15972 27028 15978
rect 26976 15914 27028 15920
rect 26988 14414 27016 15914
rect 27540 15162 27568 16526
rect 27712 15496 27764 15502
rect 27712 15438 27764 15444
rect 27528 15156 27580 15162
rect 27528 15098 27580 15104
rect 27620 15156 27672 15162
rect 27620 15098 27672 15104
rect 27632 14822 27660 15098
rect 27724 14822 27752 15438
rect 27804 14952 27856 14958
rect 27804 14894 27856 14900
rect 27620 14816 27672 14822
rect 27620 14758 27672 14764
rect 27712 14816 27764 14822
rect 27712 14758 27764 14764
rect 26976 14408 27028 14414
rect 26976 14350 27028 14356
rect 26792 13388 26844 13394
rect 26792 13330 26844 13336
rect 26988 3670 27016 14350
rect 27436 13388 27488 13394
rect 27436 13330 27488 13336
rect 27448 13258 27476 13330
rect 27620 13320 27672 13326
rect 27620 13262 27672 13268
rect 27436 13252 27488 13258
rect 27436 13194 27488 13200
rect 27344 12776 27396 12782
rect 27344 12718 27396 12724
rect 27356 11762 27384 12718
rect 27344 11756 27396 11762
rect 27344 11698 27396 11704
rect 27252 4072 27304 4078
rect 27252 4014 27304 4020
rect 26976 3664 27028 3670
rect 26976 3606 27028 3612
rect 26240 3392 26292 3398
rect 26240 3334 26292 3340
rect 25872 2576 25924 2582
rect 25872 2518 25924 2524
rect 26252 2514 26280 3334
rect 26988 3058 27016 3606
rect 27264 3466 27292 4014
rect 27448 4010 27476 13194
rect 27632 12850 27660 13262
rect 27620 12844 27672 12850
rect 27620 12786 27672 12792
rect 27724 4146 27752 14758
rect 27816 14346 27844 14894
rect 27804 14340 27856 14346
rect 27804 14282 27856 14288
rect 27908 14006 27936 16662
rect 30012 16652 30064 16658
rect 30012 16594 30064 16600
rect 31300 16652 31352 16658
rect 31300 16594 31352 16600
rect 28816 16584 28868 16590
rect 28816 16526 28868 16532
rect 28828 16114 28856 16526
rect 29000 16176 29052 16182
rect 29000 16118 29052 16124
rect 28816 16108 28868 16114
rect 28816 16050 28868 16056
rect 28448 16040 28500 16046
rect 28448 15982 28500 15988
rect 28460 15706 28488 15982
rect 28540 15972 28592 15978
rect 28540 15914 28592 15920
rect 28552 15706 28580 15914
rect 28448 15700 28500 15706
rect 28448 15642 28500 15648
rect 28540 15700 28592 15706
rect 28540 15642 28592 15648
rect 27988 14340 28040 14346
rect 27988 14282 28040 14288
rect 27896 14000 27948 14006
rect 27896 13942 27948 13948
rect 28000 13938 28028 14282
rect 27988 13932 28040 13938
rect 27988 13874 28040 13880
rect 28000 13326 28028 13874
rect 29012 13870 29040 16118
rect 29092 14884 29144 14890
rect 29092 14826 29144 14832
rect 29000 13864 29052 13870
rect 29000 13806 29052 13812
rect 27988 13320 28040 13326
rect 27988 13262 28040 13268
rect 29104 7410 29132 14826
rect 30024 13938 30052 16594
rect 31312 14226 31340 16594
rect 31404 14414 31432 17206
rect 32416 17134 32444 17462
rect 32128 17128 32180 17134
rect 32128 17070 32180 17076
rect 32312 17128 32364 17134
rect 32312 17070 32364 17076
rect 32404 17128 32456 17134
rect 32404 17070 32456 17076
rect 32140 16114 32168 17070
rect 32324 16794 32352 17070
rect 32312 16788 32364 16794
rect 32312 16730 32364 16736
rect 32692 16658 32720 17870
rect 32811 17436 33119 17456
rect 32811 17434 32817 17436
rect 32873 17434 32897 17436
rect 32953 17434 32977 17436
rect 33033 17434 33057 17436
rect 33113 17434 33119 17436
rect 32873 17382 32875 17434
rect 33055 17382 33057 17434
rect 32811 17380 32817 17382
rect 32873 17380 32897 17382
rect 32953 17380 32977 17382
rect 33033 17380 33057 17382
rect 33113 17380 33119 17382
rect 32811 17360 33119 17380
rect 33520 17066 33548 19200
rect 34704 17128 34756 17134
rect 34704 17070 34756 17076
rect 34888 17128 34940 17134
rect 34888 17070 34940 17076
rect 33508 17060 33560 17066
rect 33508 17002 33560 17008
rect 32680 16652 32732 16658
rect 32680 16594 32732 16600
rect 32220 16584 32272 16590
rect 32220 16526 32272 16532
rect 32128 16108 32180 16114
rect 32128 16050 32180 16056
rect 32232 16046 32260 16526
rect 32404 16516 32456 16522
rect 32404 16458 32456 16464
rect 32416 16250 32444 16458
rect 33784 16448 33836 16454
rect 33784 16390 33836 16396
rect 32811 16348 33119 16368
rect 32811 16346 32817 16348
rect 32873 16346 32897 16348
rect 32953 16346 32977 16348
rect 33033 16346 33057 16348
rect 33113 16346 33119 16348
rect 32873 16294 32875 16346
rect 33055 16294 33057 16346
rect 32811 16292 32817 16294
rect 32873 16292 32897 16294
rect 32953 16292 32977 16294
rect 33033 16292 33057 16294
rect 33113 16292 33119 16294
rect 32811 16272 33119 16292
rect 32404 16244 32456 16250
rect 32404 16186 32456 16192
rect 33796 16114 33824 16390
rect 34716 16114 34744 17070
rect 34900 16250 34928 17070
rect 35452 16658 35480 19200
rect 35440 16652 35492 16658
rect 35440 16594 35492 16600
rect 35256 16516 35308 16522
rect 35256 16458 35308 16464
rect 35268 16250 35296 16458
rect 34888 16244 34940 16250
rect 34888 16186 34940 16192
rect 35256 16244 35308 16250
rect 35256 16186 35308 16192
rect 32680 16108 32732 16114
rect 32680 16050 32732 16056
rect 33784 16108 33836 16114
rect 33784 16050 33836 16056
rect 34704 16108 34756 16114
rect 34704 16050 34756 16056
rect 32220 16040 32272 16046
rect 32220 15982 32272 15988
rect 31668 15020 31720 15026
rect 31668 14962 31720 14968
rect 31484 14816 31536 14822
rect 31484 14758 31536 14764
rect 31392 14408 31444 14414
rect 31392 14350 31444 14356
rect 31312 14198 31432 14226
rect 30012 13932 30064 13938
rect 30012 13874 30064 13880
rect 31404 13870 31432 14198
rect 31392 13864 31444 13870
rect 31392 13806 31444 13812
rect 29736 7880 29788 7886
rect 29736 7822 29788 7828
rect 29748 7410 29776 7822
rect 29092 7404 29144 7410
rect 29092 7346 29144 7352
rect 29736 7404 29788 7410
rect 29736 7346 29788 7352
rect 27988 5636 28040 5642
rect 27988 5578 28040 5584
rect 28000 5234 28028 5578
rect 27988 5228 28040 5234
rect 27988 5170 28040 5176
rect 28080 5024 28132 5030
rect 28080 4966 28132 4972
rect 27896 4616 27948 4622
rect 27896 4558 27948 4564
rect 27908 4146 27936 4558
rect 28092 4214 28120 4966
rect 29000 4616 29052 4622
rect 29000 4558 29052 4564
rect 28080 4208 28132 4214
rect 28080 4150 28132 4156
rect 27712 4140 27764 4146
rect 27712 4082 27764 4088
rect 27896 4140 27948 4146
rect 27896 4082 27948 4088
rect 28356 4072 28408 4078
rect 28356 4014 28408 4020
rect 27436 4004 27488 4010
rect 27436 3946 27488 3952
rect 27712 3596 27764 3602
rect 27712 3538 27764 3544
rect 27068 3460 27120 3466
rect 27068 3402 27120 3408
rect 27252 3460 27304 3466
rect 27252 3402 27304 3408
rect 27080 3194 27108 3402
rect 27068 3188 27120 3194
rect 27068 3130 27120 3136
rect 26976 3052 27028 3058
rect 26976 2994 27028 3000
rect 26424 2848 26476 2854
rect 26424 2790 26476 2796
rect 26436 2514 26464 2790
rect 20812 2508 20864 2514
rect 20812 2450 20864 2456
rect 21088 2508 21140 2514
rect 21088 2450 21140 2456
rect 21272 2508 21324 2514
rect 21272 2450 21324 2456
rect 22468 2508 22520 2514
rect 23664 2508 23716 2514
rect 22520 2468 22600 2496
rect 22468 2450 22520 2456
rect 20824 1970 20852 2450
rect 20812 1964 20864 1970
rect 20812 1906 20864 1912
rect 22572 800 22600 2468
rect 23664 2450 23716 2456
rect 23848 2508 23900 2514
rect 23848 2450 23900 2456
rect 26240 2508 26292 2514
rect 26240 2450 26292 2456
rect 26424 2508 26476 2514
rect 26424 2450 26476 2456
rect 24584 2372 24636 2378
rect 24584 2314 24636 2320
rect 24596 2038 24624 2314
rect 24584 2032 24636 2038
rect 24584 1974 24636 1980
rect 27724 800 27752 3538
rect 28368 800 28396 4014
rect 28816 3528 28868 3534
rect 28816 3470 28868 3476
rect 28828 3058 28856 3470
rect 28816 3052 28868 3058
rect 28816 2994 28868 3000
rect 29012 2514 29040 4558
rect 29104 2990 29132 7346
rect 31404 3058 31432 13806
rect 31496 5234 31524 14758
rect 31680 14414 31708 14962
rect 32692 14958 32720 16050
rect 32811 15260 33119 15280
rect 32811 15258 32817 15260
rect 32873 15258 32897 15260
rect 32953 15258 32977 15260
rect 33033 15258 33057 15260
rect 33113 15258 33119 15260
rect 32873 15206 32875 15258
rect 33055 15206 33057 15258
rect 32811 15204 32817 15206
rect 32873 15204 32897 15206
rect 32953 15204 32977 15206
rect 33033 15204 33057 15206
rect 33113 15204 33119 15206
rect 32811 15184 33119 15204
rect 33796 15162 33824 16050
rect 35624 15904 35676 15910
rect 35624 15846 35676 15852
rect 35636 15570 35664 15846
rect 36096 15570 36124 19200
rect 37280 17128 37332 17134
rect 37280 17070 37332 17076
rect 37464 17128 37516 17134
rect 37464 17070 37516 17076
rect 36912 16584 36964 16590
rect 36912 16526 36964 16532
rect 36924 16114 36952 16526
rect 37292 16114 37320 17070
rect 37476 16794 37504 17070
rect 38028 16998 38056 19200
rect 39960 17270 39988 19200
rect 39948 17264 40000 17270
rect 39948 17206 40000 17212
rect 40604 17134 40632 19200
rect 39948 17128 40000 17134
rect 39948 17070 40000 17076
rect 40132 17128 40184 17134
rect 40132 17070 40184 17076
rect 40592 17128 40644 17134
rect 40592 17070 40644 17076
rect 38016 16992 38068 16998
rect 38016 16934 38068 16940
rect 39960 16794 39988 17070
rect 37464 16788 37516 16794
rect 37464 16730 37516 16736
rect 39948 16788 40000 16794
rect 39948 16730 40000 16736
rect 40144 16590 40172 17070
rect 40684 16992 40736 16998
rect 40684 16934 40736 16940
rect 40696 16726 40724 16934
rect 40776 16892 41084 16912
rect 40776 16890 40782 16892
rect 40838 16890 40862 16892
rect 40918 16890 40942 16892
rect 40998 16890 41022 16892
rect 41078 16890 41084 16892
rect 40838 16838 40840 16890
rect 41020 16838 41022 16890
rect 40776 16836 40782 16838
rect 40838 16836 40862 16838
rect 40918 16836 40942 16838
rect 40998 16836 41022 16838
rect 41078 16836 41084 16838
rect 40776 16816 41084 16836
rect 40684 16720 40736 16726
rect 40684 16662 40736 16668
rect 37372 16584 37424 16590
rect 37372 16526 37424 16532
rect 38936 16584 38988 16590
rect 38936 16526 38988 16532
rect 39856 16584 39908 16590
rect 39856 16526 39908 16532
rect 40132 16584 40184 16590
rect 40132 16526 40184 16532
rect 36912 16108 36964 16114
rect 36912 16050 36964 16056
rect 37280 16108 37332 16114
rect 37280 16050 37332 16056
rect 35624 15564 35676 15570
rect 35624 15506 35676 15512
rect 36084 15564 36136 15570
rect 36084 15506 36136 15512
rect 35900 15428 35952 15434
rect 35900 15370 35952 15376
rect 35912 15162 35940 15370
rect 33784 15156 33836 15162
rect 33784 15098 33836 15104
rect 35900 15156 35952 15162
rect 35900 15098 35952 15104
rect 35992 15020 36044 15026
rect 35992 14962 36044 14968
rect 32680 14952 32732 14958
rect 32680 14894 32732 14900
rect 31668 14408 31720 14414
rect 31668 14350 31720 14356
rect 32692 12714 32720 14894
rect 33232 14340 33284 14346
rect 33232 14282 33284 14288
rect 32811 14172 33119 14192
rect 32811 14170 32817 14172
rect 32873 14170 32897 14172
rect 32953 14170 32977 14172
rect 33033 14170 33057 14172
rect 33113 14170 33119 14172
rect 32873 14118 32875 14170
rect 33055 14118 33057 14170
rect 32811 14116 32817 14118
rect 32873 14116 32897 14118
rect 32953 14116 32977 14118
rect 33033 14116 33057 14118
rect 33113 14116 33119 14118
rect 32811 14096 33119 14116
rect 32811 13084 33119 13104
rect 32811 13082 32817 13084
rect 32873 13082 32897 13084
rect 32953 13082 32977 13084
rect 33033 13082 33057 13084
rect 33113 13082 33119 13084
rect 32873 13030 32875 13082
rect 33055 13030 33057 13082
rect 32811 13028 32817 13030
rect 32873 13028 32897 13030
rect 32953 13028 32977 13030
rect 33033 13028 33057 13030
rect 33113 13028 33119 13030
rect 32811 13008 33119 13028
rect 32680 12708 32732 12714
rect 32680 12650 32732 12656
rect 32692 5250 32720 12650
rect 32811 11996 33119 12016
rect 32811 11994 32817 11996
rect 32873 11994 32897 11996
rect 32953 11994 32977 11996
rect 33033 11994 33057 11996
rect 33113 11994 33119 11996
rect 32873 11942 32875 11994
rect 33055 11942 33057 11994
rect 32811 11940 32817 11942
rect 32873 11940 32897 11942
rect 32953 11940 32977 11942
rect 33033 11940 33057 11942
rect 33113 11940 33119 11942
rect 32811 11920 33119 11940
rect 32811 10908 33119 10928
rect 32811 10906 32817 10908
rect 32873 10906 32897 10908
rect 32953 10906 32977 10908
rect 33033 10906 33057 10908
rect 33113 10906 33119 10908
rect 32873 10854 32875 10906
rect 33055 10854 33057 10906
rect 32811 10852 32817 10854
rect 32873 10852 32897 10854
rect 32953 10852 32977 10854
rect 33033 10852 33057 10854
rect 33113 10852 33119 10854
rect 32811 10832 33119 10852
rect 32811 9820 33119 9840
rect 32811 9818 32817 9820
rect 32873 9818 32897 9820
rect 32953 9818 32977 9820
rect 33033 9818 33057 9820
rect 33113 9818 33119 9820
rect 32873 9766 32875 9818
rect 33055 9766 33057 9818
rect 32811 9764 32817 9766
rect 32873 9764 32897 9766
rect 32953 9764 32977 9766
rect 33033 9764 33057 9766
rect 33113 9764 33119 9766
rect 32811 9744 33119 9764
rect 32811 8732 33119 8752
rect 32811 8730 32817 8732
rect 32873 8730 32897 8732
rect 32953 8730 32977 8732
rect 33033 8730 33057 8732
rect 33113 8730 33119 8732
rect 32873 8678 32875 8730
rect 33055 8678 33057 8730
rect 32811 8676 32817 8678
rect 32873 8676 32897 8678
rect 32953 8676 32977 8678
rect 33033 8676 33057 8678
rect 33113 8676 33119 8678
rect 32811 8656 33119 8676
rect 33244 7886 33272 14282
rect 36004 14278 36032 14962
rect 35992 14272 36044 14278
rect 35992 14214 36044 14220
rect 34704 13932 34756 13938
rect 34704 13874 34756 13880
rect 33232 7880 33284 7886
rect 33232 7822 33284 7828
rect 33876 7744 33928 7750
rect 33876 7686 33928 7692
rect 32811 7644 33119 7664
rect 32811 7642 32817 7644
rect 32873 7642 32897 7644
rect 32953 7642 32977 7644
rect 33033 7642 33057 7644
rect 33113 7642 33119 7644
rect 32873 7590 32875 7642
rect 33055 7590 33057 7642
rect 32811 7588 32817 7590
rect 32873 7588 32897 7590
rect 32953 7588 32977 7590
rect 33033 7588 33057 7590
rect 33113 7588 33119 7590
rect 32811 7568 33119 7588
rect 33888 7478 33916 7686
rect 33876 7472 33928 7478
rect 33876 7414 33928 7420
rect 33692 7336 33744 7342
rect 33692 7278 33744 7284
rect 34612 7336 34664 7342
rect 34612 7278 34664 7284
rect 33704 7002 33732 7278
rect 33692 6996 33744 7002
rect 33692 6938 33744 6944
rect 32811 6556 33119 6576
rect 32811 6554 32817 6556
rect 32873 6554 32897 6556
rect 32953 6554 32977 6556
rect 33033 6554 33057 6556
rect 33113 6554 33119 6556
rect 32873 6502 32875 6554
rect 33055 6502 33057 6554
rect 32811 6500 32817 6502
rect 32873 6500 32897 6502
rect 32953 6500 32977 6502
rect 33033 6500 33057 6502
rect 33113 6500 33119 6502
rect 32811 6480 33119 6500
rect 32811 5468 33119 5488
rect 32811 5466 32817 5468
rect 32873 5466 32897 5468
rect 32953 5466 32977 5468
rect 33033 5466 33057 5468
rect 33113 5466 33119 5468
rect 32873 5414 32875 5466
rect 33055 5414 33057 5466
rect 32811 5412 32817 5414
rect 32873 5412 32897 5414
rect 32953 5412 32977 5414
rect 33033 5412 33057 5414
rect 33113 5412 33119 5414
rect 32811 5392 33119 5412
rect 31484 5228 31536 5234
rect 32692 5222 32812 5250
rect 31484 5170 31536 5176
rect 32680 5024 32732 5030
rect 32680 4966 32732 4972
rect 32036 4616 32088 4622
rect 32036 4558 32088 4564
rect 31576 3936 31628 3942
rect 31576 3878 31628 3884
rect 31588 3058 31616 3878
rect 32048 3602 32076 4558
rect 32692 4146 32720 4966
rect 32784 4622 32812 5222
rect 32772 4616 32824 4622
rect 32772 4558 32824 4564
rect 34520 4616 34572 4622
rect 34520 4558 34572 4564
rect 33140 4480 33192 4486
rect 33140 4422 33192 4428
rect 32811 4380 33119 4400
rect 32811 4378 32817 4380
rect 32873 4378 32897 4380
rect 32953 4378 32977 4380
rect 33033 4378 33057 4380
rect 33113 4378 33119 4380
rect 32873 4326 32875 4378
rect 33055 4326 33057 4378
rect 32811 4324 32817 4326
rect 32873 4324 32897 4326
rect 32953 4324 32977 4326
rect 33033 4324 33057 4326
rect 33113 4324 33119 4326
rect 32811 4304 33119 4324
rect 33152 4214 33180 4422
rect 33140 4208 33192 4214
rect 33140 4150 33192 4156
rect 32128 4140 32180 4146
rect 32128 4082 32180 4088
rect 32680 4140 32732 4146
rect 32680 4082 32732 4088
rect 32140 4010 32168 4082
rect 33508 4072 33560 4078
rect 33508 4014 33560 4020
rect 32128 4004 32180 4010
rect 32128 3946 32180 3952
rect 32140 3738 32168 3946
rect 32220 3936 32272 3942
rect 32220 3878 32272 3884
rect 32128 3732 32180 3738
rect 32128 3674 32180 3680
rect 32232 3602 32260 3878
rect 32036 3596 32088 3602
rect 32036 3538 32088 3544
rect 32220 3596 32272 3602
rect 32220 3538 32272 3544
rect 32680 3596 32732 3602
rect 32680 3538 32732 3544
rect 31944 3528 31996 3534
rect 31944 3470 31996 3476
rect 31392 3052 31444 3058
rect 31392 2994 31444 3000
rect 31576 3052 31628 3058
rect 31576 2994 31628 3000
rect 29092 2984 29144 2990
rect 29092 2926 29144 2932
rect 29644 2984 29696 2990
rect 29644 2926 29696 2932
rect 28816 2508 28868 2514
rect 28816 2450 28868 2456
rect 29000 2508 29052 2514
rect 29000 2450 29052 2456
rect 28828 1442 28856 2450
rect 29104 2446 29132 2926
rect 29092 2440 29144 2446
rect 29092 2382 29144 2388
rect 28828 1414 29040 1442
rect 29012 800 29040 1414
rect 29656 800 29684 2926
rect 31576 2576 31628 2582
rect 31576 2518 31628 2524
rect 31588 800 31616 2518
rect 31956 2514 31984 3470
rect 31944 2508 31996 2514
rect 31944 2450 31996 2456
rect 32220 1964 32272 1970
rect 32220 1906 32272 1912
rect 32232 800 32260 1906
rect 32692 1714 32720 3538
rect 32811 3292 33119 3312
rect 32811 3290 32817 3292
rect 32873 3290 32897 3292
rect 32953 3290 32977 3292
rect 33033 3290 33057 3292
rect 33113 3290 33119 3292
rect 32873 3238 32875 3290
rect 33055 3238 33057 3290
rect 32811 3236 32817 3238
rect 32873 3236 32897 3238
rect 32953 3236 32977 3238
rect 33033 3236 33057 3238
rect 33113 3236 33119 3238
rect 32811 3216 33119 3236
rect 32811 2204 33119 2224
rect 32811 2202 32817 2204
rect 32873 2202 32897 2204
rect 32953 2202 32977 2204
rect 33033 2202 33057 2204
rect 33113 2202 33119 2204
rect 32873 2150 32875 2202
rect 33055 2150 33057 2202
rect 32811 2148 32817 2150
rect 32873 2148 32897 2150
rect 32953 2148 32977 2150
rect 33033 2148 33057 2150
rect 33113 2148 33119 2150
rect 32811 2128 33119 2148
rect 32692 1686 32904 1714
rect 32876 800 32904 1686
rect 33520 800 33548 4014
rect 33968 2984 34020 2990
rect 33968 2926 34020 2932
rect 33980 1358 34008 2926
rect 34532 2514 34560 4558
rect 34520 2508 34572 2514
rect 34520 2450 34572 2456
rect 34624 2394 34652 7278
rect 34716 4622 34744 13874
rect 37384 13190 37412 16526
rect 38948 16114 38976 16526
rect 39120 16448 39172 16454
rect 39120 16390 39172 16396
rect 38936 16108 38988 16114
rect 38936 16050 38988 16056
rect 39132 16046 39160 16390
rect 39120 16040 39172 16046
rect 39120 15982 39172 15988
rect 39868 14482 39896 16526
rect 41236 15904 41288 15910
rect 41236 15846 41288 15852
rect 40776 15804 41084 15824
rect 40776 15802 40782 15804
rect 40838 15802 40862 15804
rect 40918 15802 40942 15804
rect 40998 15802 41022 15804
rect 41078 15802 41084 15804
rect 40838 15750 40840 15802
rect 41020 15750 41022 15802
rect 40776 15748 40782 15750
rect 40838 15748 40862 15750
rect 40918 15748 40942 15750
rect 40998 15748 41022 15750
rect 41078 15748 41084 15750
rect 40776 15728 41084 15748
rect 41248 15570 41276 15846
rect 41892 15570 41920 19200
rect 43180 17134 43208 19200
rect 42156 17128 42208 17134
rect 42156 17070 42208 17076
rect 42708 17128 42760 17134
rect 42708 17070 42760 17076
rect 43168 17128 43220 17134
rect 43168 17070 43220 17076
rect 42168 16794 42196 17070
rect 42156 16788 42208 16794
rect 42156 16730 42208 16736
rect 42432 16720 42484 16726
rect 42432 16662 42484 16668
rect 42444 16114 42472 16662
rect 42720 16250 42748 17070
rect 43824 16658 43852 19200
rect 46754 19136 46810 19145
rect 46754 19071 46810 19080
rect 45558 17776 45614 17785
rect 45558 17711 45614 17720
rect 44732 17128 44784 17134
rect 44732 17070 44784 17076
rect 45376 17128 45428 17134
rect 45376 17070 45428 17076
rect 43260 16652 43312 16658
rect 43260 16594 43312 16600
rect 43812 16652 43864 16658
rect 43812 16594 43864 16600
rect 43168 16448 43220 16454
rect 43168 16390 43220 16396
rect 42708 16244 42760 16250
rect 42708 16186 42760 16192
rect 43180 16114 43208 16390
rect 42432 16108 42484 16114
rect 42432 16050 42484 16056
rect 43168 16108 43220 16114
rect 43168 16050 43220 16056
rect 42800 16040 42852 16046
rect 42800 15982 42852 15988
rect 42812 15706 42840 15982
rect 42800 15700 42852 15706
rect 42800 15642 42852 15648
rect 41236 15564 41288 15570
rect 41236 15506 41288 15512
rect 41880 15564 41932 15570
rect 41880 15506 41932 15512
rect 40132 15496 40184 15502
rect 40132 15438 40184 15444
rect 39856 14476 39908 14482
rect 39856 14418 39908 14424
rect 36544 13184 36596 13190
rect 36544 13126 36596 13132
rect 37372 13184 37424 13190
rect 37372 13126 37424 13132
rect 34704 4616 34756 4622
rect 34704 4558 34756 4564
rect 35900 4616 35952 4622
rect 35900 4558 35952 4564
rect 34716 3534 34744 4558
rect 34796 4480 34848 4486
rect 34796 4422 34848 4428
rect 34704 3528 34756 3534
rect 34704 3470 34756 3476
rect 34808 2582 34836 4422
rect 34888 3936 34940 3942
rect 34888 3878 34940 3884
rect 34900 3058 34928 3878
rect 35912 3602 35940 4558
rect 36556 4146 36584 13126
rect 40040 10056 40092 10062
rect 40040 9998 40092 10004
rect 40052 9586 40080 9998
rect 40040 9580 40092 9586
rect 40040 9522 40092 9528
rect 37280 4616 37332 4622
rect 37280 4558 37332 4564
rect 37292 4146 37320 4558
rect 40144 4146 40172 15438
rect 40776 14716 41084 14736
rect 40776 14714 40782 14716
rect 40838 14714 40862 14716
rect 40918 14714 40942 14716
rect 40998 14714 41022 14716
rect 41078 14714 41084 14716
rect 40838 14662 40840 14714
rect 41020 14662 41022 14714
rect 40776 14660 40782 14662
rect 40838 14660 40862 14662
rect 40918 14660 40942 14662
rect 40998 14660 41022 14662
rect 41078 14660 41084 14662
rect 40776 14640 41084 14660
rect 40776 13628 41084 13648
rect 40776 13626 40782 13628
rect 40838 13626 40862 13628
rect 40918 13626 40942 13628
rect 40998 13626 41022 13628
rect 41078 13626 41084 13628
rect 40838 13574 40840 13626
rect 41020 13574 41022 13626
rect 40776 13572 40782 13574
rect 40838 13572 40862 13574
rect 40918 13572 40942 13574
rect 40998 13572 41022 13574
rect 41078 13572 41084 13574
rect 40776 13552 41084 13572
rect 42340 12776 42392 12782
rect 42340 12718 42392 12724
rect 40776 12540 41084 12560
rect 40776 12538 40782 12540
rect 40838 12538 40862 12540
rect 40918 12538 40942 12540
rect 40998 12538 41022 12540
rect 41078 12538 41084 12540
rect 40838 12486 40840 12538
rect 41020 12486 41022 12538
rect 40776 12484 40782 12486
rect 40838 12484 40862 12486
rect 40918 12484 40942 12486
rect 40998 12484 41022 12486
rect 41078 12484 41084 12486
rect 40776 12464 41084 12484
rect 40776 11452 41084 11472
rect 40776 11450 40782 11452
rect 40838 11450 40862 11452
rect 40918 11450 40942 11452
rect 40998 11450 41022 11452
rect 41078 11450 41084 11452
rect 40838 11398 40840 11450
rect 41020 11398 41022 11450
rect 40776 11396 40782 11398
rect 40838 11396 40862 11398
rect 40918 11396 40942 11398
rect 40998 11396 41022 11398
rect 41078 11396 41084 11398
rect 40776 11376 41084 11396
rect 40776 10364 41084 10384
rect 40776 10362 40782 10364
rect 40838 10362 40862 10364
rect 40918 10362 40942 10364
rect 40998 10362 41022 10364
rect 41078 10362 41084 10364
rect 40838 10310 40840 10362
rect 41020 10310 41022 10362
rect 40776 10308 40782 10310
rect 40838 10308 40862 10310
rect 40918 10308 40942 10310
rect 40998 10308 41022 10310
rect 41078 10308 41084 10310
rect 40776 10288 41084 10308
rect 40224 9512 40276 9518
rect 40224 9454 40276 9460
rect 40592 9512 40644 9518
rect 40592 9454 40644 9460
rect 40236 9178 40264 9454
rect 40224 9172 40276 9178
rect 40224 9114 40276 9120
rect 36544 4140 36596 4146
rect 36544 4082 36596 4088
rect 37280 4140 37332 4146
rect 37280 4082 37332 4088
rect 40132 4140 40184 4146
rect 40132 4082 40184 4088
rect 37556 4072 37608 4078
rect 37556 4014 37608 4020
rect 36084 3936 36136 3942
rect 36084 3878 36136 3884
rect 36096 3602 36124 3878
rect 35900 3596 35952 3602
rect 35900 3538 35952 3544
rect 36084 3596 36136 3602
rect 36084 3538 36136 3544
rect 36728 3596 36780 3602
rect 36728 3538 36780 3544
rect 35164 3460 35216 3466
rect 35164 3402 35216 3408
rect 35072 3392 35124 3398
rect 35072 3334 35124 3340
rect 35084 3126 35112 3334
rect 35176 3126 35204 3402
rect 35072 3120 35124 3126
rect 35072 3062 35124 3068
rect 35164 3120 35216 3126
rect 35164 3062 35216 3068
rect 34888 3052 34940 3058
rect 34888 2994 34940 3000
rect 36084 2984 36136 2990
rect 36084 2926 36136 2932
rect 34796 2576 34848 2582
rect 34796 2518 34848 2524
rect 34624 2366 34836 2394
rect 33968 1352 34020 1358
rect 33968 1294 34020 1300
rect 34808 800 34836 2366
rect 36096 800 36124 2926
rect 36740 800 36768 3538
rect 37280 3528 37332 3534
rect 37280 3470 37332 3476
rect 37292 2514 37320 3470
rect 37372 3052 37424 3058
rect 37372 2994 37424 3000
rect 37384 2650 37412 2994
rect 37464 2848 37516 2854
rect 37464 2790 37516 2796
rect 37372 2644 37424 2650
rect 37372 2586 37424 2592
rect 37476 2514 37504 2790
rect 37280 2508 37332 2514
rect 37280 2450 37332 2456
rect 37464 2508 37516 2514
rect 37464 2450 37516 2456
rect 37568 2122 37596 4014
rect 39948 3936 40000 3942
rect 39948 3878 40000 3884
rect 39120 3528 39172 3534
rect 39120 3470 39172 3476
rect 39856 3528 39908 3534
rect 39856 3470 39908 3476
rect 39132 3058 39160 3470
rect 39868 3194 39896 3470
rect 39856 3188 39908 3194
rect 39856 3130 39908 3136
rect 39120 3052 39172 3058
rect 39120 2994 39172 3000
rect 39960 2514 39988 3878
rect 40132 3392 40184 3398
rect 40132 3334 40184 3340
rect 40144 2514 40172 3334
rect 39948 2508 40000 2514
rect 39948 2450 40000 2456
rect 40132 2508 40184 2514
rect 40132 2450 40184 2456
rect 39304 2372 39356 2378
rect 39304 2314 39356 2320
rect 37384 2094 37596 2122
rect 37384 800 37412 2094
rect 39316 800 39344 2314
rect 40604 800 40632 9454
rect 40776 9276 41084 9296
rect 40776 9274 40782 9276
rect 40838 9274 40862 9276
rect 40918 9274 40942 9276
rect 40998 9274 41022 9276
rect 41078 9274 41084 9276
rect 40838 9222 40840 9274
rect 41020 9222 41022 9274
rect 40776 9220 40782 9222
rect 40838 9220 40862 9222
rect 40918 9220 40942 9222
rect 40998 9220 41022 9222
rect 41078 9220 41084 9222
rect 40776 9200 41084 9220
rect 40776 8188 41084 8208
rect 40776 8186 40782 8188
rect 40838 8186 40862 8188
rect 40918 8186 40942 8188
rect 40998 8186 41022 8188
rect 41078 8186 41084 8188
rect 40838 8134 40840 8186
rect 41020 8134 41022 8186
rect 40776 8132 40782 8134
rect 40838 8132 40862 8134
rect 40918 8132 40942 8134
rect 40998 8132 41022 8134
rect 41078 8132 41084 8134
rect 40776 8112 41084 8132
rect 40776 7100 41084 7120
rect 40776 7098 40782 7100
rect 40838 7098 40862 7100
rect 40918 7098 40942 7100
rect 40998 7098 41022 7100
rect 41078 7098 41084 7100
rect 40838 7046 40840 7098
rect 41020 7046 41022 7098
rect 40776 7044 40782 7046
rect 40838 7044 40862 7046
rect 40918 7044 40942 7046
rect 40998 7044 41022 7046
rect 41078 7044 41084 7046
rect 40776 7024 41084 7044
rect 40776 6012 41084 6032
rect 40776 6010 40782 6012
rect 40838 6010 40862 6012
rect 40918 6010 40942 6012
rect 40998 6010 41022 6012
rect 41078 6010 41084 6012
rect 40838 5958 40840 6010
rect 41020 5958 41022 6010
rect 40776 5956 40782 5958
rect 40838 5956 40862 5958
rect 40918 5956 40942 5958
rect 40998 5956 41022 5958
rect 41078 5956 41084 5958
rect 40776 5936 41084 5956
rect 40776 4924 41084 4944
rect 40776 4922 40782 4924
rect 40838 4922 40862 4924
rect 40918 4922 40942 4924
rect 40998 4922 41022 4924
rect 41078 4922 41084 4924
rect 40838 4870 40840 4922
rect 41020 4870 41022 4922
rect 40776 4868 40782 4870
rect 40838 4868 40862 4870
rect 40918 4868 40942 4870
rect 40998 4868 41022 4870
rect 41078 4868 41084 4870
rect 40776 4848 41084 4868
rect 42352 4622 42380 12718
rect 43180 6914 43208 16050
rect 43272 15706 43300 16594
rect 43444 16516 43496 16522
rect 43444 16458 43496 16464
rect 43456 16250 43484 16458
rect 43444 16244 43496 16250
rect 43444 16186 43496 16192
rect 44744 16114 44772 17070
rect 45388 16794 45416 17070
rect 45376 16788 45428 16794
rect 45376 16730 45428 16736
rect 45572 16182 45600 17711
rect 46570 17096 46626 17105
rect 46570 17031 46626 17040
rect 46584 16726 46612 17031
rect 46572 16720 46624 16726
rect 46572 16662 46624 16668
rect 45560 16176 45612 16182
rect 45560 16118 45612 16124
rect 44732 16108 44784 16114
rect 44732 16050 44784 16056
rect 45376 16040 45428 16046
rect 45376 15982 45428 15988
rect 45388 15706 45416 15982
rect 45560 15972 45612 15978
rect 45560 15914 45612 15920
rect 43260 15700 43312 15706
rect 43260 15642 43312 15648
rect 45376 15700 45428 15706
rect 45376 15642 45428 15648
rect 45572 15026 45600 15914
rect 46768 15570 46796 19071
rect 47044 17270 47072 19200
rect 47688 17898 47716 19200
rect 47596 17870 47716 17898
rect 47032 17264 47084 17270
rect 47032 17206 47084 17212
rect 47492 16992 47544 16998
rect 47492 16934 47544 16940
rect 47504 16574 47532 16934
rect 47320 16546 47532 16574
rect 46846 16416 46902 16425
rect 46846 16351 46902 16360
rect 46860 16046 46888 16351
rect 47320 16114 47348 16546
rect 47308 16108 47360 16114
rect 47308 16050 47360 16056
rect 46848 16040 46900 16046
rect 46848 15982 46900 15988
rect 46756 15564 46808 15570
rect 46756 15506 46808 15512
rect 45560 15020 45612 15026
rect 45560 14962 45612 14968
rect 46756 15020 46808 15026
rect 46756 14962 46808 14968
rect 46296 14816 46348 14822
rect 46296 14758 46348 14764
rect 46480 14816 46532 14822
rect 46480 14758 46532 14764
rect 46308 14482 46336 14758
rect 46492 14482 46520 14758
rect 46296 14476 46348 14482
rect 46296 14418 46348 14424
rect 46480 14476 46532 14482
rect 46480 14418 46532 14424
rect 45192 14408 45244 14414
rect 45192 14350 45244 14356
rect 45204 13938 45232 14350
rect 45192 13932 45244 13938
rect 45192 13874 45244 13880
rect 45192 12776 45244 12782
rect 45192 12718 45244 12724
rect 45204 12442 45232 12718
rect 45192 12436 45244 12442
rect 45192 12378 45244 12384
rect 46572 11688 46624 11694
rect 46572 11630 46624 11636
rect 46584 10810 46612 11630
rect 46768 11506 46796 14962
rect 46940 14952 46992 14958
rect 46940 14894 46992 14900
rect 46848 13864 46900 13870
rect 46848 13806 46900 13812
rect 46860 13705 46888 13806
rect 46846 13696 46902 13705
rect 46846 13631 46902 13640
rect 46952 13190 46980 14894
rect 47032 13932 47084 13938
rect 47032 13874 47084 13880
rect 46940 13184 46992 13190
rect 46940 13126 46992 13132
rect 46848 12776 46900 12782
rect 46848 12718 46900 12724
rect 46860 12345 46888 12718
rect 46846 12336 46902 12345
rect 46846 12271 46902 12280
rect 46848 11688 46900 11694
rect 46846 11656 46848 11665
rect 46900 11656 46902 11665
rect 46846 11591 46902 11600
rect 46768 11478 46888 11506
rect 46572 10804 46624 10810
rect 46572 10746 46624 10752
rect 46664 10668 46716 10674
rect 46664 10610 46716 10616
rect 46296 10464 46348 10470
rect 46296 10406 46348 10412
rect 46308 10130 46336 10406
rect 46296 10124 46348 10130
rect 46296 10066 46348 10072
rect 46676 8974 46704 10610
rect 46664 8968 46716 8974
rect 46664 8910 46716 8916
rect 46754 7576 46810 7585
rect 46754 7511 46810 7520
rect 46768 7342 46796 7511
rect 46756 7336 46808 7342
rect 46756 7278 46808 7284
rect 46860 6914 46888 11478
rect 47044 10674 47072 13874
rect 47032 10668 47084 10674
rect 47032 10610 47084 10616
rect 43180 6886 43300 6914
rect 43272 4622 43300 6886
rect 46768 6886 46888 6914
rect 46296 6792 46348 6798
rect 46296 6734 46348 6740
rect 45192 6248 45244 6254
rect 45192 6190 45244 6196
rect 45376 6248 45428 6254
rect 45376 6190 45428 6196
rect 45204 5914 45232 6190
rect 45192 5908 45244 5914
rect 45192 5850 45244 5856
rect 44456 5024 44508 5030
rect 44456 4966 44508 4972
rect 44732 5024 44784 5030
rect 44732 4966 44784 4972
rect 42340 4616 42392 4622
rect 42340 4558 42392 4564
rect 43260 4616 43312 4622
rect 43260 4558 43312 4564
rect 43720 4616 43772 4622
rect 43720 4558 43772 4564
rect 42616 4480 42668 4486
rect 42616 4422 42668 4428
rect 43168 4480 43220 4486
rect 43168 4422 43220 4428
rect 41880 4072 41932 4078
rect 41880 4014 41932 4020
rect 40776 3836 41084 3856
rect 40776 3834 40782 3836
rect 40838 3834 40862 3836
rect 40918 3834 40942 3836
rect 40998 3834 41022 3836
rect 41078 3834 41084 3836
rect 40838 3782 40840 3834
rect 41020 3782 41022 3834
rect 40776 3780 40782 3782
rect 40838 3780 40862 3782
rect 40918 3780 40942 3782
rect 40998 3780 41022 3782
rect 41078 3780 41084 3782
rect 40776 3760 41084 3780
rect 41696 3460 41748 3466
rect 41696 3402 41748 3408
rect 41708 3194 41736 3402
rect 41892 3398 41920 4014
rect 42432 3936 42484 3942
rect 42432 3878 42484 3884
rect 42444 3534 42472 3878
rect 42432 3528 42484 3534
rect 42432 3470 42484 3476
rect 42628 3466 42656 4422
rect 43180 4078 43208 4422
rect 43168 4072 43220 4078
rect 43168 4014 43220 4020
rect 43272 4010 43300 4558
rect 43260 4004 43312 4010
rect 43260 3946 43312 3952
rect 42616 3460 42668 3466
rect 42616 3402 42668 3408
rect 41880 3392 41932 3398
rect 41880 3334 41932 3340
rect 41696 3188 41748 3194
rect 41696 3130 41748 3136
rect 41892 3058 41920 3334
rect 41880 3052 41932 3058
rect 41880 2994 41932 3000
rect 43732 2990 43760 4558
rect 43812 3596 43864 3602
rect 43812 3538 43864 3544
rect 43720 2984 43772 2990
rect 43720 2926 43772 2932
rect 40776 2748 41084 2768
rect 40776 2746 40782 2748
rect 40838 2746 40862 2748
rect 40918 2746 40942 2748
rect 40998 2746 41022 2748
rect 41078 2746 41084 2748
rect 40838 2694 40840 2746
rect 41020 2694 41022 2746
rect 40776 2692 40782 2694
rect 40838 2692 40862 2694
rect 40918 2692 40942 2694
rect 40998 2692 41022 2694
rect 41078 2692 41084 2694
rect 40776 2672 41084 2692
rect 43824 2514 43852 3538
rect 43904 2984 43956 2990
rect 43904 2926 43956 2932
rect 43812 2508 43864 2514
rect 43812 2450 43864 2456
rect 43916 1578 43944 2926
rect 44364 2916 44416 2922
rect 44364 2858 44416 2864
rect 44180 2372 44232 2378
rect 44180 2314 44232 2320
rect 43824 1550 43944 1578
rect 43824 800 43852 1550
rect 44192 1086 44220 2314
rect 44376 1578 44404 2858
rect 44468 2446 44496 4966
rect 44744 4146 44772 4966
rect 45388 4826 45416 6190
rect 45652 5704 45704 5710
rect 45652 5646 45704 5652
rect 45664 5302 45692 5646
rect 45652 5296 45704 5302
rect 45652 5238 45704 5244
rect 45376 4820 45428 4826
rect 45376 4762 45428 4768
rect 46308 4690 46336 6734
rect 46572 6248 46624 6254
rect 46572 6190 46624 6196
rect 46388 6112 46440 6118
rect 46388 6054 46440 6060
rect 46400 5166 46428 6054
rect 46388 5160 46440 5166
rect 46388 5102 46440 5108
rect 46584 4865 46612 6190
rect 46664 5772 46716 5778
rect 46664 5714 46716 5720
rect 46676 5545 46704 5714
rect 46662 5536 46718 5545
rect 46662 5471 46718 5480
rect 46570 4856 46626 4865
rect 46570 4791 46626 4800
rect 46296 4684 46348 4690
rect 46296 4626 46348 4632
rect 45468 4616 45520 4622
rect 45468 4558 45520 4564
rect 44732 4140 44784 4146
rect 44732 4082 44784 4088
rect 45100 4072 45152 4078
rect 45100 4014 45152 4020
rect 45112 3738 45140 4014
rect 45100 3732 45152 3738
rect 45100 3674 45152 3680
rect 45100 3460 45152 3466
rect 45100 3402 45152 3408
rect 44456 2440 44508 2446
rect 44456 2382 44508 2388
rect 44376 1550 44496 1578
rect 44180 1080 44232 1086
rect 44180 1022 44232 1028
rect 44468 800 44496 1550
rect 45112 800 45140 3402
rect 45480 3058 45508 4558
rect 46664 4548 46716 4554
rect 46664 4490 46716 4496
rect 46480 3936 46532 3942
rect 46480 3878 46532 3884
rect 46492 3602 46520 3878
rect 46480 3596 46532 3602
rect 46480 3538 46532 3544
rect 46676 3194 46704 4490
rect 46664 3188 46716 3194
rect 46664 3130 46716 3136
rect 46768 3058 46796 6886
rect 47320 5234 47348 16050
rect 47492 12844 47544 12850
rect 47492 12786 47544 12792
rect 47504 12714 47532 12786
rect 47492 12708 47544 12714
rect 47492 12650 47544 12656
rect 47400 11756 47452 11762
rect 47400 11698 47452 11704
rect 47412 10674 47440 11698
rect 47400 10668 47452 10674
rect 47400 10610 47452 10616
rect 47308 5228 47360 5234
rect 47308 5170 47360 5176
rect 46848 5160 46900 5166
rect 46848 5102 46900 5108
rect 46860 4185 46888 5102
rect 46846 4176 46902 4185
rect 46846 4111 46902 4120
rect 47032 4072 47084 4078
rect 47032 4014 47084 4020
rect 46848 4004 46900 4010
rect 46848 3946 46900 3952
rect 46860 3505 46888 3946
rect 46846 3496 46902 3505
rect 46846 3431 46902 3440
rect 45468 3052 45520 3058
rect 45468 2994 45520 3000
rect 46756 3052 46808 3058
rect 46756 2994 46808 3000
rect 46572 2916 46624 2922
rect 46572 2858 46624 2864
rect 45560 2848 45612 2854
rect 45560 2790 45612 2796
rect 45572 2378 45600 2790
rect 45744 2576 45796 2582
rect 45744 2518 45796 2524
rect 45652 2440 45704 2446
rect 45652 2382 45704 2388
rect 45560 2372 45612 2378
rect 45560 2314 45612 2320
rect 45664 1465 45692 2382
rect 45650 1456 45706 1465
rect 45650 1391 45706 1400
rect 45756 800 45784 2518
rect 46584 2514 46612 2858
rect 46572 2508 46624 2514
rect 46572 2450 46624 2456
rect 46664 1352 46716 1358
rect 46664 1294 46716 1300
rect -10 0 102 800
rect 634 0 746 800
rect 1278 0 1390 800
rect 1922 0 2034 800
rect 2566 0 2678 800
rect 3210 0 3322 800
rect 3854 0 3966 800
rect 4498 0 4610 800
rect 5142 0 5254 800
rect 5786 0 5898 800
rect 6430 0 6542 800
rect 7074 0 7186 800
rect 7718 0 7830 800
rect 8362 0 8474 800
rect 9006 0 9118 800
rect 9650 0 9762 800
rect 10294 0 10406 800
rect 10938 0 11050 800
rect 11582 0 11694 800
rect 12226 0 12338 800
rect 12870 0 12982 800
rect 13514 0 13626 800
rect 14158 0 14270 800
rect 14802 0 14914 800
rect 15446 0 15558 800
rect 16090 0 16202 800
rect 16734 0 16846 800
rect 17378 0 17490 800
rect 18022 0 18134 800
rect 18666 0 18778 800
rect 19310 0 19422 800
rect 19954 0 20066 800
rect 20598 0 20710 800
rect 21242 0 21354 800
rect 21886 0 21998 800
rect 22530 0 22642 800
rect 23174 0 23286 800
rect 23818 0 23930 800
rect 24462 0 24574 800
rect 25106 0 25218 800
rect 25750 0 25862 800
rect 26394 0 26506 800
rect 27038 0 27150 800
rect 27682 0 27794 800
rect 28326 0 28438 800
rect 28970 0 29082 800
rect 29614 0 29726 800
rect 30258 0 30370 800
rect 30902 0 31014 800
rect 31546 0 31658 800
rect 32190 0 32302 800
rect 32834 0 32946 800
rect 33478 0 33590 800
rect 34766 0 34878 800
rect 35410 0 35522 800
rect 36054 0 36166 800
rect 36698 0 36810 800
rect 37342 0 37454 800
rect 37986 0 38098 800
rect 38630 0 38742 800
rect 39274 0 39386 800
rect 39918 0 40030 800
rect 40562 0 40674 800
rect 41206 0 41318 800
rect 41850 0 41962 800
rect 42494 0 42606 800
rect 43138 0 43250 800
rect 43782 0 43894 800
rect 44426 0 44538 800
rect 45070 0 45182 800
rect 45714 0 45826 800
rect 46358 0 46470 800
rect 46676 105 46704 1294
rect 46848 1080 46900 1086
rect 46848 1022 46900 1028
rect 46860 785 46888 1022
rect 47044 800 47072 4014
rect 47412 3058 47440 10610
rect 47504 6322 47532 12650
rect 47596 12306 47624 17870
rect 47768 16992 47820 16998
rect 47768 16934 47820 16940
rect 47676 16516 47728 16522
rect 47676 16458 47728 16464
rect 47688 16250 47716 16458
rect 47676 16244 47728 16250
rect 47676 16186 47728 16192
rect 47780 15570 47808 16934
rect 48332 16590 48360 19200
rect 48320 16584 48372 16590
rect 48320 16526 48372 16532
rect 47768 15564 47820 15570
rect 47768 15506 47820 15512
rect 47952 15428 48004 15434
rect 47952 15370 48004 15376
rect 47964 15162 47992 15370
rect 47952 15156 48004 15162
rect 47952 15098 48004 15104
rect 48134 15056 48190 15065
rect 48134 14991 48190 15000
rect 48148 14482 48176 14991
rect 48136 14476 48188 14482
rect 48136 14418 48188 14424
rect 48136 13252 48188 13258
rect 48136 13194 48188 13200
rect 48148 13025 48176 13194
rect 48134 13016 48190 13025
rect 48134 12951 48190 12960
rect 47584 12300 47636 12306
rect 47584 12242 47636 12248
rect 47676 12164 47728 12170
rect 47676 12106 47728 12112
rect 47688 11898 47716 12106
rect 47676 11892 47728 11898
rect 47676 11834 47728 11840
rect 47676 11076 47728 11082
rect 47676 11018 47728 11024
rect 48136 11076 48188 11082
rect 48136 11018 48188 11024
rect 47688 10810 47716 11018
rect 48148 10985 48176 11018
rect 48134 10976 48190 10985
rect 48134 10911 48190 10920
rect 47676 10804 47728 10810
rect 47676 10746 47728 10752
rect 48134 10296 48190 10305
rect 48134 10231 48190 10240
rect 48148 10130 48176 10231
rect 48136 10124 48188 10130
rect 48136 10066 48188 10072
rect 47676 9988 47728 9994
rect 47676 9930 47728 9936
rect 47688 9654 47716 9930
rect 47676 9648 47728 9654
rect 47676 9590 47728 9596
rect 47584 9580 47636 9586
rect 47584 9522 47636 9528
rect 47492 6316 47544 6322
rect 47492 6258 47544 6264
rect 47596 4146 47624 9522
rect 48136 6792 48188 6798
rect 48136 6734 48188 6740
rect 48148 5778 48176 6734
rect 48136 5772 48188 5778
rect 48136 5714 48188 5720
rect 47952 5636 48004 5642
rect 47952 5578 48004 5584
rect 47964 5370 47992 5578
rect 47952 5364 48004 5370
rect 47952 5306 48004 5312
rect 48320 4548 48372 4554
rect 48320 4490 48372 4496
rect 47584 4140 47636 4146
rect 47584 4082 47636 4088
rect 47596 3670 47624 4082
rect 47584 3664 47636 3670
rect 47584 3606 47636 3612
rect 48136 3460 48188 3466
rect 48136 3402 48188 3408
rect 47400 3052 47452 3058
rect 47400 2994 47452 3000
rect 47676 2848 47728 2854
rect 48148 2825 48176 3402
rect 47676 2790 47728 2796
rect 48134 2816 48190 2825
rect 47688 2514 47716 2790
rect 48134 2751 48190 2760
rect 47676 2508 47728 2514
rect 47676 2450 47728 2456
rect 47676 2304 47728 2310
rect 47676 2246 47728 2252
rect 47688 800 47716 2246
rect 48332 800 48360 4490
rect 49608 2916 49660 2922
rect 49608 2858 49660 2864
rect 49620 800 49648 2858
rect 46846 776 46902 785
rect 46846 711 46902 720
rect 46662 96 46718 105
rect 46662 31 46718 40
rect 47002 0 47114 800
rect 47646 0 47758 800
rect 48290 0 48402 800
rect 48934 0 49046 800
rect 49578 0 49690 800
<< via2 >>
rect 1398 17720 1454 17776
rect 4066 17040 4122 17096
rect 2778 15680 2834 15736
rect 2778 14320 2834 14376
rect 2778 12960 2834 13016
rect 4066 12300 4122 12336
rect 4066 12280 4068 12300
rect 4068 12280 4120 12300
rect 4120 12280 4122 12300
rect 2778 10920 2834 10976
rect 3422 10240 3478 10296
rect 2778 8200 2834 8256
rect 3422 7520 3478 7576
rect 2778 6840 2834 6896
rect 1398 4800 1454 4856
rect 2778 5480 2834 5536
rect 2778 4120 2834 4176
rect 3974 3440 4030 3496
rect 8921 16890 8977 16892
rect 9001 16890 9057 16892
rect 9081 16890 9137 16892
rect 9161 16890 9217 16892
rect 8921 16838 8967 16890
rect 8967 16838 8977 16890
rect 9001 16838 9031 16890
rect 9031 16838 9043 16890
rect 9043 16838 9057 16890
rect 9081 16838 9095 16890
rect 9095 16838 9107 16890
rect 9107 16838 9137 16890
rect 9161 16838 9171 16890
rect 9171 16838 9217 16890
rect 8921 16836 8977 16838
rect 9001 16836 9057 16838
rect 9081 16836 9137 16838
rect 9161 16836 9217 16838
rect 8921 15802 8977 15804
rect 9001 15802 9057 15804
rect 9081 15802 9137 15804
rect 9161 15802 9217 15804
rect 8921 15750 8967 15802
rect 8967 15750 8977 15802
rect 9001 15750 9031 15802
rect 9031 15750 9043 15802
rect 9043 15750 9057 15802
rect 9081 15750 9095 15802
rect 9095 15750 9107 15802
rect 9107 15750 9137 15802
rect 9161 15750 9171 15802
rect 9171 15750 9217 15802
rect 8921 15748 8977 15750
rect 9001 15748 9057 15750
rect 9081 15748 9137 15750
rect 9161 15748 9217 15750
rect 8921 14714 8977 14716
rect 9001 14714 9057 14716
rect 9081 14714 9137 14716
rect 9161 14714 9217 14716
rect 8921 14662 8967 14714
rect 8967 14662 8977 14714
rect 9001 14662 9031 14714
rect 9031 14662 9043 14714
rect 9043 14662 9057 14714
rect 9081 14662 9095 14714
rect 9095 14662 9107 14714
rect 9107 14662 9137 14714
rect 9161 14662 9171 14714
rect 9171 14662 9217 14714
rect 8921 14660 8977 14662
rect 9001 14660 9057 14662
rect 9081 14660 9137 14662
rect 9161 14660 9217 14662
rect 8921 13626 8977 13628
rect 9001 13626 9057 13628
rect 9081 13626 9137 13628
rect 9161 13626 9217 13628
rect 8921 13574 8967 13626
rect 8967 13574 8977 13626
rect 9001 13574 9031 13626
rect 9031 13574 9043 13626
rect 9043 13574 9057 13626
rect 9081 13574 9095 13626
rect 9095 13574 9107 13626
rect 9107 13574 9137 13626
rect 9161 13574 9171 13626
rect 9171 13574 9217 13626
rect 8921 13572 8977 13574
rect 9001 13572 9057 13574
rect 9081 13572 9137 13574
rect 9161 13572 9217 13574
rect 8921 12538 8977 12540
rect 9001 12538 9057 12540
rect 9081 12538 9137 12540
rect 9161 12538 9217 12540
rect 8921 12486 8967 12538
rect 8967 12486 8977 12538
rect 9001 12486 9031 12538
rect 9031 12486 9043 12538
rect 9043 12486 9057 12538
rect 9081 12486 9095 12538
rect 9095 12486 9107 12538
rect 9107 12486 9137 12538
rect 9161 12486 9171 12538
rect 9171 12486 9217 12538
rect 8921 12484 8977 12486
rect 9001 12484 9057 12486
rect 9081 12484 9137 12486
rect 9161 12484 9217 12486
rect 2870 2760 2926 2816
rect 3422 2080 3478 2136
rect 3514 1400 3570 1456
rect 8921 11450 8977 11452
rect 9001 11450 9057 11452
rect 9081 11450 9137 11452
rect 9161 11450 9217 11452
rect 8921 11398 8967 11450
rect 8967 11398 8977 11450
rect 9001 11398 9031 11450
rect 9031 11398 9043 11450
rect 9043 11398 9057 11450
rect 9081 11398 9095 11450
rect 9095 11398 9107 11450
rect 9107 11398 9137 11450
rect 9161 11398 9171 11450
rect 9171 11398 9217 11450
rect 8921 11396 8977 11398
rect 9001 11396 9057 11398
rect 9081 11396 9137 11398
rect 9161 11396 9217 11398
rect 8921 10362 8977 10364
rect 9001 10362 9057 10364
rect 9081 10362 9137 10364
rect 9161 10362 9217 10364
rect 8921 10310 8967 10362
rect 8967 10310 8977 10362
rect 9001 10310 9031 10362
rect 9031 10310 9043 10362
rect 9043 10310 9057 10362
rect 9081 10310 9095 10362
rect 9095 10310 9107 10362
rect 9107 10310 9137 10362
rect 9161 10310 9171 10362
rect 9171 10310 9217 10362
rect 8921 10308 8977 10310
rect 9001 10308 9057 10310
rect 9081 10308 9137 10310
rect 9161 10308 9217 10310
rect 8921 9274 8977 9276
rect 9001 9274 9057 9276
rect 9081 9274 9137 9276
rect 9161 9274 9217 9276
rect 8921 9222 8967 9274
rect 8967 9222 8977 9274
rect 9001 9222 9031 9274
rect 9031 9222 9043 9274
rect 9043 9222 9057 9274
rect 9081 9222 9095 9274
rect 9095 9222 9107 9274
rect 9107 9222 9137 9274
rect 9161 9222 9171 9274
rect 9171 9222 9217 9274
rect 8921 9220 8977 9222
rect 9001 9220 9057 9222
rect 9081 9220 9137 9222
rect 9161 9220 9217 9222
rect 8921 8186 8977 8188
rect 9001 8186 9057 8188
rect 9081 8186 9137 8188
rect 9161 8186 9217 8188
rect 8921 8134 8967 8186
rect 8967 8134 8977 8186
rect 9001 8134 9031 8186
rect 9031 8134 9043 8186
rect 9043 8134 9057 8186
rect 9081 8134 9095 8186
rect 9095 8134 9107 8186
rect 9107 8134 9137 8186
rect 9161 8134 9171 8186
rect 9171 8134 9217 8186
rect 8921 8132 8977 8134
rect 9001 8132 9057 8134
rect 9081 8132 9137 8134
rect 9161 8132 9217 8134
rect 8921 7098 8977 7100
rect 9001 7098 9057 7100
rect 9081 7098 9137 7100
rect 9161 7098 9217 7100
rect 8921 7046 8967 7098
rect 8967 7046 8977 7098
rect 9001 7046 9031 7098
rect 9031 7046 9043 7098
rect 9043 7046 9057 7098
rect 9081 7046 9095 7098
rect 9095 7046 9107 7098
rect 9107 7046 9137 7098
rect 9161 7046 9171 7098
rect 9171 7046 9217 7098
rect 8921 7044 8977 7046
rect 9001 7044 9057 7046
rect 9081 7044 9137 7046
rect 9161 7044 9217 7046
rect 8921 6010 8977 6012
rect 9001 6010 9057 6012
rect 9081 6010 9137 6012
rect 9161 6010 9217 6012
rect 8921 5958 8967 6010
rect 8967 5958 8977 6010
rect 9001 5958 9031 6010
rect 9031 5958 9043 6010
rect 9043 5958 9057 6010
rect 9081 5958 9095 6010
rect 9095 5958 9107 6010
rect 9107 5958 9137 6010
rect 9161 5958 9171 6010
rect 9171 5958 9217 6010
rect 8921 5956 8977 5958
rect 9001 5956 9057 5958
rect 9081 5956 9137 5958
rect 9161 5956 9217 5958
rect 8921 4922 8977 4924
rect 9001 4922 9057 4924
rect 9081 4922 9137 4924
rect 9161 4922 9217 4924
rect 8921 4870 8967 4922
rect 8967 4870 8977 4922
rect 9001 4870 9031 4922
rect 9031 4870 9043 4922
rect 9043 4870 9057 4922
rect 9081 4870 9095 4922
rect 9095 4870 9107 4922
rect 9107 4870 9137 4922
rect 9161 4870 9171 4922
rect 9171 4870 9217 4922
rect 8921 4868 8977 4870
rect 9001 4868 9057 4870
rect 9081 4868 9137 4870
rect 9161 4868 9217 4870
rect 8921 3834 8977 3836
rect 9001 3834 9057 3836
rect 9081 3834 9137 3836
rect 9161 3834 9217 3836
rect 8921 3782 8967 3834
rect 8967 3782 8977 3834
rect 9001 3782 9031 3834
rect 9031 3782 9043 3834
rect 9043 3782 9057 3834
rect 9081 3782 9095 3834
rect 9095 3782 9107 3834
rect 9107 3782 9137 3834
rect 9161 3782 9171 3834
rect 9171 3782 9217 3834
rect 8921 3780 8977 3782
rect 9001 3780 9057 3782
rect 9081 3780 9137 3782
rect 9161 3780 9217 3782
rect 8921 2746 8977 2748
rect 9001 2746 9057 2748
rect 9081 2746 9137 2748
rect 9161 2746 9217 2748
rect 8921 2694 8967 2746
rect 8967 2694 8977 2746
rect 9001 2694 9031 2746
rect 9031 2694 9043 2746
rect 9043 2694 9057 2746
rect 9081 2694 9095 2746
rect 9095 2694 9107 2746
rect 9107 2694 9137 2746
rect 9161 2694 9171 2746
rect 9171 2694 9217 2746
rect 8921 2692 8977 2694
rect 9001 2692 9057 2694
rect 9081 2692 9137 2694
rect 9161 2692 9217 2694
rect 16886 17434 16942 17436
rect 16966 17434 17022 17436
rect 17046 17434 17102 17436
rect 17126 17434 17182 17436
rect 16886 17382 16932 17434
rect 16932 17382 16942 17434
rect 16966 17382 16996 17434
rect 16996 17382 17008 17434
rect 17008 17382 17022 17434
rect 17046 17382 17060 17434
rect 17060 17382 17072 17434
rect 17072 17382 17102 17434
rect 17126 17382 17136 17434
rect 17136 17382 17182 17434
rect 16886 17380 16942 17382
rect 16966 17380 17022 17382
rect 17046 17380 17102 17382
rect 17126 17380 17182 17382
rect 16886 16346 16942 16348
rect 16966 16346 17022 16348
rect 17046 16346 17102 16348
rect 17126 16346 17182 16348
rect 16886 16294 16932 16346
rect 16932 16294 16942 16346
rect 16966 16294 16996 16346
rect 16996 16294 17008 16346
rect 17008 16294 17022 16346
rect 17046 16294 17060 16346
rect 17060 16294 17072 16346
rect 17072 16294 17102 16346
rect 17126 16294 17136 16346
rect 17136 16294 17182 16346
rect 16886 16292 16942 16294
rect 16966 16292 17022 16294
rect 17046 16292 17102 16294
rect 17126 16292 17182 16294
rect 16886 15258 16942 15260
rect 16966 15258 17022 15260
rect 17046 15258 17102 15260
rect 17126 15258 17182 15260
rect 16886 15206 16932 15258
rect 16932 15206 16942 15258
rect 16966 15206 16996 15258
rect 16996 15206 17008 15258
rect 17008 15206 17022 15258
rect 17046 15206 17060 15258
rect 17060 15206 17072 15258
rect 17072 15206 17102 15258
rect 17126 15206 17136 15258
rect 17136 15206 17182 15258
rect 16886 15204 16942 15206
rect 16966 15204 17022 15206
rect 17046 15204 17102 15206
rect 17126 15204 17182 15206
rect 16886 14170 16942 14172
rect 16966 14170 17022 14172
rect 17046 14170 17102 14172
rect 17126 14170 17182 14172
rect 16886 14118 16932 14170
rect 16932 14118 16942 14170
rect 16966 14118 16996 14170
rect 16996 14118 17008 14170
rect 17008 14118 17022 14170
rect 17046 14118 17060 14170
rect 17060 14118 17072 14170
rect 17072 14118 17102 14170
rect 17126 14118 17136 14170
rect 17136 14118 17182 14170
rect 16886 14116 16942 14118
rect 16966 14116 17022 14118
rect 17046 14116 17102 14118
rect 17126 14116 17182 14118
rect 16886 13082 16942 13084
rect 16966 13082 17022 13084
rect 17046 13082 17102 13084
rect 17126 13082 17182 13084
rect 16886 13030 16932 13082
rect 16932 13030 16942 13082
rect 16966 13030 16996 13082
rect 16996 13030 17008 13082
rect 17008 13030 17022 13082
rect 17046 13030 17060 13082
rect 17060 13030 17072 13082
rect 17072 13030 17102 13082
rect 17126 13030 17136 13082
rect 17136 13030 17182 13082
rect 16886 13028 16942 13030
rect 16966 13028 17022 13030
rect 17046 13028 17102 13030
rect 17126 13028 17182 13030
rect 16886 11994 16942 11996
rect 16966 11994 17022 11996
rect 17046 11994 17102 11996
rect 17126 11994 17182 11996
rect 16886 11942 16932 11994
rect 16932 11942 16942 11994
rect 16966 11942 16996 11994
rect 16996 11942 17008 11994
rect 17008 11942 17022 11994
rect 17046 11942 17060 11994
rect 17060 11942 17072 11994
rect 17072 11942 17102 11994
rect 17126 11942 17136 11994
rect 17136 11942 17182 11994
rect 16886 11940 16942 11942
rect 16966 11940 17022 11942
rect 17046 11940 17102 11942
rect 17126 11940 17182 11942
rect 16886 10906 16942 10908
rect 16966 10906 17022 10908
rect 17046 10906 17102 10908
rect 17126 10906 17182 10908
rect 16886 10854 16932 10906
rect 16932 10854 16942 10906
rect 16966 10854 16996 10906
rect 16996 10854 17008 10906
rect 17008 10854 17022 10906
rect 17046 10854 17060 10906
rect 17060 10854 17072 10906
rect 17072 10854 17102 10906
rect 17126 10854 17136 10906
rect 17136 10854 17182 10906
rect 16886 10852 16942 10854
rect 16966 10852 17022 10854
rect 17046 10852 17102 10854
rect 17126 10852 17182 10854
rect 16886 9818 16942 9820
rect 16966 9818 17022 9820
rect 17046 9818 17102 9820
rect 17126 9818 17182 9820
rect 16886 9766 16932 9818
rect 16932 9766 16942 9818
rect 16966 9766 16996 9818
rect 16996 9766 17008 9818
rect 17008 9766 17022 9818
rect 17046 9766 17060 9818
rect 17060 9766 17072 9818
rect 17072 9766 17102 9818
rect 17126 9766 17136 9818
rect 17136 9766 17182 9818
rect 16886 9764 16942 9766
rect 16966 9764 17022 9766
rect 17046 9764 17102 9766
rect 17126 9764 17182 9766
rect 16886 8730 16942 8732
rect 16966 8730 17022 8732
rect 17046 8730 17102 8732
rect 17126 8730 17182 8732
rect 16886 8678 16932 8730
rect 16932 8678 16942 8730
rect 16966 8678 16996 8730
rect 16996 8678 17008 8730
rect 17008 8678 17022 8730
rect 17046 8678 17060 8730
rect 17060 8678 17072 8730
rect 17072 8678 17102 8730
rect 17126 8678 17136 8730
rect 17136 8678 17182 8730
rect 16886 8676 16942 8678
rect 16966 8676 17022 8678
rect 17046 8676 17102 8678
rect 17126 8676 17182 8678
rect 16886 7642 16942 7644
rect 16966 7642 17022 7644
rect 17046 7642 17102 7644
rect 17126 7642 17182 7644
rect 16886 7590 16932 7642
rect 16932 7590 16942 7642
rect 16966 7590 16996 7642
rect 16996 7590 17008 7642
rect 17008 7590 17022 7642
rect 17046 7590 17060 7642
rect 17060 7590 17072 7642
rect 17072 7590 17102 7642
rect 17126 7590 17136 7642
rect 17136 7590 17182 7642
rect 16886 7588 16942 7590
rect 16966 7588 17022 7590
rect 17046 7588 17102 7590
rect 17126 7588 17182 7590
rect 16886 6554 16942 6556
rect 16966 6554 17022 6556
rect 17046 6554 17102 6556
rect 17126 6554 17182 6556
rect 16886 6502 16932 6554
rect 16932 6502 16942 6554
rect 16966 6502 16996 6554
rect 16996 6502 17008 6554
rect 17008 6502 17022 6554
rect 17046 6502 17060 6554
rect 17060 6502 17072 6554
rect 17072 6502 17102 6554
rect 17126 6502 17136 6554
rect 17136 6502 17182 6554
rect 16886 6500 16942 6502
rect 16966 6500 17022 6502
rect 17046 6500 17102 6502
rect 17126 6500 17182 6502
rect 16886 5466 16942 5468
rect 16966 5466 17022 5468
rect 17046 5466 17102 5468
rect 17126 5466 17182 5468
rect 16886 5414 16932 5466
rect 16932 5414 16942 5466
rect 16966 5414 16996 5466
rect 16996 5414 17008 5466
rect 17008 5414 17022 5466
rect 17046 5414 17060 5466
rect 17060 5414 17072 5466
rect 17072 5414 17102 5466
rect 17126 5414 17136 5466
rect 17136 5414 17182 5466
rect 16886 5412 16942 5414
rect 16966 5412 17022 5414
rect 17046 5412 17102 5414
rect 17126 5412 17182 5414
rect 16886 4378 16942 4380
rect 16966 4378 17022 4380
rect 17046 4378 17102 4380
rect 17126 4378 17182 4380
rect 16886 4326 16932 4378
rect 16932 4326 16942 4378
rect 16966 4326 16996 4378
rect 16996 4326 17008 4378
rect 17008 4326 17022 4378
rect 17046 4326 17060 4378
rect 17060 4326 17072 4378
rect 17072 4326 17102 4378
rect 17126 4326 17136 4378
rect 17136 4326 17182 4378
rect 16886 4324 16942 4326
rect 16966 4324 17022 4326
rect 17046 4324 17102 4326
rect 17126 4324 17182 4326
rect 16886 3290 16942 3292
rect 16966 3290 17022 3292
rect 17046 3290 17102 3292
rect 17126 3290 17182 3292
rect 16886 3238 16932 3290
rect 16932 3238 16942 3290
rect 16966 3238 16996 3290
rect 16996 3238 17008 3290
rect 17008 3238 17022 3290
rect 17046 3238 17060 3290
rect 17060 3238 17072 3290
rect 17072 3238 17102 3290
rect 17126 3238 17136 3290
rect 17136 3238 17182 3290
rect 16886 3236 16942 3238
rect 16966 3236 17022 3238
rect 17046 3236 17102 3238
rect 17126 3236 17182 3238
rect 16886 2202 16942 2204
rect 16966 2202 17022 2204
rect 17046 2202 17102 2204
rect 17126 2202 17182 2204
rect 16886 2150 16932 2202
rect 16932 2150 16942 2202
rect 16966 2150 16996 2202
rect 16996 2150 17008 2202
rect 17008 2150 17022 2202
rect 17046 2150 17060 2202
rect 17060 2150 17072 2202
rect 17072 2150 17102 2202
rect 17126 2150 17136 2202
rect 17136 2150 17182 2202
rect 16886 2148 16942 2150
rect 16966 2148 17022 2150
rect 17046 2148 17102 2150
rect 17126 2148 17182 2150
rect 24852 16890 24908 16892
rect 24932 16890 24988 16892
rect 25012 16890 25068 16892
rect 25092 16890 25148 16892
rect 24852 16838 24898 16890
rect 24898 16838 24908 16890
rect 24932 16838 24962 16890
rect 24962 16838 24974 16890
rect 24974 16838 24988 16890
rect 25012 16838 25026 16890
rect 25026 16838 25038 16890
rect 25038 16838 25068 16890
rect 25092 16838 25102 16890
rect 25102 16838 25148 16890
rect 24852 16836 24908 16838
rect 24932 16836 24988 16838
rect 25012 16836 25068 16838
rect 25092 16836 25148 16838
rect 24852 15802 24908 15804
rect 24932 15802 24988 15804
rect 25012 15802 25068 15804
rect 25092 15802 25148 15804
rect 24852 15750 24898 15802
rect 24898 15750 24908 15802
rect 24932 15750 24962 15802
rect 24962 15750 24974 15802
rect 24974 15750 24988 15802
rect 25012 15750 25026 15802
rect 25026 15750 25038 15802
rect 25038 15750 25068 15802
rect 25092 15750 25102 15802
rect 25102 15750 25148 15802
rect 24852 15748 24908 15750
rect 24932 15748 24988 15750
rect 25012 15748 25068 15750
rect 25092 15748 25148 15750
rect 24852 14714 24908 14716
rect 24932 14714 24988 14716
rect 25012 14714 25068 14716
rect 25092 14714 25148 14716
rect 24852 14662 24898 14714
rect 24898 14662 24908 14714
rect 24932 14662 24962 14714
rect 24962 14662 24974 14714
rect 24974 14662 24988 14714
rect 25012 14662 25026 14714
rect 25026 14662 25038 14714
rect 25038 14662 25068 14714
rect 25092 14662 25102 14714
rect 25102 14662 25148 14714
rect 24852 14660 24908 14662
rect 24932 14660 24988 14662
rect 25012 14660 25068 14662
rect 25092 14660 25148 14662
rect 24852 13626 24908 13628
rect 24932 13626 24988 13628
rect 25012 13626 25068 13628
rect 25092 13626 25148 13628
rect 24852 13574 24898 13626
rect 24898 13574 24908 13626
rect 24932 13574 24962 13626
rect 24962 13574 24974 13626
rect 24974 13574 24988 13626
rect 25012 13574 25026 13626
rect 25026 13574 25038 13626
rect 25038 13574 25068 13626
rect 25092 13574 25102 13626
rect 25102 13574 25148 13626
rect 24852 13572 24908 13574
rect 24932 13572 24988 13574
rect 25012 13572 25068 13574
rect 25092 13572 25148 13574
rect 24852 12538 24908 12540
rect 24932 12538 24988 12540
rect 25012 12538 25068 12540
rect 25092 12538 25148 12540
rect 24852 12486 24898 12538
rect 24898 12486 24908 12538
rect 24932 12486 24962 12538
rect 24962 12486 24974 12538
rect 24974 12486 24988 12538
rect 25012 12486 25026 12538
rect 25026 12486 25038 12538
rect 25038 12486 25068 12538
rect 25092 12486 25102 12538
rect 25102 12486 25148 12538
rect 24852 12484 24908 12486
rect 24932 12484 24988 12486
rect 25012 12484 25068 12486
rect 25092 12484 25148 12486
rect 24852 11450 24908 11452
rect 24932 11450 24988 11452
rect 25012 11450 25068 11452
rect 25092 11450 25148 11452
rect 24852 11398 24898 11450
rect 24898 11398 24908 11450
rect 24932 11398 24962 11450
rect 24962 11398 24974 11450
rect 24974 11398 24988 11450
rect 25012 11398 25026 11450
rect 25026 11398 25038 11450
rect 25038 11398 25068 11450
rect 25092 11398 25102 11450
rect 25102 11398 25148 11450
rect 24852 11396 24908 11398
rect 24932 11396 24988 11398
rect 25012 11396 25068 11398
rect 25092 11396 25148 11398
rect 24852 10362 24908 10364
rect 24932 10362 24988 10364
rect 25012 10362 25068 10364
rect 25092 10362 25148 10364
rect 24852 10310 24898 10362
rect 24898 10310 24908 10362
rect 24932 10310 24962 10362
rect 24962 10310 24974 10362
rect 24974 10310 24988 10362
rect 25012 10310 25026 10362
rect 25026 10310 25038 10362
rect 25038 10310 25068 10362
rect 25092 10310 25102 10362
rect 25102 10310 25148 10362
rect 24852 10308 24908 10310
rect 24932 10308 24988 10310
rect 25012 10308 25068 10310
rect 25092 10308 25148 10310
rect 24852 9274 24908 9276
rect 24932 9274 24988 9276
rect 25012 9274 25068 9276
rect 25092 9274 25148 9276
rect 24852 9222 24898 9274
rect 24898 9222 24908 9274
rect 24932 9222 24962 9274
rect 24962 9222 24974 9274
rect 24974 9222 24988 9274
rect 25012 9222 25026 9274
rect 25026 9222 25038 9274
rect 25038 9222 25068 9274
rect 25092 9222 25102 9274
rect 25102 9222 25148 9274
rect 24852 9220 24908 9222
rect 24932 9220 24988 9222
rect 25012 9220 25068 9222
rect 25092 9220 25148 9222
rect 24852 8186 24908 8188
rect 24932 8186 24988 8188
rect 25012 8186 25068 8188
rect 25092 8186 25148 8188
rect 24852 8134 24898 8186
rect 24898 8134 24908 8186
rect 24932 8134 24962 8186
rect 24962 8134 24974 8186
rect 24974 8134 24988 8186
rect 25012 8134 25026 8186
rect 25026 8134 25038 8186
rect 25038 8134 25068 8186
rect 25092 8134 25102 8186
rect 25102 8134 25148 8186
rect 24852 8132 24908 8134
rect 24932 8132 24988 8134
rect 25012 8132 25068 8134
rect 25092 8132 25148 8134
rect 24852 7098 24908 7100
rect 24932 7098 24988 7100
rect 25012 7098 25068 7100
rect 25092 7098 25148 7100
rect 24852 7046 24898 7098
rect 24898 7046 24908 7098
rect 24932 7046 24962 7098
rect 24962 7046 24974 7098
rect 24974 7046 24988 7098
rect 25012 7046 25026 7098
rect 25026 7046 25038 7098
rect 25038 7046 25068 7098
rect 25092 7046 25102 7098
rect 25102 7046 25148 7098
rect 24852 7044 24908 7046
rect 24932 7044 24988 7046
rect 25012 7044 25068 7046
rect 25092 7044 25148 7046
rect 24852 6010 24908 6012
rect 24932 6010 24988 6012
rect 25012 6010 25068 6012
rect 25092 6010 25148 6012
rect 24852 5958 24898 6010
rect 24898 5958 24908 6010
rect 24932 5958 24962 6010
rect 24962 5958 24974 6010
rect 24974 5958 24988 6010
rect 25012 5958 25026 6010
rect 25026 5958 25038 6010
rect 25038 5958 25068 6010
rect 25092 5958 25102 6010
rect 25102 5958 25148 6010
rect 24852 5956 24908 5958
rect 24932 5956 24988 5958
rect 25012 5956 25068 5958
rect 25092 5956 25148 5958
rect 24852 4922 24908 4924
rect 24932 4922 24988 4924
rect 25012 4922 25068 4924
rect 25092 4922 25148 4924
rect 24852 4870 24898 4922
rect 24898 4870 24908 4922
rect 24932 4870 24962 4922
rect 24962 4870 24974 4922
rect 24974 4870 24988 4922
rect 25012 4870 25026 4922
rect 25026 4870 25038 4922
rect 25038 4870 25068 4922
rect 25092 4870 25102 4922
rect 25102 4870 25148 4922
rect 24852 4868 24908 4870
rect 24932 4868 24988 4870
rect 25012 4868 25068 4870
rect 25092 4868 25148 4870
rect 24852 3834 24908 3836
rect 24932 3834 24988 3836
rect 25012 3834 25068 3836
rect 25092 3834 25148 3836
rect 24852 3782 24898 3834
rect 24898 3782 24908 3834
rect 24932 3782 24962 3834
rect 24962 3782 24974 3834
rect 24974 3782 24988 3834
rect 25012 3782 25026 3834
rect 25026 3782 25038 3834
rect 25038 3782 25068 3834
rect 25092 3782 25102 3834
rect 25102 3782 25148 3834
rect 24852 3780 24908 3782
rect 24932 3780 24988 3782
rect 25012 3780 25068 3782
rect 25092 3780 25148 3782
rect 24852 2746 24908 2748
rect 24932 2746 24988 2748
rect 25012 2746 25068 2748
rect 25092 2746 25148 2748
rect 24852 2694 24898 2746
rect 24898 2694 24908 2746
rect 24932 2694 24962 2746
rect 24962 2694 24974 2746
rect 24974 2694 24988 2746
rect 25012 2694 25026 2746
rect 25026 2694 25038 2746
rect 25038 2694 25068 2746
rect 25092 2694 25102 2746
rect 25102 2694 25148 2746
rect 24852 2692 24908 2694
rect 24932 2692 24988 2694
rect 25012 2692 25068 2694
rect 25092 2692 25148 2694
rect 32817 17434 32873 17436
rect 32897 17434 32953 17436
rect 32977 17434 33033 17436
rect 33057 17434 33113 17436
rect 32817 17382 32863 17434
rect 32863 17382 32873 17434
rect 32897 17382 32927 17434
rect 32927 17382 32939 17434
rect 32939 17382 32953 17434
rect 32977 17382 32991 17434
rect 32991 17382 33003 17434
rect 33003 17382 33033 17434
rect 33057 17382 33067 17434
rect 33067 17382 33113 17434
rect 32817 17380 32873 17382
rect 32897 17380 32953 17382
rect 32977 17380 33033 17382
rect 33057 17380 33113 17382
rect 32817 16346 32873 16348
rect 32897 16346 32953 16348
rect 32977 16346 33033 16348
rect 33057 16346 33113 16348
rect 32817 16294 32863 16346
rect 32863 16294 32873 16346
rect 32897 16294 32927 16346
rect 32927 16294 32939 16346
rect 32939 16294 32953 16346
rect 32977 16294 32991 16346
rect 32991 16294 33003 16346
rect 33003 16294 33033 16346
rect 33057 16294 33067 16346
rect 33067 16294 33113 16346
rect 32817 16292 32873 16294
rect 32897 16292 32953 16294
rect 32977 16292 33033 16294
rect 33057 16292 33113 16294
rect 32817 15258 32873 15260
rect 32897 15258 32953 15260
rect 32977 15258 33033 15260
rect 33057 15258 33113 15260
rect 32817 15206 32863 15258
rect 32863 15206 32873 15258
rect 32897 15206 32927 15258
rect 32927 15206 32939 15258
rect 32939 15206 32953 15258
rect 32977 15206 32991 15258
rect 32991 15206 33003 15258
rect 33003 15206 33033 15258
rect 33057 15206 33067 15258
rect 33067 15206 33113 15258
rect 32817 15204 32873 15206
rect 32897 15204 32953 15206
rect 32977 15204 33033 15206
rect 33057 15204 33113 15206
rect 40782 16890 40838 16892
rect 40862 16890 40918 16892
rect 40942 16890 40998 16892
rect 41022 16890 41078 16892
rect 40782 16838 40828 16890
rect 40828 16838 40838 16890
rect 40862 16838 40892 16890
rect 40892 16838 40904 16890
rect 40904 16838 40918 16890
rect 40942 16838 40956 16890
rect 40956 16838 40968 16890
rect 40968 16838 40998 16890
rect 41022 16838 41032 16890
rect 41032 16838 41078 16890
rect 40782 16836 40838 16838
rect 40862 16836 40918 16838
rect 40942 16836 40998 16838
rect 41022 16836 41078 16838
rect 32817 14170 32873 14172
rect 32897 14170 32953 14172
rect 32977 14170 33033 14172
rect 33057 14170 33113 14172
rect 32817 14118 32863 14170
rect 32863 14118 32873 14170
rect 32897 14118 32927 14170
rect 32927 14118 32939 14170
rect 32939 14118 32953 14170
rect 32977 14118 32991 14170
rect 32991 14118 33003 14170
rect 33003 14118 33033 14170
rect 33057 14118 33067 14170
rect 33067 14118 33113 14170
rect 32817 14116 32873 14118
rect 32897 14116 32953 14118
rect 32977 14116 33033 14118
rect 33057 14116 33113 14118
rect 32817 13082 32873 13084
rect 32897 13082 32953 13084
rect 32977 13082 33033 13084
rect 33057 13082 33113 13084
rect 32817 13030 32863 13082
rect 32863 13030 32873 13082
rect 32897 13030 32927 13082
rect 32927 13030 32939 13082
rect 32939 13030 32953 13082
rect 32977 13030 32991 13082
rect 32991 13030 33003 13082
rect 33003 13030 33033 13082
rect 33057 13030 33067 13082
rect 33067 13030 33113 13082
rect 32817 13028 32873 13030
rect 32897 13028 32953 13030
rect 32977 13028 33033 13030
rect 33057 13028 33113 13030
rect 32817 11994 32873 11996
rect 32897 11994 32953 11996
rect 32977 11994 33033 11996
rect 33057 11994 33113 11996
rect 32817 11942 32863 11994
rect 32863 11942 32873 11994
rect 32897 11942 32927 11994
rect 32927 11942 32939 11994
rect 32939 11942 32953 11994
rect 32977 11942 32991 11994
rect 32991 11942 33003 11994
rect 33003 11942 33033 11994
rect 33057 11942 33067 11994
rect 33067 11942 33113 11994
rect 32817 11940 32873 11942
rect 32897 11940 32953 11942
rect 32977 11940 33033 11942
rect 33057 11940 33113 11942
rect 32817 10906 32873 10908
rect 32897 10906 32953 10908
rect 32977 10906 33033 10908
rect 33057 10906 33113 10908
rect 32817 10854 32863 10906
rect 32863 10854 32873 10906
rect 32897 10854 32927 10906
rect 32927 10854 32939 10906
rect 32939 10854 32953 10906
rect 32977 10854 32991 10906
rect 32991 10854 33003 10906
rect 33003 10854 33033 10906
rect 33057 10854 33067 10906
rect 33067 10854 33113 10906
rect 32817 10852 32873 10854
rect 32897 10852 32953 10854
rect 32977 10852 33033 10854
rect 33057 10852 33113 10854
rect 32817 9818 32873 9820
rect 32897 9818 32953 9820
rect 32977 9818 33033 9820
rect 33057 9818 33113 9820
rect 32817 9766 32863 9818
rect 32863 9766 32873 9818
rect 32897 9766 32927 9818
rect 32927 9766 32939 9818
rect 32939 9766 32953 9818
rect 32977 9766 32991 9818
rect 32991 9766 33003 9818
rect 33003 9766 33033 9818
rect 33057 9766 33067 9818
rect 33067 9766 33113 9818
rect 32817 9764 32873 9766
rect 32897 9764 32953 9766
rect 32977 9764 33033 9766
rect 33057 9764 33113 9766
rect 32817 8730 32873 8732
rect 32897 8730 32953 8732
rect 32977 8730 33033 8732
rect 33057 8730 33113 8732
rect 32817 8678 32863 8730
rect 32863 8678 32873 8730
rect 32897 8678 32927 8730
rect 32927 8678 32939 8730
rect 32939 8678 32953 8730
rect 32977 8678 32991 8730
rect 32991 8678 33003 8730
rect 33003 8678 33033 8730
rect 33057 8678 33067 8730
rect 33067 8678 33113 8730
rect 32817 8676 32873 8678
rect 32897 8676 32953 8678
rect 32977 8676 33033 8678
rect 33057 8676 33113 8678
rect 32817 7642 32873 7644
rect 32897 7642 32953 7644
rect 32977 7642 33033 7644
rect 33057 7642 33113 7644
rect 32817 7590 32863 7642
rect 32863 7590 32873 7642
rect 32897 7590 32927 7642
rect 32927 7590 32939 7642
rect 32939 7590 32953 7642
rect 32977 7590 32991 7642
rect 32991 7590 33003 7642
rect 33003 7590 33033 7642
rect 33057 7590 33067 7642
rect 33067 7590 33113 7642
rect 32817 7588 32873 7590
rect 32897 7588 32953 7590
rect 32977 7588 33033 7590
rect 33057 7588 33113 7590
rect 32817 6554 32873 6556
rect 32897 6554 32953 6556
rect 32977 6554 33033 6556
rect 33057 6554 33113 6556
rect 32817 6502 32863 6554
rect 32863 6502 32873 6554
rect 32897 6502 32927 6554
rect 32927 6502 32939 6554
rect 32939 6502 32953 6554
rect 32977 6502 32991 6554
rect 32991 6502 33003 6554
rect 33003 6502 33033 6554
rect 33057 6502 33067 6554
rect 33067 6502 33113 6554
rect 32817 6500 32873 6502
rect 32897 6500 32953 6502
rect 32977 6500 33033 6502
rect 33057 6500 33113 6502
rect 32817 5466 32873 5468
rect 32897 5466 32953 5468
rect 32977 5466 33033 5468
rect 33057 5466 33113 5468
rect 32817 5414 32863 5466
rect 32863 5414 32873 5466
rect 32897 5414 32927 5466
rect 32927 5414 32939 5466
rect 32939 5414 32953 5466
rect 32977 5414 32991 5466
rect 32991 5414 33003 5466
rect 33003 5414 33033 5466
rect 33057 5414 33067 5466
rect 33067 5414 33113 5466
rect 32817 5412 32873 5414
rect 32897 5412 32953 5414
rect 32977 5412 33033 5414
rect 33057 5412 33113 5414
rect 32817 4378 32873 4380
rect 32897 4378 32953 4380
rect 32977 4378 33033 4380
rect 33057 4378 33113 4380
rect 32817 4326 32863 4378
rect 32863 4326 32873 4378
rect 32897 4326 32927 4378
rect 32927 4326 32939 4378
rect 32939 4326 32953 4378
rect 32977 4326 32991 4378
rect 32991 4326 33003 4378
rect 33003 4326 33033 4378
rect 33057 4326 33067 4378
rect 33067 4326 33113 4378
rect 32817 4324 32873 4326
rect 32897 4324 32953 4326
rect 32977 4324 33033 4326
rect 33057 4324 33113 4326
rect 32817 3290 32873 3292
rect 32897 3290 32953 3292
rect 32977 3290 33033 3292
rect 33057 3290 33113 3292
rect 32817 3238 32863 3290
rect 32863 3238 32873 3290
rect 32897 3238 32927 3290
rect 32927 3238 32939 3290
rect 32939 3238 32953 3290
rect 32977 3238 32991 3290
rect 32991 3238 33003 3290
rect 33003 3238 33033 3290
rect 33057 3238 33067 3290
rect 33067 3238 33113 3290
rect 32817 3236 32873 3238
rect 32897 3236 32953 3238
rect 32977 3236 33033 3238
rect 33057 3236 33113 3238
rect 32817 2202 32873 2204
rect 32897 2202 32953 2204
rect 32977 2202 33033 2204
rect 33057 2202 33113 2204
rect 32817 2150 32863 2202
rect 32863 2150 32873 2202
rect 32897 2150 32927 2202
rect 32927 2150 32939 2202
rect 32939 2150 32953 2202
rect 32977 2150 32991 2202
rect 32991 2150 33003 2202
rect 33003 2150 33033 2202
rect 33057 2150 33067 2202
rect 33067 2150 33113 2202
rect 32817 2148 32873 2150
rect 32897 2148 32953 2150
rect 32977 2148 33033 2150
rect 33057 2148 33113 2150
rect 40782 15802 40838 15804
rect 40862 15802 40918 15804
rect 40942 15802 40998 15804
rect 41022 15802 41078 15804
rect 40782 15750 40828 15802
rect 40828 15750 40838 15802
rect 40862 15750 40892 15802
rect 40892 15750 40904 15802
rect 40904 15750 40918 15802
rect 40942 15750 40956 15802
rect 40956 15750 40968 15802
rect 40968 15750 40998 15802
rect 41022 15750 41032 15802
rect 41032 15750 41078 15802
rect 40782 15748 40838 15750
rect 40862 15748 40918 15750
rect 40942 15748 40998 15750
rect 41022 15748 41078 15750
rect 46754 19080 46810 19136
rect 45558 17720 45614 17776
rect 40782 14714 40838 14716
rect 40862 14714 40918 14716
rect 40942 14714 40998 14716
rect 41022 14714 41078 14716
rect 40782 14662 40828 14714
rect 40828 14662 40838 14714
rect 40862 14662 40892 14714
rect 40892 14662 40904 14714
rect 40904 14662 40918 14714
rect 40942 14662 40956 14714
rect 40956 14662 40968 14714
rect 40968 14662 40998 14714
rect 41022 14662 41032 14714
rect 41032 14662 41078 14714
rect 40782 14660 40838 14662
rect 40862 14660 40918 14662
rect 40942 14660 40998 14662
rect 41022 14660 41078 14662
rect 40782 13626 40838 13628
rect 40862 13626 40918 13628
rect 40942 13626 40998 13628
rect 41022 13626 41078 13628
rect 40782 13574 40828 13626
rect 40828 13574 40838 13626
rect 40862 13574 40892 13626
rect 40892 13574 40904 13626
rect 40904 13574 40918 13626
rect 40942 13574 40956 13626
rect 40956 13574 40968 13626
rect 40968 13574 40998 13626
rect 41022 13574 41032 13626
rect 41032 13574 41078 13626
rect 40782 13572 40838 13574
rect 40862 13572 40918 13574
rect 40942 13572 40998 13574
rect 41022 13572 41078 13574
rect 40782 12538 40838 12540
rect 40862 12538 40918 12540
rect 40942 12538 40998 12540
rect 41022 12538 41078 12540
rect 40782 12486 40828 12538
rect 40828 12486 40838 12538
rect 40862 12486 40892 12538
rect 40892 12486 40904 12538
rect 40904 12486 40918 12538
rect 40942 12486 40956 12538
rect 40956 12486 40968 12538
rect 40968 12486 40998 12538
rect 41022 12486 41032 12538
rect 41032 12486 41078 12538
rect 40782 12484 40838 12486
rect 40862 12484 40918 12486
rect 40942 12484 40998 12486
rect 41022 12484 41078 12486
rect 40782 11450 40838 11452
rect 40862 11450 40918 11452
rect 40942 11450 40998 11452
rect 41022 11450 41078 11452
rect 40782 11398 40828 11450
rect 40828 11398 40838 11450
rect 40862 11398 40892 11450
rect 40892 11398 40904 11450
rect 40904 11398 40918 11450
rect 40942 11398 40956 11450
rect 40956 11398 40968 11450
rect 40968 11398 40998 11450
rect 41022 11398 41032 11450
rect 41032 11398 41078 11450
rect 40782 11396 40838 11398
rect 40862 11396 40918 11398
rect 40942 11396 40998 11398
rect 41022 11396 41078 11398
rect 40782 10362 40838 10364
rect 40862 10362 40918 10364
rect 40942 10362 40998 10364
rect 41022 10362 41078 10364
rect 40782 10310 40828 10362
rect 40828 10310 40838 10362
rect 40862 10310 40892 10362
rect 40892 10310 40904 10362
rect 40904 10310 40918 10362
rect 40942 10310 40956 10362
rect 40956 10310 40968 10362
rect 40968 10310 40998 10362
rect 41022 10310 41032 10362
rect 41032 10310 41078 10362
rect 40782 10308 40838 10310
rect 40862 10308 40918 10310
rect 40942 10308 40998 10310
rect 41022 10308 41078 10310
rect 40782 9274 40838 9276
rect 40862 9274 40918 9276
rect 40942 9274 40998 9276
rect 41022 9274 41078 9276
rect 40782 9222 40828 9274
rect 40828 9222 40838 9274
rect 40862 9222 40892 9274
rect 40892 9222 40904 9274
rect 40904 9222 40918 9274
rect 40942 9222 40956 9274
rect 40956 9222 40968 9274
rect 40968 9222 40998 9274
rect 41022 9222 41032 9274
rect 41032 9222 41078 9274
rect 40782 9220 40838 9222
rect 40862 9220 40918 9222
rect 40942 9220 40998 9222
rect 41022 9220 41078 9222
rect 40782 8186 40838 8188
rect 40862 8186 40918 8188
rect 40942 8186 40998 8188
rect 41022 8186 41078 8188
rect 40782 8134 40828 8186
rect 40828 8134 40838 8186
rect 40862 8134 40892 8186
rect 40892 8134 40904 8186
rect 40904 8134 40918 8186
rect 40942 8134 40956 8186
rect 40956 8134 40968 8186
rect 40968 8134 40998 8186
rect 41022 8134 41032 8186
rect 41032 8134 41078 8186
rect 40782 8132 40838 8134
rect 40862 8132 40918 8134
rect 40942 8132 40998 8134
rect 41022 8132 41078 8134
rect 40782 7098 40838 7100
rect 40862 7098 40918 7100
rect 40942 7098 40998 7100
rect 41022 7098 41078 7100
rect 40782 7046 40828 7098
rect 40828 7046 40838 7098
rect 40862 7046 40892 7098
rect 40892 7046 40904 7098
rect 40904 7046 40918 7098
rect 40942 7046 40956 7098
rect 40956 7046 40968 7098
rect 40968 7046 40998 7098
rect 41022 7046 41032 7098
rect 41032 7046 41078 7098
rect 40782 7044 40838 7046
rect 40862 7044 40918 7046
rect 40942 7044 40998 7046
rect 41022 7044 41078 7046
rect 40782 6010 40838 6012
rect 40862 6010 40918 6012
rect 40942 6010 40998 6012
rect 41022 6010 41078 6012
rect 40782 5958 40828 6010
rect 40828 5958 40838 6010
rect 40862 5958 40892 6010
rect 40892 5958 40904 6010
rect 40904 5958 40918 6010
rect 40942 5958 40956 6010
rect 40956 5958 40968 6010
rect 40968 5958 40998 6010
rect 41022 5958 41032 6010
rect 41032 5958 41078 6010
rect 40782 5956 40838 5958
rect 40862 5956 40918 5958
rect 40942 5956 40998 5958
rect 41022 5956 41078 5958
rect 40782 4922 40838 4924
rect 40862 4922 40918 4924
rect 40942 4922 40998 4924
rect 41022 4922 41078 4924
rect 40782 4870 40828 4922
rect 40828 4870 40838 4922
rect 40862 4870 40892 4922
rect 40892 4870 40904 4922
rect 40904 4870 40918 4922
rect 40942 4870 40956 4922
rect 40956 4870 40968 4922
rect 40968 4870 40998 4922
rect 41022 4870 41032 4922
rect 41032 4870 41078 4922
rect 40782 4868 40838 4870
rect 40862 4868 40918 4870
rect 40942 4868 40998 4870
rect 41022 4868 41078 4870
rect 46570 17040 46626 17096
rect 46846 16360 46902 16416
rect 46846 13640 46902 13696
rect 46846 12280 46902 12336
rect 46846 11636 46848 11656
rect 46848 11636 46900 11656
rect 46900 11636 46902 11656
rect 46846 11600 46902 11636
rect 46754 7520 46810 7576
rect 40782 3834 40838 3836
rect 40862 3834 40918 3836
rect 40942 3834 40998 3836
rect 41022 3834 41078 3836
rect 40782 3782 40828 3834
rect 40828 3782 40838 3834
rect 40862 3782 40892 3834
rect 40892 3782 40904 3834
rect 40904 3782 40918 3834
rect 40942 3782 40956 3834
rect 40956 3782 40968 3834
rect 40968 3782 40998 3834
rect 41022 3782 41032 3834
rect 41032 3782 41078 3834
rect 40782 3780 40838 3782
rect 40862 3780 40918 3782
rect 40942 3780 40998 3782
rect 41022 3780 41078 3782
rect 40782 2746 40838 2748
rect 40862 2746 40918 2748
rect 40942 2746 40998 2748
rect 41022 2746 41078 2748
rect 40782 2694 40828 2746
rect 40828 2694 40838 2746
rect 40862 2694 40892 2746
rect 40892 2694 40904 2746
rect 40904 2694 40918 2746
rect 40942 2694 40956 2746
rect 40956 2694 40968 2746
rect 40968 2694 40998 2746
rect 41022 2694 41032 2746
rect 41032 2694 41078 2746
rect 40782 2692 40838 2694
rect 40862 2692 40918 2694
rect 40942 2692 40998 2694
rect 41022 2692 41078 2694
rect 46662 5480 46718 5536
rect 46570 4800 46626 4856
rect 46846 4120 46902 4176
rect 46846 3440 46902 3496
rect 45650 1400 45706 1456
rect 48134 15000 48190 15056
rect 48134 12960 48190 13016
rect 48134 10920 48190 10976
rect 48134 10240 48190 10296
rect 48134 2760 48190 2816
rect 46846 720 46902 776
rect 46662 40 46718 96
<< metal3 >>
rect 0 19668 800 19908
rect 0 18988 800 19228
rect 46749 19138 46815 19141
rect 49200 19138 50000 19228
rect 46749 19136 50000 19138
rect 46749 19080 46754 19136
rect 46810 19080 50000 19136
rect 46749 19078 50000 19080
rect 46749 19075 46815 19078
rect 49200 18988 50000 19078
rect 0 18308 800 18548
rect 49200 18308 50000 18548
rect 0 17778 800 17868
rect 1393 17778 1459 17781
rect 0 17776 1459 17778
rect 0 17720 1398 17776
rect 1454 17720 1459 17776
rect 0 17718 1459 17720
rect 0 17628 800 17718
rect 1393 17715 1459 17718
rect 45553 17778 45619 17781
rect 49200 17778 50000 17868
rect 45553 17776 50000 17778
rect 45553 17720 45558 17776
rect 45614 17720 50000 17776
rect 45553 17718 50000 17720
rect 45553 17715 45619 17718
rect 49200 17628 50000 17718
rect 16874 17440 17194 17441
rect 16874 17376 16882 17440
rect 16946 17376 16962 17440
rect 17026 17376 17042 17440
rect 17106 17376 17122 17440
rect 17186 17376 17194 17440
rect 16874 17375 17194 17376
rect 32805 17440 33125 17441
rect 32805 17376 32813 17440
rect 32877 17376 32893 17440
rect 32957 17376 32973 17440
rect 33037 17376 33053 17440
rect 33117 17376 33125 17440
rect 32805 17375 33125 17376
rect 0 17098 800 17188
rect 4061 17098 4127 17101
rect 0 17096 4127 17098
rect 0 17040 4066 17096
rect 4122 17040 4127 17096
rect 0 17038 4127 17040
rect 0 16948 800 17038
rect 4061 17035 4127 17038
rect 46565 17098 46631 17101
rect 49200 17098 50000 17188
rect 46565 17096 50000 17098
rect 46565 17040 46570 17096
rect 46626 17040 50000 17096
rect 46565 17038 50000 17040
rect 46565 17035 46631 17038
rect 49200 16948 50000 17038
rect 8909 16896 9229 16897
rect 8909 16832 8917 16896
rect 8981 16832 8997 16896
rect 9061 16832 9077 16896
rect 9141 16832 9157 16896
rect 9221 16832 9229 16896
rect 8909 16831 9229 16832
rect 24840 16896 25160 16897
rect 24840 16832 24848 16896
rect 24912 16832 24928 16896
rect 24992 16832 25008 16896
rect 25072 16832 25088 16896
rect 25152 16832 25160 16896
rect 24840 16831 25160 16832
rect 40770 16896 41090 16897
rect 40770 16832 40778 16896
rect 40842 16832 40858 16896
rect 40922 16832 40938 16896
rect 41002 16832 41018 16896
rect 41082 16832 41090 16896
rect 40770 16831 41090 16832
rect 0 16268 800 16508
rect 46841 16418 46907 16421
rect 49200 16418 50000 16508
rect 46841 16416 50000 16418
rect 46841 16360 46846 16416
rect 46902 16360 50000 16416
rect 46841 16358 50000 16360
rect 46841 16355 46907 16358
rect 16874 16352 17194 16353
rect 16874 16288 16882 16352
rect 16946 16288 16962 16352
rect 17026 16288 17042 16352
rect 17106 16288 17122 16352
rect 17186 16288 17194 16352
rect 16874 16287 17194 16288
rect 32805 16352 33125 16353
rect 32805 16288 32813 16352
rect 32877 16288 32893 16352
rect 32957 16288 32973 16352
rect 33037 16288 33053 16352
rect 33117 16288 33125 16352
rect 32805 16287 33125 16288
rect 49200 16268 50000 16358
rect 0 15738 800 15828
rect 8909 15808 9229 15809
rect 8909 15744 8917 15808
rect 8981 15744 8997 15808
rect 9061 15744 9077 15808
rect 9141 15744 9157 15808
rect 9221 15744 9229 15808
rect 8909 15743 9229 15744
rect 24840 15808 25160 15809
rect 24840 15744 24848 15808
rect 24912 15744 24928 15808
rect 24992 15744 25008 15808
rect 25072 15744 25088 15808
rect 25152 15744 25160 15808
rect 24840 15743 25160 15744
rect 40770 15808 41090 15809
rect 40770 15744 40778 15808
rect 40842 15744 40858 15808
rect 40922 15744 40938 15808
rect 41002 15744 41018 15808
rect 41082 15744 41090 15808
rect 40770 15743 41090 15744
rect 2773 15738 2839 15741
rect 0 15736 2839 15738
rect 0 15680 2778 15736
rect 2834 15680 2839 15736
rect 0 15678 2839 15680
rect 0 15588 800 15678
rect 2773 15675 2839 15678
rect 49200 15588 50000 15828
rect 16874 15264 17194 15265
rect 16874 15200 16882 15264
rect 16946 15200 16962 15264
rect 17026 15200 17042 15264
rect 17106 15200 17122 15264
rect 17186 15200 17194 15264
rect 16874 15199 17194 15200
rect 32805 15264 33125 15265
rect 32805 15200 32813 15264
rect 32877 15200 32893 15264
rect 32957 15200 32973 15264
rect 33037 15200 33053 15264
rect 33117 15200 33125 15264
rect 32805 15199 33125 15200
rect 0 14908 800 15148
rect 48129 15058 48195 15061
rect 49200 15058 50000 15148
rect 48129 15056 50000 15058
rect 48129 15000 48134 15056
rect 48190 15000 50000 15056
rect 48129 14998 50000 15000
rect 48129 14995 48195 14998
rect 49200 14908 50000 14998
rect 8909 14720 9229 14721
rect 8909 14656 8917 14720
rect 8981 14656 8997 14720
rect 9061 14656 9077 14720
rect 9141 14656 9157 14720
rect 9221 14656 9229 14720
rect 8909 14655 9229 14656
rect 24840 14720 25160 14721
rect 24840 14656 24848 14720
rect 24912 14656 24928 14720
rect 24992 14656 25008 14720
rect 25072 14656 25088 14720
rect 25152 14656 25160 14720
rect 24840 14655 25160 14656
rect 40770 14720 41090 14721
rect 40770 14656 40778 14720
rect 40842 14656 40858 14720
rect 40922 14656 40938 14720
rect 41002 14656 41018 14720
rect 41082 14656 41090 14720
rect 40770 14655 41090 14656
rect 0 14378 800 14468
rect 2773 14378 2839 14381
rect 0 14376 2839 14378
rect 0 14320 2778 14376
rect 2834 14320 2839 14376
rect 0 14318 2839 14320
rect 0 14228 800 14318
rect 2773 14315 2839 14318
rect 49200 14228 50000 14468
rect 16874 14176 17194 14177
rect 16874 14112 16882 14176
rect 16946 14112 16962 14176
rect 17026 14112 17042 14176
rect 17106 14112 17122 14176
rect 17186 14112 17194 14176
rect 16874 14111 17194 14112
rect 32805 14176 33125 14177
rect 32805 14112 32813 14176
rect 32877 14112 32893 14176
rect 32957 14112 32973 14176
rect 33037 14112 33053 14176
rect 33117 14112 33125 14176
rect 32805 14111 33125 14112
rect 0 13548 800 13788
rect 46841 13698 46907 13701
rect 49200 13698 50000 13788
rect 46841 13696 50000 13698
rect 46841 13640 46846 13696
rect 46902 13640 50000 13696
rect 46841 13638 50000 13640
rect 46841 13635 46907 13638
rect 8909 13632 9229 13633
rect 8909 13568 8917 13632
rect 8981 13568 8997 13632
rect 9061 13568 9077 13632
rect 9141 13568 9157 13632
rect 9221 13568 9229 13632
rect 8909 13567 9229 13568
rect 24840 13632 25160 13633
rect 24840 13568 24848 13632
rect 24912 13568 24928 13632
rect 24992 13568 25008 13632
rect 25072 13568 25088 13632
rect 25152 13568 25160 13632
rect 24840 13567 25160 13568
rect 40770 13632 41090 13633
rect 40770 13568 40778 13632
rect 40842 13568 40858 13632
rect 40922 13568 40938 13632
rect 41002 13568 41018 13632
rect 41082 13568 41090 13632
rect 40770 13567 41090 13568
rect 49200 13548 50000 13638
rect 0 13018 800 13108
rect 16874 13088 17194 13089
rect 16874 13024 16882 13088
rect 16946 13024 16962 13088
rect 17026 13024 17042 13088
rect 17106 13024 17122 13088
rect 17186 13024 17194 13088
rect 16874 13023 17194 13024
rect 32805 13088 33125 13089
rect 32805 13024 32813 13088
rect 32877 13024 32893 13088
rect 32957 13024 32973 13088
rect 33037 13024 33053 13088
rect 33117 13024 33125 13088
rect 32805 13023 33125 13024
rect 2773 13018 2839 13021
rect 0 13016 2839 13018
rect 0 12960 2778 13016
rect 2834 12960 2839 13016
rect 0 12958 2839 12960
rect 0 12868 800 12958
rect 2773 12955 2839 12958
rect 48129 13018 48195 13021
rect 49200 13018 50000 13108
rect 48129 13016 50000 13018
rect 48129 12960 48134 13016
rect 48190 12960 50000 13016
rect 48129 12958 50000 12960
rect 48129 12955 48195 12958
rect 49200 12868 50000 12958
rect 8909 12544 9229 12545
rect 8909 12480 8917 12544
rect 8981 12480 8997 12544
rect 9061 12480 9077 12544
rect 9141 12480 9157 12544
rect 9221 12480 9229 12544
rect 8909 12479 9229 12480
rect 24840 12544 25160 12545
rect 24840 12480 24848 12544
rect 24912 12480 24928 12544
rect 24992 12480 25008 12544
rect 25072 12480 25088 12544
rect 25152 12480 25160 12544
rect 24840 12479 25160 12480
rect 40770 12544 41090 12545
rect 40770 12480 40778 12544
rect 40842 12480 40858 12544
rect 40922 12480 40938 12544
rect 41002 12480 41018 12544
rect 41082 12480 41090 12544
rect 40770 12479 41090 12480
rect 0 12338 800 12428
rect 4061 12338 4127 12341
rect 0 12336 4127 12338
rect 0 12280 4066 12336
rect 4122 12280 4127 12336
rect 0 12278 4127 12280
rect 0 12188 800 12278
rect 4061 12275 4127 12278
rect 46841 12338 46907 12341
rect 49200 12338 50000 12428
rect 46841 12336 50000 12338
rect 46841 12280 46846 12336
rect 46902 12280 50000 12336
rect 46841 12278 50000 12280
rect 46841 12275 46907 12278
rect 49200 12188 50000 12278
rect 16874 12000 17194 12001
rect 16874 11936 16882 12000
rect 16946 11936 16962 12000
rect 17026 11936 17042 12000
rect 17106 11936 17122 12000
rect 17186 11936 17194 12000
rect 16874 11935 17194 11936
rect 32805 12000 33125 12001
rect 32805 11936 32813 12000
rect 32877 11936 32893 12000
rect 32957 11936 32973 12000
rect 33037 11936 33053 12000
rect 33117 11936 33125 12000
rect 32805 11935 33125 11936
rect 0 11508 800 11748
rect 46841 11658 46907 11661
rect 49200 11658 50000 11748
rect 46841 11656 50000 11658
rect 46841 11600 46846 11656
rect 46902 11600 50000 11656
rect 46841 11598 50000 11600
rect 46841 11595 46907 11598
rect 49200 11508 50000 11598
rect 8909 11456 9229 11457
rect 8909 11392 8917 11456
rect 8981 11392 8997 11456
rect 9061 11392 9077 11456
rect 9141 11392 9157 11456
rect 9221 11392 9229 11456
rect 8909 11391 9229 11392
rect 24840 11456 25160 11457
rect 24840 11392 24848 11456
rect 24912 11392 24928 11456
rect 24992 11392 25008 11456
rect 25072 11392 25088 11456
rect 25152 11392 25160 11456
rect 24840 11391 25160 11392
rect 40770 11456 41090 11457
rect 40770 11392 40778 11456
rect 40842 11392 40858 11456
rect 40922 11392 40938 11456
rect 41002 11392 41018 11456
rect 41082 11392 41090 11456
rect 40770 11391 41090 11392
rect 0 10978 800 11068
rect 2773 10978 2839 10981
rect 0 10976 2839 10978
rect 0 10920 2778 10976
rect 2834 10920 2839 10976
rect 0 10918 2839 10920
rect 0 10828 800 10918
rect 2773 10915 2839 10918
rect 48129 10978 48195 10981
rect 49200 10978 50000 11068
rect 48129 10976 50000 10978
rect 48129 10920 48134 10976
rect 48190 10920 50000 10976
rect 48129 10918 50000 10920
rect 48129 10915 48195 10918
rect 16874 10912 17194 10913
rect 16874 10848 16882 10912
rect 16946 10848 16962 10912
rect 17026 10848 17042 10912
rect 17106 10848 17122 10912
rect 17186 10848 17194 10912
rect 16874 10847 17194 10848
rect 32805 10912 33125 10913
rect 32805 10848 32813 10912
rect 32877 10848 32893 10912
rect 32957 10848 32973 10912
rect 33037 10848 33053 10912
rect 33117 10848 33125 10912
rect 32805 10847 33125 10848
rect 49200 10828 50000 10918
rect 0 10298 800 10388
rect 8909 10368 9229 10369
rect 8909 10304 8917 10368
rect 8981 10304 8997 10368
rect 9061 10304 9077 10368
rect 9141 10304 9157 10368
rect 9221 10304 9229 10368
rect 8909 10303 9229 10304
rect 24840 10368 25160 10369
rect 24840 10304 24848 10368
rect 24912 10304 24928 10368
rect 24992 10304 25008 10368
rect 25072 10304 25088 10368
rect 25152 10304 25160 10368
rect 24840 10303 25160 10304
rect 40770 10368 41090 10369
rect 40770 10304 40778 10368
rect 40842 10304 40858 10368
rect 40922 10304 40938 10368
rect 41002 10304 41018 10368
rect 41082 10304 41090 10368
rect 40770 10303 41090 10304
rect 3417 10298 3483 10301
rect 0 10296 3483 10298
rect 0 10240 3422 10296
rect 3478 10240 3483 10296
rect 0 10238 3483 10240
rect 0 10148 800 10238
rect 3417 10235 3483 10238
rect 48129 10298 48195 10301
rect 49200 10298 50000 10388
rect 48129 10296 50000 10298
rect 48129 10240 48134 10296
rect 48190 10240 50000 10296
rect 48129 10238 50000 10240
rect 48129 10235 48195 10238
rect 49200 10148 50000 10238
rect 16874 9824 17194 9825
rect 16874 9760 16882 9824
rect 16946 9760 16962 9824
rect 17026 9760 17042 9824
rect 17106 9760 17122 9824
rect 17186 9760 17194 9824
rect 16874 9759 17194 9760
rect 32805 9824 33125 9825
rect 32805 9760 32813 9824
rect 32877 9760 32893 9824
rect 32957 9760 32973 9824
rect 33037 9760 33053 9824
rect 33117 9760 33125 9824
rect 32805 9759 33125 9760
rect 0 9468 800 9708
rect 49200 9468 50000 9708
rect 8909 9280 9229 9281
rect 8909 9216 8917 9280
rect 8981 9216 8997 9280
rect 9061 9216 9077 9280
rect 9141 9216 9157 9280
rect 9221 9216 9229 9280
rect 8909 9215 9229 9216
rect 24840 9280 25160 9281
rect 24840 9216 24848 9280
rect 24912 9216 24928 9280
rect 24992 9216 25008 9280
rect 25072 9216 25088 9280
rect 25152 9216 25160 9280
rect 24840 9215 25160 9216
rect 40770 9280 41090 9281
rect 40770 9216 40778 9280
rect 40842 9216 40858 9280
rect 40922 9216 40938 9280
rect 41002 9216 41018 9280
rect 41082 9216 41090 9280
rect 40770 9215 41090 9216
rect 0 8788 800 9028
rect 49200 8788 50000 9028
rect 16874 8736 17194 8737
rect 16874 8672 16882 8736
rect 16946 8672 16962 8736
rect 17026 8672 17042 8736
rect 17106 8672 17122 8736
rect 17186 8672 17194 8736
rect 16874 8671 17194 8672
rect 32805 8736 33125 8737
rect 32805 8672 32813 8736
rect 32877 8672 32893 8736
rect 32957 8672 32973 8736
rect 33037 8672 33053 8736
rect 33117 8672 33125 8736
rect 32805 8671 33125 8672
rect 0 8258 800 8348
rect 2773 8258 2839 8261
rect 0 8256 2839 8258
rect 0 8200 2778 8256
rect 2834 8200 2839 8256
rect 0 8198 2839 8200
rect 0 8108 800 8198
rect 2773 8195 2839 8198
rect 8909 8192 9229 8193
rect 8909 8128 8917 8192
rect 8981 8128 8997 8192
rect 9061 8128 9077 8192
rect 9141 8128 9157 8192
rect 9221 8128 9229 8192
rect 8909 8127 9229 8128
rect 24840 8192 25160 8193
rect 24840 8128 24848 8192
rect 24912 8128 24928 8192
rect 24992 8128 25008 8192
rect 25072 8128 25088 8192
rect 25152 8128 25160 8192
rect 24840 8127 25160 8128
rect 40770 8192 41090 8193
rect 40770 8128 40778 8192
rect 40842 8128 40858 8192
rect 40922 8128 40938 8192
rect 41002 8128 41018 8192
rect 41082 8128 41090 8192
rect 40770 8127 41090 8128
rect 49200 8108 50000 8348
rect 0 7578 800 7668
rect 16874 7648 17194 7649
rect 16874 7584 16882 7648
rect 16946 7584 16962 7648
rect 17026 7584 17042 7648
rect 17106 7584 17122 7648
rect 17186 7584 17194 7648
rect 16874 7583 17194 7584
rect 32805 7648 33125 7649
rect 32805 7584 32813 7648
rect 32877 7584 32893 7648
rect 32957 7584 32973 7648
rect 33037 7584 33053 7648
rect 33117 7584 33125 7648
rect 32805 7583 33125 7584
rect 3417 7578 3483 7581
rect 0 7576 3483 7578
rect 0 7520 3422 7576
rect 3478 7520 3483 7576
rect 0 7518 3483 7520
rect 0 7428 800 7518
rect 3417 7515 3483 7518
rect 46749 7578 46815 7581
rect 49200 7578 50000 7668
rect 46749 7576 50000 7578
rect 46749 7520 46754 7576
rect 46810 7520 50000 7576
rect 46749 7518 50000 7520
rect 46749 7515 46815 7518
rect 49200 7428 50000 7518
rect 8909 7104 9229 7105
rect 8909 7040 8917 7104
rect 8981 7040 8997 7104
rect 9061 7040 9077 7104
rect 9141 7040 9157 7104
rect 9221 7040 9229 7104
rect 8909 7039 9229 7040
rect 24840 7104 25160 7105
rect 24840 7040 24848 7104
rect 24912 7040 24928 7104
rect 24992 7040 25008 7104
rect 25072 7040 25088 7104
rect 25152 7040 25160 7104
rect 24840 7039 25160 7040
rect 40770 7104 41090 7105
rect 40770 7040 40778 7104
rect 40842 7040 40858 7104
rect 40922 7040 40938 7104
rect 41002 7040 41018 7104
rect 41082 7040 41090 7104
rect 40770 7039 41090 7040
rect 0 6898 800 6988
rect 2773 6898 2839 6901
rect 0 6896 2839 6898
rect 0 6840 2778 6896
rect 2834 6840 2839 6896
rect 0 6838 2839 6840
rect 0 6748 800 6838
rect 2773 6835 2839 6838
rect 49200 6748 50000 6988
rect 16874 6560 17194 6561
rect 16874 6496 16882 6560
rect 16946 6496 16962 6560
rect 17026 6496 17042 6560
rect 17106 6496 17122 6560
rect 17186 6496 17194 6560
rect 16874 6495 17194 6496
rect 32805 6560 33125 6561
rect 32805 6496 32813 6560
rect 32877 6496 32893 6560
rect 32957 6496 32973 6560
rect 33037 6496 33053 6560
rect 33117 6496 33125 6560
rect 32805 6495 33125 6496
rect 0 6068 800 6308
rect 49200 6068 50000 6308
rect 8909 6016 9229 6017
rect 8909 5952 8917 6016
rect 8981 5952 8997 6016
rect 9061 5952 9077 6016
rect 9141 5952 9157 6016
rect 9221 5952 9229 6016
rect 8909 5951 9229 5952
rect 24840 6016 25160 6017
rect 24840 5952 24848 6016
rect 24912 5952 24928 6016
rect 24992 5952 25008 6016
rect 25072 5952 25088 6016
rect 25152 5952 25160 6016
rect 24840 5951 25160 5952
rect 40770 6016 41090 6017
rect 40770 5952 40778 6016
rect 40842 5952 40858 6016
rect 40922 5952 40938 6016
rect 41002 5952 41018 6016
rect 41082 5952 41090 6016
rect 40770 5951 41090 5952
rect 0 5538 800 5628
rect 2773 5538 2839 5541
rect 0 5536 2839 5538
rect 0 5480 2778 5536
rect 2834 5480 2839 5536
rect 0 5478 2839 5480
rect 0 5388 800 5478
rect 2773 5475 2839 5478
rect 46657 5538 46723 5541
rect 49200 5538 50000 5628
rect 46657 5536 50000 5538
rect 46657 5480 46662 5536
rect 46718 5480 50000 5536
rect 46657 5478 50000 5480
rect 46657 5475 46723 5478
rect 16874 5472 17194 5473
rect 16874 5408 16882 5472
rect 16946 5408 16962 5472
rect 17026 5408 17042 5472
rect 17106 5408 17122 5472
rect 17186 5408 17194 5472
rect 16874 5407 17194 5408
rect 32805 5472 33125 5473
rect 32805 5408 32813 5472
rect 32877 5408 32893 5472
rect 32957 5408 32973 5472
rect 33037 5408 33053 5472
rect 33117 5408 33125 5472
rect 32805 5407 33125 5408
rect 49200 5388 50000 5478
rect 0 4858 800 4948
rect 8909 4928 9229 4929
rect 8909 4864 8917 4928
rect 8981 4864 8997 4928
rect 9061 4864 9077 4928
rect 9141 4864 9157 4928
rect 9221 4864 9229 4928
rect 8909 4863 9229 4864
rect 24840 4928 25160 4929
rect 24840 4864 24848 4928
rect 24912 4864 24928 4928
rect 24992 4864 25008 4928
rect 25072 4864 25088 4928
rect 25152 4864 25160 4928
rect 24840 4863 25160 4864
rect 40770 4928 41090 4929
rect 40770 4864 40778 4928
rect 40842 4864 40858 4928
rect 40922 4864 40938 4928
rect 41002 4864 41018 4928
rect 41082 4864 41090 4928
rect 40770 4863 41090 4864
rect 1393 4858 1459 4861
rect 0 4856 1459 4858
rect 0 4800 1398 4856
rect 1454 4800 1459 4856
rect 0 4798 1459 4800
rect 0 4708 800 4798
rect 1393 4795 1459 4798
rect 46565 4858 46631 4861
rect 49200 4858 50000 4948
rect 46565 4856 50000 4858
rect 46565 4800 46570 4856
rect 46626 4800 50000 4856
rect 46565 4798 50000 4800
rect 46565 4795 46631 4798
rect 49200 4708 50000 4798
rect 16874 4384 17194 4385
rect 16874 4320 16882 4384
rect 16946 4320 16962 4384
rect 17026 4320 17042 4384
rect 17106 4320 17122 4384
rect 17186 4320 17194 4384
rect 16874 4319 17194 4320
rect 32805 4384 33125 4385
rect 32805 4320 32813 4384
rect 32877 4320 32893 4384
rect 32957 4320 32973 4384
rect 33037 4320 33053 4384
rect 33117 4320 33125 4384
rect 32805 4319 33125 4320
rect 0 4178 800 4268
rect 2773 4178 2839 4181
rect 0 4176 2839 4178
rect 0 4120 2778 4176
rect 2834 4120 2839 4176
rect 0 4118 2839 4120
rect 0 4028 800 4118
rect 2773 4115 2839 4118
rect 46841 4178 46907 4181
rect 49200 4178 50000 4268
rect 46841 4176 50000 4178
rect 46841 4120 46846 4176
rect 46902 4120 50000 4176
rect 46841 4118 50000 4120
rect 46841 4115 46907 4118
rect 49200 4028 50000 4118
rect 8909 3840 9229 3841
rect 8909 3776 8917 3840
rect 8981 3776 8997 3840
rect 9061 3776 9077 3840
rect 9141 3776 9157 3840
rect 9221 3776 9229 3840
rect 8909 3775 9229 3776
rect 24840 3840 25160 3841
rect 24840 3776 24848 3840
rect 24912 3776 24928 3840
rect 24992 3776 25008 3840
rect 25072 3776 25088 3840
rect 25152 3776 25160 3840
rect 24840 3775 25160 3776
rect 40770 3840 41090 3841
rect 40770 3776 40778 3840
rect 40842 3776 40858 3840
rect 40922 3776 40938 3840
rect 41002 3776 41018 3840
rect 41082 3776 41090 3840
rect 40770 3775 41090 3776
rect 0 3498 800 3588
rect 3969 3498 4035 3501
rect 0 3496 4035 3498
rect 0 3440 3974 3496
rect 4030 3440 4035 3496
rect 0 3438 4035 3440
rect 0 3348 800 3438
rect 3969 3435 4035 3438
rect 46841 3498 46907 3501
rect 49200 3498 50000 3588
rect 46841 3496 50000 3498
rect 46841 3440 46846 3496
rect 46902 3440 50000 3496
rect 46841 3438 50000 3440
rect 46841 3435 46907 3438
rect 49200 3348 50000 3438
rect 16874 3296 17194 3297
rect 16874 3232 16882 3296
rect 16946 3232 16962 3296
rect 17026 3232 17042 3296
rect 17106 3232 17122 3296
rect 17186 3232 17194 3296
rect 16874 3231 17194 3232
rect 32805 3296 33125 3297
rect 32805 3232 32813 3296
rect 32877 3232 32893 3296
rect 32957 3232 32973 3296
rect 33037 3232 33053 3296
rect 33117 3232 33125 3296
rect 32805 3231 33125 3232
rect 0 2818 800 2908
rect 2865 2818 2931 2821
rect 0 2816 2931 2818
rect 0 2760 2870 2816
rect 2926 2760 2931 2816
rect 0 2758 2931 2760
rect 0 2668 800 2758
rect 2865 2755 2931 2758
rect 48129 2818 48195 2821
rect 49200 2818 50000 2908
rect 48129 2816 50000 2818
rect 48129 2760 48134 2816
rect 48190 2760 50000 2816
rect 48129 2758 50000 2760
rect 48129 2755 48195 2758
rect 8909 2752 9229 2753
rect 8909 2688 8917 2752
rect 8981 2688 8997 2752
rect 9061 2688 9077 2752
rect 9141 2688 9157 2752
rect 9221 2688 9229 2752
rect 8909 2687 9229 2688
rect 24840 2752 25160 2753
rect 24840 2688 24848 2752
rect 24912 2688 24928 2752
rect 24992 2688 25008 2752
rect 25072 2688 25088 2752
rect 25152 2688 25160 2752
rect 24840 2687 25160 2688
rect 40770 2752 41090 2753
rect 40770 2688 40778 2752
rect 40842 2688 40858 2752
rect 40922 2688 40938 2752
rect 41002 2688 41018 2752
rect 41082 2688 41090 2752
rect 40770 2687 41090 2688
rect 49200 2668 50000 2758
rect 0 2138 800 2228
rect 16874 2208 17194 2209
rect 16874 2144 16882 2208
rect 16946 2144 16962 2208
rect 17026 2144 17042 2208
rect 17106 2144 17122 2208
rect 17186 2144 17194 2208
rect 16874 2143 17194 2144
rect 32805 2208 33125 2209
rect 32805 2144 32813 2208
rect 32877 2144 32893 2208
rect 32957 2144 32973 2208
rect 33037 2144 33053 2208
rect 33117 2144 33125 2208
rect 32805 2143 33125 2144
rect 3417 2138 3483 2141
rect 0 2136 3483 2138
rect 0 2080 3422 2136
rect 3478 2080 3483 2136
rect 0 2078 3483 2080
rect 0 1988 800 2078
rect 3417 2075 3483 2078
rect 49200 1988 50000 2228
rect 0 1458 800 1548
rect 3509 1458 3575 1461
rect 0 1456 3575 1458
rect 0 1400 3514 1456
rect 3570 1400 3575 1456
rect 0 1398 3575 1400
rect 0 1308 800 1398
rect 3509 1395 3575 1398
rect 45645 1458 45711 1461
rect 49200 1458 50000 1548
rect 45645 1456 50000 1458
rect 45645 1400 45650 1456
rect 45706 1400 50000 1456
rect 45645 1398 50000 1400
rect 45645 1395 45711 1398
rect 49200 1308 50000 1398
rect 0 628 800 868
rect 46841 778 46907 781
rect 49200 778 50000 868
rect 46841 776 50000 778
rect 46841 720 46846 776
rect 46902 720 50000 776
rect 46841 718 50000 720
rect 46841 715 46907 718
rect 49200 628 50000 718
rect 46657 98 46723 101
rect 49200 98 50000 188
rect 46657 96 50000 98
rect 46657 40 46662 96
rect 46718 40 50000 96
rect 46657 38 50000 40
rect 46657 35 46723 38
rect 49200 -52 50000 38
<< via3 >>
rect 16882 17436 16946 17440
rect 16882 17380 16886 17436
rect 16886 17380 16942 17436
rect 16942 17380 16946 17436
rect 16882 17376 16946 17380
rect 16962 17436 17026 17440
rect 16962 17380 16966 17436
rect 16966 17380 17022 17436
rect 17022 17380 17026 17436
rect 16962 17376 17026 17380
rect 17042 17436 17106 17440
rect 17042 17380 17046 17436
rect 17046 17380 17102 17436
rect 17102 17380 17106 17436
rect 17042 17376 17106 17380
rect 17122 17436 17186 17440
rect 17122 17380 17126 17436
rect 17126 17380 17182 17436
rect 17182 17380 17186 17436
rect 17122 17376 17186 17380
rect 32813 17436 32877 17440
rect 32813 17380 32817 17436
rect 32817 17380 32873 17436
rect 32873 17380 32877 17436
rect 32813 17376 32877 17380
rect 32893 17436 32957 17440
rect 32893 17380 32897 17436
rect 32897 17380 32953 17436
rect 32953 17380 32957 17436
rect 32893 17376 32957 17380
rect 32973 17436 33037 17440
rect 32973 17380 32977 17436
rect 32977 17380 33033 17436
rect 33033 17380 33037 17436
rect 32973 17376 33037 17380
rect 33053 17436 33117 17440
rect 33053 17380 33057 17436
rect 33057 17380 33113 17436
rect 33113 17380 33117 17436
rect 33053 17376 33117 17380
rect 8917 16892 8981 16896
rect 8917 16836 8921 16892
rect 8921 16836 8977 16892
rect 8977 16836 8981 16892
rect 8917 16832 8981 16836
rect 8997 16892 9061 16896
rect 8997 16836 9001 16892
rect 9001 16836 9057 16892
rect 9057 16836 9061 16892
rect 8997 16832 9061 16836
rect 9077 16892 9141 16896
rect 9077 16836 9081 16892
rect 9081 16836 9137 16892
rect 9137 16836 9141 16892
rect 9077 16832 9141 16836
rect 9157 16892 9221 16896
rect 9157 16836 9161 16892
rect 9161 16836 9217 16892
rect 9217 16836 9221 16892
rect 9157 16832 9221 16836
rect 24848 16892 24912 16896
rect 24848 16836 24852 16892
rect 24852 16836 24908 16892
rect 24908 16836 24912 16892
rect 24848 16832 24912 16836
rect 24928 16892 24992 16896
rect 24928 16836 24932 16892
rect 24932 16836 24988 16892
rect 24988 16836 24992 16892
rect 24928 16832 24992 16836
rect 25008 16892 25072 16896
rect 25008 16836 25012 16892
rect 25012 16836 25068 16892
rect 25068 16836 25072 16892
rect 25008 16832 25072 16836
rect 25088 16892 25152 16896
rect 25088 16836 25092 16892
rect 25092 16836 25148 16892
rect 25148 16836 25152 16892
rect 25088 16832 25152 16836
rect 40778 16892 40842 16896
rect 40778 16836 40782 16892
rect 40782 16836 40838 16892
rect 40838 16836 40842 16892
rect 40778 16832 40842 16836
rect 40858 16892 40922 16896
rect 40858 16836 40862 16892
rect 40862 16836 40918 16892
rect 40918 16836 40922 16892
rect 40858 16832 40922 16836
rect 40938 16892 41002 16896
rect 40938 16836 40942 16892
rect 40942 16836 40998 16892
rect 40998 16836 41002 16892
rect 40938 16832 41002 16836
rect 41018 16892 41082 16896
rect 41018 16836 41022 16892
rect 41022 16836 41078 16892
rect 41078 16836 41082 16892
rect 41018 16832 41082 16836
rect 16882 16348 16946 16352
rect 16882 16292 16886 16348
rect 16886 16292 16942 16348
rect 16942 16292 16946 16348
rect 16882 16288 16946 16292
rect 16962 16348 17026 16352
rect 16962 16292 16966 16348
rect 16966 16292 17022 16348
rect 17022 16292 17026 16348
rect 16962 16288 17026 16292
rect 17042 16348 17106 16352
rect 17042 16292 17046 16348
rect 17046 16292 17102 16348
rect 17102 16292 17106 16348
rect 17042 16288 17106 16292
rect 17122 16348 17186 16352
rect 17122 16292 17126 16348
rect 17126 16292 17182 16348
rect 17182 16292 17186 16348
rect 17122 16288 17186 16292
rect 32813 16348 32877 16352
rect 32813 16292 32817 16348
rect 32817 16292 32873 16348
rect 32873 16292 32877 16348
rect 32813 16288 32877 16292
rect 32893 16348 32957 16352
rect 32893 16292 32897 16348
rect 32897 16292 32953 16348
rect 32953 16292 32957 16348
rect 32893 16288 32957 16292
rect 32973 16348 33037 16352
rect 32973 16292 32977 16348
rect 32977 16292 33033 16348
rect 33033 16292 33037 16348
rect 32973 16288 33037 16292
rect 33053 16348 33117 16352
rect 33053 16292 33057 16348
rect 33057 16292 33113 16348
rect 33113 16292 33117 16348
rect 33053 16288 33117 16292
rect 8917 15804 8981 15808
rect 8917 15748 8921 15804
rect 8921 15748 8977 15804
rect 8977 15748 8981 15804
rect 8917 15744 8981 15748
rect 8997 15804 9061 15808
rect 8997 15748 9001 15804
rect 9001 15748 9057 15804
rect 9057 15748 9061 15804
rect 8997 15744 9061 15748
rect 9077 15804 9141 15808
rect 9077 15748 9081 15804
rect 9081 15748 9137 15804
rect 9137 15748 9141 15804
rect 9077 15744 9141 15748
rect 9157 15804 9221 15808
rect 9157 15748 9161 15804
rect 9161 15748 9217 15804
rect 9217 15748 9221 15804
rect 9157 15744 9221 15748
rect 24848 15804 24912 15808
rect 24848 15748 24852 15804
rect 24852 15748 24908 15804
rect 24908 15748 24912 15804
rect 24848 15744 24912 15748
rect 24928 15804 24992 15808
rect 24928 15748 24932 15804
rect 24932 15748 24988 15804
rect 24988 15748 24992 15804
rect 24928 15744 24992 15748
rect 25008 15804 25072 15808
rect 25008 15748 25012 15804
rect 25012 15748 25068 15804
rect 25068 15748 25072 15804
rect 25008 15744 25072 15748
rect 25088 15804 25152 15808
rect 25088 15748 25092 15804
rect 25092 15748 25148 15804
rect 25148 15748 25152 15804
rect 25088 15744 25152 15748
rect 40778 15804 40842 15808
rect 40778 15748 40782 15804
rect 40782 15748 40838 15804
rect 40838 15748 40842 15804
rect 40778 15744 40842 15748
rect 40858 15804 40922 15808
rect 40858 15748 40862 15804
rect 40862 15748 40918 15804
rect 40918 15748 40922 15804
rect 40858 15744 40922 15748
rect 40938 15804 41002 15808
rect 40938 15748 40942 15804
rect 40942 15748 40998 15804
rect 40998 15748 41002 15804
rect 40938 15744 41002 15748
rect 41018 15804 41082 15808
rect 41018 15748 41022 15804
rect 41022 15748 41078 15804
rect 41078 15748 41082 15804
rect 41018 15744 41082 15748
rect 16882 15260 16946 15264
rect 16882 15204 16886 15260
rect 16886 15204 16942 15260
rect 16942 15204 16946 15260
rect 16882 15200 16946 15204
rect 16962 15260 17026 15264
rect 16962 15204 16966 15260
rect 16966 15204 17022 15260
rect 17022 15204 17026 15260
rect 16962 15200 17026 15204
rect 17042 15260 17106 15264
rect 17042 15204 17046 15260
rect 17046 15204 17102 15260
rect 17102 15204 17106 15260
rect 17042 15200 17106 15204
rect 17122 15260 17186 15264
rect 17122 15204 17126 15260
rect 17126 15204 17182 15260
rect 17182 15204 17186 15260
rect 17122 15200 17186 15204
rect 32813 15260 32877 15264
rect 32813 15204 32817 15260
rect 32817 15204 32873 15260
rect 32873 15204 32877 15260
rect 32813 15200 32877 15204
rect 32893 15260 32957 15264
rect 32893 15204 32897 15260
rect 32897 15204 32953 15260
rect 32953 15204 32957 15260
rect 32893 15200 32957 15204
rect 32973 15260 33037 15264
rect 32973 15204 32977 15260
rect 32977 15204 33033 15260
rect 33033 15204 33037 15260
rect 32973 15200 33037 15204
rect 33053 15260 33117 15264
rect 33053 15204 33057 15260
rect 33057 15204 33113 15260
rect 33113 15204 33117 15260
rect 33053 15200 33117 15204
rect 8917 14716 8981 14720
rect 8917 14660 8921 14716
rect 8921 14660 8977 14716
rect 8977 14660 8981 14716
rect 8917 14656 8981 14660
rect 8997 14716 9061 14720
rect 8997 14660 9001 14716
rect 9001 14660 9057 14716
rect 9057 14660 9061 14716
rect 8997 14656 9061 14660
rect 9077 14716 9141 14720
rect 9077 14660 9081 14716
rect 9081 14660 9137 14716
rect 9137 14660 9141 14716
rect 9077 14656 9141 14660
rect 9157 14716 9221 14720
rect 9157 14660 9161 14716
rect 9161 14660 9217 14716
rect 9217 14660 9221 14716
rect 9157 14656 9221 14660
rect 24848 14716 24912 14720
rect 24848 14660 24852 14716
rect 24852 14660 24908 14716
rect 24908 14660 24912 14716
rect 24848 14656 24912 14660
rect 24928 14716 24992 14720
rect 24928 14660 24932 14716
rect 24932 14660 24988 14716
rect 24988 14660 24992 14716
rect 24928 14656 24992 14660
rect 25008 14716 25072 14720
rect 25008 14660 25012 14716
rect 25012 14660 25068 14716
rect 25068 14660 25072 14716
rect 25008 14656 25072 14660
rect 25088 14716 25152 14720
rect 25088 14660 25092 14716
rect 25092 14660 25148 14716
rect 25148 14660 25152 14716
rect 25088 14656 25152 14660
rect 40778 14716 40842 14720
rect 40778 14660 40782 14716
rect 40782 14660 40838 14716
rect 40838 14660 40842 14716
rect 40778 14656 40842 14660
rect 40858 14716 40922 14720
rect 40858 14660 40862 14716
rect 40862 14660 40918 14716
rect 40918 14660 40922 14716
rect 40858 14656 40922 14660
rect 40938 14716 41002 14720
rect 40938 14660 40942 14716
rect 40942 14660 40998 14716
rect 40998 14660 41002 14716
rect 40938 14656 41002 14660
rect 41018 14716 41082 14720
rect 41018 14660 41022 14716
rect 41022 14660 41078 14716
rect 41078 14660 41082 14716
rect 41018 14656 41082 14660
rect 16882 14172 16946 14176
rect 16882 14116 16886 14172
rect 16886 14116 16942 14172
rect 16942 14116 16946 14172
rect 16882 14112 16946 14116
rect 16962 14172 17026 14176
rect 16962 14116 16966 14172
rect 16966 14116 17022 14172
rect 17022 14116 17026 14172
rect 16962 14112 17026 14116
rect 17042 14172 17106 14176
rect 17042 14116 17046 14172
rect 17046 14116 17102 14172
rect 17102 14116 17106 14172
rect 17042 14112 17106 14116
rect 17122 14172 17186 14176
rect 17122 14116 17126 14172
rect 17126 14116 17182 14172
rect 17182 14116 17186 14172
rect 17122 14112 17186 14116
rect 32813 14172 32877 14176
rect 32813 14116 32817 14172
rect 32817 14116 32873 14172
rect 32873 14116 32877 14172
rect 32813 14112 32877 14116
rect 32893 14172 32957 14176
rect 32893 14116 32897 14172
rect 32897 14116 32953 14172
rect 32953 14116 32957 14172
rect 32893 14112 32957 14116
rect 32973 14172 33037 14176
rect 32973 14116 32977 14172
rect 32977 14116 33033 14172
rect 33033 14116 33037 14172
rect 32973 14112 33037 14116
rect 33053 14172 33117 14176
rect 33053 14116 33057 14172
rect 33057 14116 33113 14172
rect 33113 14116 33117 14172
rect 33053 14112 33117 14116
rect 8917 13628 8981 13632
rect 8917 13572 8921 13628
rect 8921 13572 8977 13628
rect 8977 13572 8981 13628
rect 8917 13568 8981 13572
rect 8997 13628 9061 13632
rect 8997 13572 9001 13628
rect 9001 13572 9057 13628
rect 9057 13572 9061 13628
rect 8997 13568 9061 13572
rect 9077 13628 9141 13632
rect 9077 13572 9081 13628
rect 9081 13572 9137 13628
rect 9137 13572 9141 13628
rect 9077 13568 9141 13572
rect 9157 13628 9221 13632
rect 9157 13572 9161 13628
rect 9161 13572 9217 13628
rect 9217 13572 9221 13628
rect 9157 13568 9221 13572
rect 24848 13628 24912 13632
rect 24848 13572 24852 13628
rect 24852 13572 24908 13628
rect 24908 13572 24912 13628
rect 24848 13568 24912 13572
rect 24928 13628 24992 13632
rect 24928 13572 24932 13628
rect 24932 13572 24988 13628
rect 24988 13572 24992 13628
rect 24928 13568 24992 13572
rect 25008 13628 25072 13632
rect 25008 13572 25012 13628
rect 25012 13572 25068 13628
rect 25068 13572 25072 13628
rect 25008 13568 25072 13572
rect 25088 13628 25152 13632
rect 25088 13572 25092 13628
rect 25092 13572 25148 13628
rect 25148 13572 25152 13628
rect 25088 13568 25152 13572
rect 40778 13628 40842 13632
rect 40778 13572 40782 13628
rect 40782 13572 40838 13628
rect 40838 13572 40842 13628
rect 40778 13568 40842 13572
rect 40858 13628 40922 13632
rect 40858 13572 40862 13628
rect 40862 13572 40918 13628
rect 40918 13572 40922 13628
rect 40858 13568 40922 13572
rect 40938 13628 41002 13632
rect 40938 13572 40942 13628
rect 40942 13572 40998 13628
rect 40998 13572 41002 13628
rect 40938 13568 41002 13572
rect 41018 13628 41082 13632
rect 41018 13572 41022 13628
rect 41022 13572 41078 13628
rect 41078 13572 41082 13628
rect 41018 13568 41082 13572
rect 16882 13084 16946 13088
rect 16882 13028 16886 13084
rect 16886 13028 16942 13084
rect 16942 13028 16946 13084
rect 16882 13024 16946 13028
rect 16962 13084 17026 13088
rect 16962 13028 16966 13084
rect 16966 13028 17022 13084
rect 17022 13028 17026 13084
rect 16962 13024 17026 13028
rect 17042 13084 17106 13088
rect 17042 13028 17046 13084
rect 17046 13028 17102 13084
rect 17102 13028 17106 13084
rect 17042 13024 17106 13028
rect 17122 13084 17186 13088
rect 17122 13028 17126 13084
rect 17126 13028 17182 13084
rect 17182 13028 17186 13084
rect 17122 13024 17186 13028
rect 32813 13084 32877 13088
rect 32813 13028 32817 13084
rect 32817 13028 32873 13084
rect 32873 13028 32877 13084
rect 32813 13024 32877 13028
rect 32893 13084 32957 13088
rect 32893 13028 32897 13084
rect 32897 13028 32953 13084
rect 32953 13028 32957 13084
rect 32893 13024 32957 13028
rect 32973 13084 33037 13088
rect 32973 13028 32977 13084
rect 32977 13028 33033 13084
rect 33033 13028 33037 13084
rect 32973 13024 33037 13028
rect 33053 13084 33117 13088
rect 33053 13028 33057 13084
rect 33057 13028 33113 13084
rect 33113 13028 33117 13084
rect 33053 13024 33117 13028
rect 8917 12540 8981 12544
rect 8917 12484 8921 12540
rect 8921 12484 8977 12540
rect 8977 12484 8981 12540
rect 8917 12480 8981 12484
rect 8997 12540 9061 12544
rect 8997 12484 9001 12540
rect 9001 12484 9057 12540
rect 9057 12484 9061 12540
rect 8997 12480 9061 12484
rect 9077 12540 9141 12544
rect 9077 12484 9081 12540
rect 9081 12484 9137 12540
rect 9137 12484 9141 12540
rect 9077 12480 9141 12484
rect 9157 12540 9221 12544
rect 9157 12484 9161 12540
rect 9161 12484 9217 12540
rect 9217 12484 9221 12540
rect 9157 12480 9221 12484
rect 24848 12540 24912 12544
rect 24848 12484 24852 12540
rect 24852 12484 24908 12540
rect 24908 12484 24912 12540
rect 24848 12480 24912 12484
rect 24928 12540 24992 12544
rect 24928 12484 24932 12540
rect 24932 12484 24988 12540
rect 24988 12484 24992 12540
rect 24928 12480 24992 12484
rect 25008 12540 25072 12544
rect 25008 12484 25012 12540
rect 25012 12484 25068 12540
rect 25068 12484 25072 12540
rect 25008 12480 25072 12484
rect 25088 12540 25152 12544
rect 25088 12484 25092 12540
rect 25092 12484 25148 12540
rect 25148 12484 25152 12540
rect 25088 12480 25152 12484
rect 40778 12540 40842 12544
rect 40778 12484 40782 12540
rect 40782 12484 40838 12540
rect 40838 12484 40842 12540
rect 40778 12480 40842 12484
rect 40858 12540 40922 12544
rect 40858 12484 40862 12540
rect 40862 12484 40918 12540
rect 40918 12484 40922 12540
rect 40858 12480 40922 12484
rect 40938 12540 41002 12544
rect 40938 12484 40942 12540
rect 40942 12484 40998 12540
rect 40998 12484 41002 12540
rect 40938 12480 41002 12484
rect 41018 12540 41082 12544
rect 41018 12484 41022 12540
rect 41022 12484 41078 12540
rect 41078 12484 41082 12540
rect 41018 12480 41082 12484
rect 16882 11996 16946 12000
rect 16882 11940 16886 11996
rect 16886 11940 16942 11996
rect 16942 11940 16946 11996
rect 16882 11936 16946 11940
rect 16962 11996 17026 12000
rect 16962 11940 16966 11996
rect 16966 11940 17022 11996
rect 17022 11940 17026 11996
rect 16962 11936 17026 11940
rect 17042 11996 17106 12000
rect 17042 11940 17046 11996
rect 17046 11940 17102 11996
rect 17102 11940 17106 11996
rect 17042 11936 17106 11940
rect 17122 11996 17186 12000
rect 17122 11940 17126 11996
rect 17126 11940 17182 11996
rect 17182 11940 17186 11996
rect 17122 11936 17186 11940
rect 32813 11996 32877 12000
rect 32813 11940 32817 11996
rect 32817 11940 32873 11996
rect 32873 11940 32877 11996
rect 32813 11936 32877 11940
rect 32893 11996 32957 12000
rect 32893 11940 32897 11996
rect 32897 11940 32953 11996
rect 32953 11940 32957 11996
rect 32893 11936 32957 11940
rect 32973 11996 33037 12000
rect 32973 11940 32977 11996
rect 32977 11940 33033 11996
rect 33033 11940 33037 11996
rect 32973 11936 33037 11940
rect 33053 11996 33117 12000
rect 33053 11940 33057 11996
rect 33057 11940 33113 11996
rect 33113 11940 33117 11996
rect 33053 11936 33117 11940
rect 8917 11452 8981 11456
rect 8917 11396 8921 11452
rect 8921 11396 8977 11452
rect 8977 11396 8981 11452
rect 8917 11392 8981 11396
rect 8997 11452 9061 11456
rect 8997 11396 9001 11452
rect 9001 11396 9057 11452
rect 9057 11396 9061 11452
rect 8997 11392 9061 11396
rect 9077 11452 9141 11456
rect 9077 11396 9081 11452
rect 9081 11396 9137 11452
rect 9137 11396 9141 11452
rect 9077 11392 9141 11396
rect 9157 11452 9221 11456
rect 9157 11396 9161 11452
rect 9161 11396 9217 11452
rect 9217 11396 9221 11452
rect 9157 11392 9221 11396
rect 24848 11452 24912 11456
rect 24848 11396 24852 11452
rect 24852 11396 24908 11452
rect 24908 11396 24912 11452
rect 24848 11392 24912 11396
rect 24928 11452 24992 11456
rect 24928 11396 24932 11452
rect 24932 11396 24988 11452
rect 24988 11396 24992 11452
rect 24928 11392 24992 11396
rect 25008 11452 25072 11456
rect 25008 11396 25012 11452
rect 25012 11396 25068 11452
rect 25068 11396 25072 11452
rect 25008 11392 25072 11396
rect 25088 11452 25152 11456
rect 25088 11396 25092 11452
rect 25092 11396 25148 11452
rect 25148 11396 25152 11452
rect 25088 11392 25152 11396
rect 40778 11452 40842 11456
rect 40778 11396 40782 11452
rect 40782 11396 40838 11452
rect 40838 11396 40842 11452
rect 40778 11392 40842 11396
rect 40858 11452 40922 11456
rect 40858 11396 40862 11452
rect 40862 11396 40918 11452
rect 40918 11396 40922 11452
rect 40858 11392 40922 11396
rect 40938 11452 41002 11456
rect 40938 11396 40942 11452
rect 40942 11396 40998 11452
rect 40998 11396 41002 11452
rect 40938 11392 41002 11396
rect 41018 11452 41082 11456
rect 41018 11396 41022 11452
rect 41022 11396 41078 11452
rect 41078 11396 41082 11452
rect 41018 11392 41082 11396
rect 16882 10908 16946 10912
rect 16882 10852 16886 10908
rect 16886 10852 16942 10908
rect 16942 10852 16946 10908
rect 16882 10848 16946 10852
rect 16962 10908 17026 10912
rect 16962 10852 16966 10908
rect 16966 10852 17022 10908
rect 17022 10852 17026 10908
rect 16962 10848 17026 10852
rect 17042 10908 17106 10912
rect 17042 10852 17046 10908
rect 17046 10852 17102 10908
rect 17102 10852 17106 10908
rect 17042 10848 17106 10852
rect 17122 10908 17186 10912
rect 17122 10852 17126 10908
rect 17126 10852 17182 10908
rect 17182 10852 17186 10908
rect 17122 10848 17186 10852
rect 32813 10908 32877 10912
rect 32813 10852 32817 10908
rect 32817 10852 32873 10908
rect 32873 10852 32877 10908
rect 32813 10848 32877 10852
rect 32893 10908 32957 10912
rect 32893 10852 32897 10908
rect 32897 10852 32953 10908
rect 32953 10852 32957 10908
rect 32893 10848 32957 10852
rect 32973 10908 33037 10912
rect 32973 10852 32977 10908
rect 32977 10852 33033 10908
rect 33033 10852 33037 10908
rect 32973 10848 33037 10852
rect 33053 10908 33117 10912
rect 33053 10852 33057 10908
rect 33057 10852 33113 10908
rect 33113 10852 33117 10908
rect 33053 10848 33117 10852
rect 8917 10364 8981 10368
rect 8917 10308 8921 10364
rect 8921 10308 8977 10364
rect 8977 10308 8981 10364
rect 8917 10304 8981 10308
rect 8997 10364 9061 10368
rect 8997 10308 9001 10364
rect 9001 10308 9057 10364
rect 9057 10308 9061 10364
rect 8997 10304 9061 10308
rect 9077 10364 9141 10368
rect 9077 10308 9081 10364
rect 9081 10308 9137 10364
rect 9137 10308 9141 10364
rect 9077 10304 9141 10308
rect 9157 10364 9221 10368
rect 9157 10308 9161 10364
rect 9161 10308 9217 10364
rect 9217 10308 9221 10364
rect 9157 10304 9221 10308
rect 24848 10364 24912 10368
rect 24848 10308 24852 10364
rect 24852 10308 24908 10364
rect 24908 10308 24912 10364
rect 24848 10304 24912 10308
rect 24928 10364 24992 10368
rect 24928 10308 24932 10364
rect 24932 10308 24988 10364
rect 24988 10308 24992 10364
rect 24928 10304 24992 10308
rect 25008 10364 25072 10368
rect 25008 10308 25012 10364
rect 25012 10308 25068 10364
rect 25068 10308 25072 10364
rect 25008 10304 25072 10308
rect 25088 10364 25152 10368
rect 25088 10308 25092 10364
rect 25092 10308 25148 10364
rect 25148 10308 25152 10364
rect 25088 10304 25152 10308
rect 40778 10364 40842 10368
rect 40778 10308 40782 10364
rect 40782 10308 40838 10364
rect 40838 10308 40842 10364
rect 40778 10304 40842 10308
rect 40858 10364 40922 10368
rect 40858 10308 40862 10364
rect 40862 10308 40918 10364
rect 40918 10308 40922 10364
rect 40858 10304 40922 10308
rect 40938 10364 41002 10368
rect 40938 10308 40942 10364
rect 40942 10308 40998 10364
rect 40998 10308 41002 10364
rect 40938 10304 41002 10308
rect 41018 10364 41082 10368
rect 41018 10308 41022 10364
rect 41022 10308 41078 10364
rect 41078 10308 41082 10364
rect 41018 10304 41082 10308
rect 16882 9820 16946 9824
rect 16882 9764 16886 9820
rect 16886 9764 16942 9820
rect 16942 9764 16946 9820
rect 16882 9760 16946 9764
rect 16962 9820 17026 9824
rect 16962 9764 16966 9820
rect 16966 9764 17022 9820
rect 17022 9764 17026 9820
rect 16962 9760 17026 9764
rect 17042 9820 17106 9824
rect 17042 9764 17046 9820
rect 17046 9764 17102 9820
rect 17102 9764 17106 9820
rect 17042 9760 17106 9764
rect 17122 9820 17186 9824
rect 17122 9764 17126 9820
rect 17126 9764 17182 9820
rect 17182 9764 17186 9820
rect 17122 9760 17186 9764
rect 32813 9820 32877 9824
rect 32813 9764 32817 9820
rect 32817 9764 32873 9820
rect 32873 9764 32877 9820
rect 32813 9760 32877 9764
rect 32893 9820 32957 9824
rect 32893 9764 32897 9820
rect 32897 9764 32953 9820
rect 32953 9764 32957 9820
rect 32893 9760 32957 9764
rect 32973 9820 33037 9824
rect 32973 9764 32977 9820
rect 32977 9764 33033 9820
rect 33033 9764 33037 9820
rect 32973 9760 33037 9764
rect 33053 9820 33117 9824
rect 33053 9764 33057 9820
rect 33057 9764 33113 9820
rect 33113 9764 33117 9820
rect 33053 9760 33117 9764
rect 8917 9276 8981 9280
rect 8917 9220 8921 9276
rect 8921 9220 8977 9276
rect 8977 9220 8981 9276
rect 8917 9216 8981 9220
rect 8997 9276 9061 9280
rect 8997 9220 9001 9276
rect 9001 9220 9057 9276
rect 9057 9220 9061 9276
rect 8997 9216 9061 9220
rect 9077 9276 9141 9280
rect 9077 9220 9081 9276
rect 9081 9220 9137 9276
rect 9137 9220 9141 9276
rect 9077 9216 9141 9220
rect 9157 9276 9221 9280
rect 9157 9220 9161 9276
rect 9161 9220 9217 9276
rect 9217 9220 9221 9276
rect 9157 9216 9221 9220
rect 24848 9276 24912 9280
rect 24848 9220 24852 9276
rect 24852 9220 24908 9276
rect 24908 9220 24912 9276
rect 24848 9216 24912 9220
rect 24928 9276 24992 9280
rect 24928 9220 24932 9276
rect 24932 9220 24988 9276
rect 24988 9220 24992 9276
rect 24928 9216 24992 9220
rect 25008 9276 25072 9280
rect 25008 9220 25012 9276
rect 25012 9220 25068 9276
rect 25068 9220 25072 9276
rect 25008 9216 25072 9220
rect 25088 9276 25152 9280
rect 25088 9220 25092 9276
rect 25092 9220 25148 9276
rect 25148 9220 25152 9276
rect 25088 9216 25152 9220
rect 40778 9276 40842 9280
rect 40778 9220 40782 9276
rect 40782 9220 40838 9276
rect 40838 9220 40842 9276
rect 40778 9216 40842 9220
rect 40858 9276 40922 9280
rect 40858 9220 40862 9276
rect 40862 9220 40918 9276
rect 40918 9220 40922 9276
rect 40858 9216 40922 9220
rect 40938 9276 41002 9280
rect 40938 9220 40942 9276
rect 40942 9220 40998 9276
rect 40998 9220 41002 9276
rect 40938 9216 41002 9220
rect 41018 9276 41082 9280
rect 41018 9220 41022 9276
rect 41022 9220 41078 9276
rect 41078 9220 41082 9276
rect 41018 9216 41082 9220
rect 16882 8732 16946 8736
rect 16882 8676 16886 8732
rect 16886 8676 16942 8732
rect 16942 8676 16946 8732
rect 16882 8672 16946 8676
rect 16962 8732 17026 8736
rect 16962 8676 16966 8732
rect 16966 8676 17022 8732
rect 17022 8676 17026 8732
rect 16962 8672 17026 8676
rect 17042 8732 17106 8736
rect 17042 8676 17046 8732
rect 17046 8676 17102 8732
rect 17102 8676 17106 8732
rect 17042 8672 17106 8676
rect 17122 8732 17186 8736
rect 17122 8676 17126 8732
rect 17126 8676 17182 8732
rect 17182 8676 17186 8732
rect 17122 8672 17186 8676
rect 32813 8732 32877 8736
rect 32813 8676 32817 8732
rect 32817 8676 32873 8732
rect 32873 8676 32877 8732
rect 32813 8672 32877 8676
rect 32893 8732 32957 8736
rect 32893 8676 32897 8732
rect 32897 8676 32953 8732
rect 32953 8676 32957 8732
rect 32893 8672 32957 8676
rect 32973 8732 33037 8736
rect 32973 8676 32977 8732
rect 32977 8676 33033 8732
rect 33033 8676 33037 8732
rect 32973 8672 33037 8676
rect 33053 8732 33117 8736
rect 33053 8676 33057 8732
rect 33057 8676 33113 8732
rect 33113 8676 33117 8732
rect 33053 8672 33117 8676
rect 8917 8188 8981 8192
rect 8917 8132 8921 8188
rect 8921 8132 8977 8188
rect 8977 8132 8981 8188
rect 8917 8128 8981 8132
rect 8997 8188 9061 8192
rect 8997 8132 9001 8188
rect 9001 8132 9057 8188
rect 9057 8132 9061 8188
rect 8997 8128 9061 8132
rect 9077 8188 9141 8192
rect 9077 8132 9081 8188
rect 9081 8132 9137 8188
rect 9137 8132 9141 8188
rect 9077 8128 9141 8132
rect 9157 8188 9221 8192
rect 9157 8132 9161 8188
rect 9161 8132 9217 8188
rect 9217 8132 9221 8188
rect 9157 8128 9221 8132
rect 24848 8188 24912 8192
rect 24848 8132 24852 8188
rect 24852 8132 24908 8188
rect 24908 8132 24912 8188
rect 24848 8128 24912 8132
rect 24928 8188 24992 8192
rect 24928 8132 24932 8188
rect 24932 8132 24988 8188
rect 24988 8132 24992 8188
rect 24928 8128 24992 8132
rect 25008 8188 25072 8192
rect 25008 8132 25012 8188
rect 25012 8132 25068 8188
rect 25068 8132 25072 8188
rect 25008 8128 25072 8132
rect 25088 8188 25152 8192
rect 25088 8132 25092 8188
rect 25092 8132 25148 8188
rect 25148 8132 25152 8188
rect 25088 8128 25152 8132
rect 40778 8188 40842 8192
rect 40778 8132 40782 8188
rect 40782 8132 40838 8188
rect 40838 8132 40842 8188
rect 40778 8128 40842 8132
rect 40858 8188 40922 8192
rect 40858 8132 40862 8188
rect 40862 8132 40918 8188
rect 40918 8132 40922 8188
rect 40858 8128 40922 8132
rect 40938 8188 41002 8192
rect 40938 8132 40942 8188
rect 40942 8132 40998 8188
rect 40998 8132 41002 8188
rect 40938 8128 41002 8132
rect 41018 8188 41082 8192
rect 41018 8132 41022 8188
rect 41022 8132 41078 8188
rect 41078 8132 41082 8188
rect 41018 8128 41082 8132
rect 16882 7644 16946 7648
rect 16882 7588 16886 7644
rect 16886 7588 16942 7644
rect 16942 7588 16946 7644
rect 16882 7584 16946 7588
rect 16962 7644 17026 7648
rect 16962 7588 16966 7644
rect 16966 7588 17022 7644
rect 17022 7588 17026 7644
rect 16962 7584 17026 7588
rect 17042 7644 17106 7648
rect 17042 7588 17046 7644
rect 17046 7588 17102 7644
rect 17102 7588 17106 7644
rect 17042 7584 17106 7588
rect 17122 7644 17186 7648
rect 17122 7588 17126 7644
rect 17126 7588 17182 7644
rect 17182 7588 17186 7644
rect 17122 7584 17186 7588
rect 32813 7644 32877 7648
rect 32813 7588 32817 7644
rect 32817 7588 32873 7644
rect 32873 7588 32877 7644
rect 32813 7584 32877 7588
rect 32893 7644 32957 7648
rect 32893 7588 32897 7644
rect 32897 7588 32953 7644
rect 32953 7588 32957 7644
rect 32893 7584 32957 7588
rect 32973 7644 33037 7648
rect 32973 7588 32977 7644
rect 32977 7588 33033 7644
rect 33033 7588 33037 7644
rect 32973 7584 33037 7588
rect 33053 7644 33117 7648
rect 33053 7588 33057 7644
rect 33057 7588 33113 7644
rect 33113 7588 33117 7644
rect 33053 7584 33117 7588
rect 8917 7100 8981 7104
rect 8917 7044 8921 7100
rect 8921 7044 8977 7100
rect 8977 7044 8981 7100
rect 8917 7040 8981 7044
rect 8997 7100 9061 7104
rect 8997 7044 9001 7100
rect 9001 7044 9057 7100
rect 9057 7044 9061 7100
rect 8997 7040 9061 7044
rect 9077 7100 9141 7104
rect 9077 7044 9081 7100
rect 9081 7044 9137 7100
rect 9137 7044 9141 7100
rect 9077 7040 9141 7044
rect 9157 7100 9221 7104
rect 9157 7044 9161 7100
rect 9161 7044 9217 7100
rect 9217 7044 9221 7100
rect 9157 7040 9221 7044
rect 24848 7100 24912 7104
rect 24848 7044 24852 7100
rect 24852 7044 24908 7100
rect 24908 7044 24912 7100
rect 24848 7040 24912 7044
rect 24928 7100 24992 7104
rect 24928 7044 24932 7100
rect 24932 7044 24988 7100
rect 24988 7044 24992 7100
rect 24928 7040 24992 7044
rect 25008 7100 25072 7104
rect 25008 7044 25012 7100
rect 25012 7044 25068 7100
rect 25068 7044 25072 7100
rect 25008 7040 25072 7044
rect 25088 7100 25152 7104
rect 25088 7044 25092 7100
rect 25092 7044 25148 7100
rect 25148 7044 25152 7100
rect 25088 7040 25152 7044
rect 40778 7100 40842 7104
rect 40778 7044 40782 7100
rect 40782 7044 40838 7100
rect 40838 7044 40842 7100
rect 40778 7040 40842 7044
rect 40858 7100 40922 7104
rect 40858 7044 40862 7100
rect 40862 7044 40918 7100
rect 40918 7044 40922 7100
rect 40858 7040 40922 7044
rect 40938 7100 41002 7104
rect 40938 7044 40942 7100
rect 40942 7044 40998 7100
rect 40998 7044 41002 7100
rect 40938 7040 41002 7044
rect 41018 7100 41082 7104
rect 41018 7044 41022 7100
rect 41022 7044 41078 7100
rect 41078 7044 41082 7100
rect 41018 7040 41082 7044
rect 16882 6556 16946 6560
rect 16882 6500 16886 6556
rect 16886 6500 16942 6556
rect 16942 6500 16946 6556
rect 16882 6496 16946 6500
rect 16962 6556 17026 6560
rect 16962 6500 16966 6556
rect 16966 6500 17022 6556
rect 17022 6500 17026 6556
rect 16962 6496 17026 6500
rect 17042 6556 17106 6560
rect 17042 6500 17046 6556
rect 17046 6500 17102 6556
rect 17102 6500 17106 6556
rect 17042 6496 17106 6500
rect 17122 6556 17186 6560
rect 17122 6500 17126 6556
rect 17126 6500 17182 6556
rect 17182 6500 17186 6556
rect 17122 6496 17186 6500
rect 32813 6556 32877 6560
rect 32813 6500 32817 6556
rect 32817 6500 32873 6556
rect 32873 6500 32877 6556
rect 32813 6496 32877 6500
rect 32893 6556 32957 6560
rect 32893 6500 32897 6556
rect 32897 6500 32953 6556
rect 32953 6500 32957 6556
rect 32893 6496 32957 6500
rect 32973 6556 33037 6560
rect 32973 6500 32977 6556
rect 32977 6500 33033 6556
rect 33033 6500 33037 6556
rect 32973 6496 33037 6500
rect 33053 6556 33117 6560
rect 33053 6500 33057 6556
rect 33057 6500 33113 6556
rect 33113 6500 33117 6556
rect 33053 6496 33117 6500
rect 8917 6012 8981 6016
rect 8917 5956 8921 6012
rect 8921 5956 8977 6012
rect 8977 5956 8981 6012
rect 8917 5952 8981 5956
rect 8997 6012 9061 6016
rect 8997 5956 9001 6012
rect 9001 5956 9057 6012
rect 9057 5956 9061 6012
rect 8997 5952 9061 5956
rect 9077 6012 9141 6016
rect 9077 5956 9081 6012
rect 9081 5956 9137 6012
rect 9137 5956 9141 6012
rect 9077 5952 9141 5956
rect 9157 6012 9221 6016
rect 9157 5956 9161 6012
rect 9161 5956 9217 6012
rect 9217 5956 9221 6012
rect 9157 5952 9221 5956
rect 24848 6012 24912 6016
rect 24848 5956 24852 6012
rect 24852 5956 24908 6012
rect 24908 5956 24912 6012
rect 24848 5952 24912 5956
rect 24928 6012 24992 6016
rect 24928 5956 24932 6012
rect 24932 5956 24988 6012
rect 24988 5956 24992 6012
rect 24928 5952 24992 5956
rect 25008 6012 25072 6016
rect 25008 5956 25012 6012
rect 25012 5956 25068 6012
rect 25068 5956 25072 6012
rect 25008 5952 25072 5956
rect 25088 6012 25152 6016
rect 25088 5956 25092 6012
rect 25092 5956 25148 6012
rect 25148 5956 25152 6012
rect 25088 5952 25152 5956
rect 40778 6012 40842 6016
rect 40778 5956 40782 6012
rect 40782 5956 40838 6012
rect 40838 5956 40842 6012
rect 40778 5952 40842 5956
rect 40858 6012 40922 6016
rect 40858 5956 40862 6012
rect 40862 5956 40918 6012
rect 40918 5956 40922 6012
rect 40858 5952 40922 5956
rect 40938 6012 41002 6016
rect 40938 5956 40942 6012
rect 40942 5956 40998 6012
rect 40998 5956 41002 6012
rect 40938 5952 41002 5956
rect 41018 6012 41082 6016
rect 41018 5956 41022 6012
rect 41022 5956 41078 6012
rect 41078 5956 41082 6012
rect 41018 5952 41082 5956
rect 16882 5468 16946 5472
rect 16882 5412 16886 5468
rect 16886 5412 16942 5468
rect 16942 5412 16946 5468
rect 16882 5408 16946 5412
rect 16962 5468 17026 5472
rect 16962 5412 16966 5468
rect 16966 5412 17022 5468
rect 17022 5412 17026 5468
rect 16962 5408 17026 5412
rect 17042 5468 17106 5472
rect 17042 5412 17046 5468
rect 17046 5412 17102 5468
rect 17102 5412 17106 5468
rect 17042 5408 17106 5412
rect 17122 5468 17186 5472
rect 17122 5412 17126 5468
rect 17126 5412 17182 5468
rect 17182 5412 17186 5468
rect 17122 5408 17186 5412
rect 32813 5468 32877 5472
rect 32813 5412 32817 5468
rect 32817 5412 32873 5468
rect 32873 5412 32877 5468
rect 32813 5408 32877 5412
rect 32893 5468 32957 5472
rect 32893 5412 32897 5468
rect 32897 5412 32953 5468
rect 32953 5412 32957 5468
rect 32893 5408 32957 5412
rect 32973 5468 33037 5472
rect 32973 5412 32977 5468
rect 32977 5412 33033 5468
rect 33033 5412 33037 5468
rect 32973 5408 33037 5412
rect 33053 5468 33117 5472
rect 33053 5412 33057 5468
rect 33057 5412 33113 5468
rect 33113 5412 33117 5468
rect 33053 5408 33117 5412
rect 8917 4924 8981 4928
rect 8917 4868 8921 4924
rect 8921 4868 8977 4924
rect 8977 4868 8981 4924
rect 8917 4864 8981 4868
rect 8997 4924 9061 4928
rect 8997 4868 9001 4924
rect 9001 4868 9057 4924
rect 9057 4868 9061 4924
rect 8997 4864 9061 4868
rect 9077 4924 9141 4928
rect 9077 4868 9081 4924
rect 9081 4868 9137 4924
rect 9137 4868 9141 4924
rect 9077 4864 9141 4868
rect 9157 4924 9221 4928
rect 9157 4868 9161 4924
rect 9161 4868 9217 4924
rect 9217 4868 9221 4924
rect 9157 4864 9221 4868
rect 24848 4924 24912 4928
rect 24848 4868 24852 4924
rect 24852 4868 24908 4924
rect 24908 4868 24912 4924
rect 24848 4864 24912 4868
rect 24928 4924 24992 4928
rect 24928 4868 24932 4924
rect 24932 4868 24988 4924
rect 24988 4868 24992 4924
rect 24928 4864 24992 4868
rect 25008 4924 25072 4928
rect 25008 4868 25012 4924
rect 25012 4868 25068 4924
rect 25068 4868 25072 4924
rect 25008 4864 25072 4868
rect 25088 4924 25152 4928
rect 25088 4868 25092 4924
rect 25092 4868 25148 4924
rect 25148 4868 25152 4924
rect 25088 4864 25152 4868
rect 40778 4924 40842 4928
rect 40778 4868 40782 4924
rect 40782 4868 40838 4924
rect 40838 4868 40842 4924
rect 40778 4864 40842 4868
rect 40858 4924 40922 4928
rect 40858 4868 40862 4924
rect 40862 4868 40918 4924
rect 40918 4868 40922 4924
rect 40858 4864 40922 4868
rect 40938 4924 41002 4928
rect 40938 4868 40942 4924
rect 40942 4868 40998 4924
rect 40998 4868 41002 4924
rect 40938 4864 41002 4868
rect 41018 4924 41082 4928
rect 41018 4868 41022 4924
rect 41022 4868 41078 4924
rect 41078 4868 41082 4924
rect 41018 4864 41082 4868
rect 16882 4380 16946 4384
rect 16882 4324 16886 4380
rect 16886 4324 16942 4380
rect 16942 4324 16946 4380
rect 16882 4320 16946 4324
rect 16962 4380 17026 4384
rect 16962 4324 16966 4380
rect 16966 4324 17022 4380
rect 17022 4324 17026 4380
rect 16962 4320 17026 4324
rect 17042 4380 17106 4384
rect 17042 4324 17046 4380
rect 17046 4324 17102 4380
rect 17102 4324 17106 4380
rect 17042 4320 17106 4324
rect 17122 4380 17186 4384
rect 17122 4324 17126 4380
rect 17126 4324 17182 4380
rect 17182 4324 17186 4380
rect 17122 4320 17186 4324
rect 32813 4380 32877 4384
rect 32813 4324 32817 4380
rect 32817 4324 32873 4380
rect 32873 4324 32877 4380
rect 32813 4320 32877 4324
rect 32893 4380 32957 4384
rect 32893 4324 32897 4380
rect 32897 4324 32953 4380
rect 32953 4324 32957 4380
rect 32893 4320 32957 4324
rect 32973 4380 33037 4384
rect 32973 4324 32977 4380
rect 32977 4324 33033 4380
rect 33033 4324 33037 4380
rect 32973 4320 33037 4324
rect 33053 4380 33117 4384
rect 33053 4324 33057 4380
rect 33057 4324 33113 4380
rect 33113 4324 33117 4380
rect 33053 4320 33117 4324
rect 8917 3836 8981 3840
rect 8917 3780 8921 3836
rect 8921 3780 8977 3836
rect 8977 3780 8981 3836
rect 8917 3776 8981 3780
rect 8997 3836 9061 3840
rect 8997 3780 9001 3836
rect 9001 3780 9057 3836
rect 9057 3780 9061 3836
rect 8997 3776 9061 3780
rect 9077 3836 9141 3840
rect 9077 3780 9081 3836
rect 9081 3780 9137 3836
rect 9137 3780 9141 3836
rect 9077 3776 9141 3780
rect 9157 3836 9221 3840
rect 9157 3780 9161 3836
rect 9161 3780 9217 3836
rect 9217 3780 9221 3836
rect 9157 3776 9221 3780
rect 24848 3836 24912 3840
rect 24848 3780 24852 3836
rect 24852 3780 24908 3836
rect 24908 3780 24912 3836
rect 24848 3776 24912 3780
rect 24928 3836 24992 3840
rect 24928 3780 24932 3836
rect 24932 3780 24988 3836
rect 24988 3780 24992 3836
rect 24928 3776 24992 3780
rect 25008 3836 25072 3840
rect 25008 3780 25012 3836
rect 25012 3780 25068 3836
rect 25068 3780 25072 3836
rect 25008 3776 25072 3780
rect 25088 3836 25152 3840
rect 25088 3780 25092 3836
rect 25092 3780 25148 3836
rect 25148 3780 25152 3836
rect 25088 3776 25152 3780
rect 40778 3836 40842 3840
rect 40778 3780 40782 3836
rect 40782 3780 40838 3836
rect 40838 3780 40842 3836
rect 40778 3776 40842 3780
rect 40858 3836 40922 3840
rect 40858 3780 40862 3836
rect 40862 3780 40918 3836
rect 40918 3780 40922 3836
rect 40858 3776 40922 3780
rect 40938 3836 41002 3840
rect 40938 3780 40942 3836
rect 40942 3780 40998 3836
rect 40998 3780 41002 3836
rect 40938 3776 41002 3780
rect 41018 3836 41082 3840
rect 41018 3780 41022 3836
rect 41022 3780 41078 3836
rect 41078 3780 41082 3836
rect 41018 3776 41082 3780
rect 16882 3292 16946 3296
rect 16882 3236 16886 3292
rect 16886 3236 16942 3292
rect 16942 3236 16946 3292
rect 16882 3232 16946 3236
rect 16962 3292 17026 3296
rect 16962 3236 16966 3292
rect 16966 3236 17022 3292
rect 17022 3236 17026 3292
rect 16962 3232 17026 3236
rect 17042 3292 17106 3296
rect 17042 3236 17046 3292
rect 17046 3236 17102 3292
rect 17102 3236 17106 3292
rect 17042 3232 17106 3236
rect 17122 3292 17186 3296
rect 17122 3236 17126 3292
rect 17126 3236 17182 3292
rect 17182 3236 17186 3292
rect 17122 3232 17186 3236
rect 32813 3292 32877 3296
rect 32813 3236 32817 3292
rect 32817 3236 32873 3292
rect 32873 3236 32877 3292
rect 32813 3232 32877 3236
rect 32893 3292 32957 3296
rect 32893 3236 32897 3292
rect 32897 3236 32953 3292
rect 32953 3236 32957 3292
rect 32893 3232 32957 3236
rect 32973 3292 33037 3296
rect 32973 3236 32977 3292
rect 32977 3236 33033 3292
rect 33033 3236 33037 3292
rect 32973 3232 33037 3236
rect 33053 3292 33117 3296
rect 33053 3236 33057 3292
rect 33057 3236 33113 3292
rect 33113 3236 33117 3292
rect 33053 3232 33117 3236
rect 8917 2748 8981 2752
rect 8917 2692 8921 2748
rect 8921 2692 8977 2748
rect 8977 2692 8981 2748
rect 8917 2688 8981 2692
rect 8997 2748 9061 2752
rect 8997 2692 9001 2748
rect 9001 2692 9057 2748
rect 9057 2692 9061 2748
rect 8997 2688 9061 2692
rect 9077 2748 9141 2752
rect 9077 2692 9081 2748
rect 9081 2692 9137 2748
rect 9137 2692 9141 2748
rect 9077 2688 9141 2692
rect 9157 2748 9221 2752
rect 9157 2692 9161 2748
rect 9161 2692 9217 2748
rect 9217 2692 9221 2748
rect 9157 2688 9221 2692
rect 24848 2748 24912 2752
rect 24848 2692 24852 2748
rect 24852 2692 24908 2748
rect 24908 2692 24912 2748
rect 24848 2688 24912 2692
rect 24928 2748 24992 2752
rect 24928 2692 24932 2748
rect 24932 2692 24988 2748
rect 24988 2692 24992 2748
rect 24928 2688 24992 2692
rect 25008 2748 25072 2752
rect 25008 2692 25012 2748
rect 25012 2692 25068 2748
rect 25068 2692 25072 2748
rect 25008 2688 25072 2692
rect 25088 2748 25152 2752
rect 25088 2692 25092 2748
rect 25092 2692 25148 2748
rect 25148 2692 25152 2748
rect 25088 2688 25152 2692
rect 40778 2748 40842 2752
rect 40778 2692 40782 2748
rect 40782 2692 40838 2748
rect 40838 2692 40842 2748
rect 40778 2688 40842 2692
rect 40858 2748 40922 2752
rect 40858 2692 40862 2748
rect 40862 2692 40918 2748
rect 40918 2692 40922 2748
rect 40858 2688 40922 2692
rect 40938 2748 41002 2752
rect 40938 2692 40942 2748
rect 40942 2692 40998 2748
rect 40998 2692 41002 2748
rect 40938 2688 41002 2692
rect 41018 2748 41082 2752
rect 41018 2692 41022 2748
rect 41022 2692 41078 2748
rect 41078 2692 41082 2748
rect 41018 2688 41082 2692
rect 16882 2204 16946 2208
rect 16882 2148 16886 2204
rect 16886 2148 16942 2204
rect 16942 2148 16946 2204
rect 16882 2144 16946 2148
rect 16962 2204 17026 2208
rect 16962 2148 16966 2204
rect 16966 2148 17022 2204
rect 17022 2148 17026 2204
rect 16962 2144 17026 2148
rect 17042 2204 17106 2208
rect 17042 2148 17046 2204
rect 17046 2148 17102 2204
rect 17102 2148 17106 2204
rect 17042 2144 17106 2148
rect 17122 2204 17186 2208
rect 17122 2148 17126 2204
rect 17126 2148 17182 2204
rect 17182 2148 17186 2204
rect 17122 2144 17186 2148
rect 32813 2204 32877 2208
rect 32813 2148 32817 2204
rect 32817 2148 32873 2204
rect 32873 2148 32877 2204
rect 32813 2144 32877 2148
rect 32893 2204 32957 2208
rect 32893 2148 32897 2204
rect 32897 2148 32953 2204
rect 32953 2148 32957 2204
rect 32893 2144 32957 2148
rect 32973 2204 33037 2208
rect 32973 2148 32977 2204
rect 32977 2148 33033 2204
rect 33033 2148 33037 2204
rect 32973 2144 33037 2148
rect 33053 2204 33117 2208
rect 33053 2148 33057 2204
rect 33057 2148 33113 2204
rect 33113 2148 33117 2204
rect 33053 2144 33117 2148
<< metal4 >>
rect 8909 16896 9230 17456
rect 8909 16832 8917 16896
rect 8981 16832 8997 16896
rect 9061 16832 9077 16896
rect 9141 16832 9157 16896
rect 9221 16832 9230 16896
rect 8909 15808 9230 16832
rect 8909 15744 8917 15808
rect 8981 15744 8997 15808
rect 9061 15744 9077 15808
rect 9141 15744 9157 15808
rect 9221 15744 9230 15808
rect 8909 14720 9230 15744
rect 8909 14656 8917 14720
rect 8981 14656 8997 14720
rect 9061 14656 9077 14720
rect 9141 14656 9157 14720
rect 9221 14656 9230 14720
rect 8909 13632 9230 14656
rect 8909 13568 8917 13632
rect 8981 13568 8997 13632
rect 9061 13568 9077 13632
rect 9141 13568 9157 13632
rect 9221 13568 9230 13632
rect 8909 12544 9230 13568
rect 8909 12480 8917 12544
rect 8981 12480 8997 12544
rect 9061 12480 9077 12544
rect 9141 12480 9157 12544
rect 9221 12480 9230 12544
rect 8909 11456 9230 12480
rect 8909 11392 8917 11456
rect 8981 11392 8997 11456
rect 9061 11392 9077 11456
rect 9141 11392 9157 11456
rect 9221 11392 9230 11456
rect 8909 10368 9230 11392
rect 8909 10304 8917 10368
rect 8981 10304 8997 10368
rect 9061 10304 9077 10368
rect 9141 10304 9157 10368
rect 9221 10304 9230 10368
rect 8909 9280 9230 10304
rect 8909 9216 8917 9280
rect 8981 9216 8997 9280
rect 9061 9216 9077 9280
rect 9141 9216 9157 9280
rect 9221 9216 9230 9280
rect 8909 8192 9230 9216
rect 8909 8128 8917 8192
rect 8981 8128 8997 8192
rect 9061 8128 9077 8192
rect 9141 8128 9157 8192
rect 9221 8128 9230 8192
rect 8909 7104 9230 8128
rect 8909 7040 8917 7104
rect 8981 7040 8997 7104
rect 9061 7040 9077 7104
rect 9141 7040 9157 7104
rect 9221 7040 9230 7104
rect 8909 6016 9230 7040
rect 8909 5952 8917 6016
rect 8981 5952 8997 6016
rect 9061 5952 9077 6016
rect 9141 5952 9157 6016
rect 9221 5952 9230 6016
rect 8909 4928 9230 5952
rect 8909 4864 8917 4928
rect 8981 4864 8997 4928
rect 9061 4864 9077 4928
rect 9141 4864 9157 4928
rect 9221 4864 9230 4928
rect 8909 3840 9230 4864
rect 8909 3776 8917 3840
rect 8981 3776 8997 3840
rect 9061 3776 9077 3840
rect 9141 3776 9157 3840
rect 9221 3776 9230 3840
rect 8909 2752 9230 3776
rect 8909 2688 8917 2752
rect 8981 2688 8997 2752
rect 9061 2688 9077 2752
rect 9141 2688 9157 2752
rect 9221 2688 9230 2752
rect 8909 2128 9230 2688
rect 16874 17440 17194 17456
rect 16874 17376 16882 17440
rect 16946 17376 16962 17440
rect 17026 17376 17042 17440
rect 17106 17376 17122 17440
rect 17186 17376 17194 17440
rect 16874 16352 17194 17376
rect 16874 16288 16882 16352
rect 16946 16288 16962 16352
rect 17026 16288 17042 16352
rect 17106 16288 17122 16352
rect 17186 16288 17194 16352
rect 16874 15264 17194 16288
rect 16874 15200 16882 15264
rect 16946 15200 16962 15264
rect 17026 15200 17042 15264
rect 17106 15200 17122 15264
rect 17186 15200 17194 15264
rect 16874 14176 17194 15200
rect 16874 14112 16882 14176
rect 16946 14112 16962 14176
rect 17026 14112 17042 14176
rect 17106 14112 17122 14176
rect 17186 14112 17194 14176
rect 16874 13088 17194 14112
rect 16874 13024 16882 13088
rect 16946 13024 16962 13088
rect 17026 13024 17042 13088
rect 17106 13024 17122 13088
rect 17186 13024 17194 13088
rect 16874 12000 17194 13024
rect 16874 11936 16882 12000
rect 16946 11936 16962 12000
rect 17026 11936 17042 12000
rect 17106 11936 17122 12000
rect 17186 11936 17194 12000
rect 16874 10912 17194 11936
rect 16874 10848 16882 10912
rect 16946 10848 16962 10912
rect 17026 10848 17042 10912
rect 17106 10848 17122 10912
rect 17186 10848 17194 10912
rect 16874 9824 17194 10848
rect 16874 9760 16882 9824
rect 16946 9760 16962 9824
rect 17026 9760 17042 9824
rect 17106 9760 17122 9824
rect 17186 9760 17194 9824
rect 16874 8736 17194 9760
rect 16874 8672 16882 8736
rect 16946 8672 16962 8736
rect 17026 8672 17042 8736
rect 17106 8672 17122 8736
rect 17186 8672 17194 8736
rect 16874 7648 17194 8672
rect 16874 7584 16882 7648
rect 16946 7584 16962 7648
rect 17026 7584 17042 7648
rect 17106 7584 17122 7648
rect 17186 7584 17194 7648
rect 16874 6560 17194 7584
rect 16874 6496 16882 6560
rect 16946 6496 16962 6560
rect 17026 6496 17042 6560
rect 17106 6496 17122 6560
rect 17186 6496 17194 6560
rect 16874 5472 17194 6496
rect 16874 5408 16882 5472
rect 16946 5408 16962 5472
rect 17026 5408 17042 5472
rect 17106 5408 17122 5472
rect 17186 5408 17194 5472
rect 16874 4384 17194 5408
rect 16874 4320 16882 4384
rect 16946 4320 16962 4384
rect 17026 4320 17042 4384
rect 17106 4320 17122 4384
rect 17186 4320 17194 4384
rect 16874 3296 17194 4320
rect 16874 3232 16882 3296
rect 16946 3232 16962 3296
rect 17026 3232 17042 3296
rect 17106 3232 17122 3296
rect 17186 3232 17194 3296
rect 16874 2208 17194 3232
rect 16874 2144 16882 2208
rect 16946 2144 16962 2208
rect 17026 2144 17042 2208
rect 17106 2144 17122 2208
rect 17186 2144 17194 2208
rect 16874 2128 17194 2144
rect 24840 16896 25160 17456
rect 24840 16832 24848 16896
rect 24912 16832 24928 16896
rect 24992 16832 25008 16896
rect 25072 16832 25088 16896
rect 25152 16832 25160 16896
rect 24840 15808 25160 16832
rect 24840 15744 24848 15808
rect 24912 15744 24928 15808
rect 24992 15744 25008 15808
rect 25072 15744 25088 15808
rect 25152 15744 25160 15808
rect 24840 14720 25160 15744
rect 24840 14656 24848 14720
rect 24912 14656 24928 14720
rect 24992 14656 25008 14720
rect 25072 14656 25088 14720
rect 25152 14656 25160 14720
rect 24840 13632 25160 14656
rect 24840 13568 24848 13632
rect 24912 13568 24928 13632
rect 24992 13568 25008 13632
rect 25072 13568 25088 13632
rect 25152 13568 25160 13632
rect 24840 12544 25160 13568
rect 24840 12480 24848 12544
rect 24912 12480 24928 12544
rect 24992 12480 25008 12544
rect 25072 12480 25088 12544
rect 25152 12480 25160 12544
rect 24840 11456 25160 12480
rect 24840 11392 24848 11456
rect 24912 11392 24928 11456
rect 24992 11392 25008 11456
rect 25072 11392 25088 11456
rect 25152 11392 25160 11456
rect 24840 10368 25160 11392
rect 24840 10304 24848 10368
rect 24912 10304 24928 10368
rect 24992 10304 25008 10368
rect 25072 10304 25088 10368
rect 25152 10304 25160 10368
rect 24840 9280 25160 10304
rect 24840 9216 24848 9280
rect 24912 9216 24928 9280
rect 24992 9216 25008 9280
rect 25072 9216 25088 9280
rect 25152 9216 25160 9280
rect 24840 8192 25160 9216
rect 24840 8128 24848 8192
rect 24912 8128 24928 8192
rect 24992 8128 25008 8192
rect 25072 8128 25088 8192
rect 25152 8128 25160 8192
rect 24840 7104 25160 8128
rect 24840 7040 24848 7104
rect 24912 7040 24928 7104
rect 24992 7040 25008 7104
rect 25072 7040 25088 7104
rect 25152 7040 25160 7104
rect 24840 6016 25160 7040
rect 24840 5952 24848 6016
rect 24912 5952 24928 6016
rect 24992 5952 25008 6016
rect 25072 5952 25088 6016
rect 25152 5952 25160 6016
rect 24840 4928 25160 5952
rect 24840 4864 24848 4928
rect 24912 4864 24928 4928
rect 24992 4864 25008 4928
rect 25072 4864 25088 4928
rect 25152 4864 25160 4928
rect 24840 3840 25160 4864
rect 24840 3776 24848 3840
rect 24912 3776 24928 3840
rect 24992 3776 25008 3840
rect 25072 3776 25088 3840
rect 25152 3776 25160 3840
rect 24840 2752 25160 3776
rect 24840 2688 24848 2752
rect 24912 2688 24928 2752
rect 24992 2688 25008 2752
rect 25072 2688 25088 2752
rect 25152 2688 25160 2752
rect 24840 2128 25160 2688
rect 32805 17440 33125 17456
rect 32805 17376 32813 17440
rect 32877 17376 32893 17440
rect 32957 17376 32973 17440
rect 33037 17376 33053 17440
rect 33117 17376 33125 17440
rect 32805 16352 33125 17376
rect 32805 16288 32813 16352
rect 32877 16288 32893 16352
rect 32957 16288 32973 16352
rect 33037 16288 33053 16352
rect 33117 16288 33125 16352
rect 32805 15264 33125 16288
rect 32805 15200 32813 15264
rect 32877 15200 32893 15264
rect 32957 15200 32973 15264
rect 33037 15200 33053 15264
rect 33117 15200 33125 15264
rect 32805 14176 33125 15200
rect 32805 14112 32813 14176
rect 32877 14112 32893 14176
rect 32957 14112 32973 14176
rect 33037 14112 33053 14176
rect 33117 14112 33125 14176
rect 32805 13088 33125 14112
rect 32805 13024 32813 13088
rect 32877 13024 32893 13088
rect 32957 13024 32973 13088
rect 33037 13024 33053 13088
rect 33117 13024 33125 13088
rect 32805 12000 33125 13024
rect 32805 11936 32813 12000
rect 32877 11936 32893 12000
rect 32957 11936 32973 12000
rect 33037 11936 33053 12000
rect 33117 11936 33125 12000
rect 32805 10912 33125 11936
rect 32805 10848 32813 10912
rect 32877 10848 32893 10912
rect 32957 10848 32973 10912
rect 33037 10848 33053 10912
rect 33117 10848 33125 10912
rect 32805 9824 33125 10848
rect 32805 9760 32813 9824
rect 32877 9760 32893 9824
rect 32957 9760 32973 9824
rect 33037 9760 33053 9824
rect 33117 9760 33125 9824
rect 32805 8736 33125 9760
rect 32805 8672 32813 8736
rect 32877 8672 32893 8736
rect 32957 8672 32973 8736
rect 33037 8672 33053 8736
rect 33117 8672 33125 8736
rect 32805 7648 33125 8672
rect 32805 7584 32813 7648
rect 32877 7584 32893 7648
rect 32957 7584 32973 7648
rect 33037 7584 33053 7648
rect 33117 7584 33125 7648
rect 32805 6560 33125 7584
rect 32805 6496 32813 6560
rect 32877 6496 32893 6560
rect 32957 6496 32973 6560
rect 33037 6496 33053 6560
rect 33117 6496 33125 6560
rect 32805 5472 33125 6496
rect 32805 5408 32813 5472
rect 32877 5408 32893 5472
rect 32957 5408 32973 5472
rect 33037 5408 33053 5472
rect 33117 5408 33125 5472
rect 32805 4384 33125 5408
rect 32805 4320 32813 4384
rect 32877 4320 32893 4384
rect 32957 4320 32973 4384
rect 33037 4320 33053 4384
rect 33117 4320 33125 4384
rect 32805 3296 33125 4320
rect 32805 3232 32813 3296
rect 32877 3232 32893 3296
rect 32957 3232 32973 3296
rect 33037 3232 33053 3296
rect 33117 3232 33125 3296
rect 32805 2208 33125 3232
rect 32805 2144 32813 2208
rect 32877 2144 32893 2208
rect 32957 2144 32973 2208
rect 33037 2144 33053 2208
rect 33117 2144 33125 2208
rect 32805 2128 33125 2144
rect 40770 16896 41091 17456
rect 40770 16832 40778 16896
rect 40842 16832 40858 16896
rect 40922 16832 40938 16896
rect 41002 16832 41018 16896
rect 41082 16832 41091 16896
rect 40770 15808 41091 16832
rect 40770 15744 40778 15808
rect 40842 15744 40858 15808
rect 40922 15744 40938 15808
rect 41002 15744 41018 15808
rect 41082 15744 41091 15808
rect 40770 14720 41091 15744
rect 40770 14656 40778 14720
rect 40842 14656 40858 14720
rect 40922 14656 40938 14720
rect 41002 14656 41018 14720
rect 41082 14656 41091 14720
rect 40770 13632 41091 14656
rect 40770 13568 40778 13632
rect 40842 13568 40858 13632
rect 40922 13568 40938 13632
rect 41002 13568 41018 13632
rect 41082 13568 41091 13632
rect 40770 12544 41091 13568
rect 40770 12480 40778 12544
rect 40842 12480 40858 12544
rect 40922 12480 40938 12544
rect 41002 12480 41018 12544
rect 41082 12480 41091 12544
rect 40770 11456 41091 12480
rect 40770 11392 40778 11456
rect 40842 11392 40858 11456
rect 40922 11392 40938 11456
rect 41002 11392 41018 11456
rect 41082 11392 41091 11456
rect 40770 10368 41091 11392
rect 40770 10304 40778 10368
rect 40842 10304 40858 10368
rect 40922 10304 40938 10368
rect 41002 10304 41018 10368
rect 41082 10304 41091 10368
rect 40770 9280 41091 10304
rect 40770 9216 40778 9280
rect 40842 9216 40858 9280
rect 40922 9216 40938 9280
rect 41002 9216 41018 9280
rect 41082 9216 41091 9280
rect 40770 8192 41091 9216
rect 40770 8128 40778 8192
rect 40842 8128 40858 8192
rect 40922 8128 40938 8192
rect 41002 8128 41018 8192
rect 41082 8128 41091 8192
rect 40770 7104 41091 8128
rect 40770 7040 40778 7104
rect 40842 7040 40858 7104
rect 40922 7040 40938 7104
rect 41002 7040 41018 7104
rect 41082 7040 41091 7104
rect 40770 6016 41091 7040
rect 40770 5952 40778 6016
rect 40842 5952 40858 6016
rect 40922 5952 40938 6016
rect 41002 5952 41018 6016
rect 41082 5952 41091 6016
rect 40770 4928 41091 5952
rect 40770 4864 40778 4928
rect 40842 4864 40858 4928
rect 40922 4864 40938 4928
rect 41002 4864 41018 4928
rect 41082 4864 41091 4928
rect 40770 3840 41091 4864
rect 40770 3776 40778 3840
rect 40842 3776 40858 3840
rect 40922 3776 40938 3840
rect 41002 3776 41018 3840
rect 41082 3776 41091 3840
rect 40770 2752 41091 3776
rect 40770 2688 40778 2752
rect 40842 2688 40858 2752
rect 40922 2688 40938 2752
rect 41002 2688 41018 2752
rect 41082 2688 41091 2752
rect 40770 2128 41091 2688
use sky130_fd_sc_hd__decap_8  FILLER_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 1380 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 2116 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 2668 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24
timestamp 1644511149
transform 1 0 3312 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 5704 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_78
timestamp 1644511149
transform 1 0 8280 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_106
timestamp 1644511149
transform 1 0 10856 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_113 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 11500 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_136
timestamp 1644511149
transform 1 0 13616 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_141 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 14076 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_163
timestamp 1644511149
transform 1 0 16100 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_167
timestamp 1644511149
transform 1 0 16468 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_190
timestamp 1644511149
transform 1 0 18584 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_197
timestamp 1644511149
transform 1 0 19228 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_220
timestamp 1644511149
transform 1 0 21344 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_225
timestamp 1644511149
transform 1 0 21804 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_248
timestamp 1644511149
transform 1 0 23920 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_253
timestamp 1644511149
transform 1 0 24380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_276
timestamp 1644511149
transform 1 0 26496 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_281
timestamp 1644511149
transform 1 0 26956 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_304
timestamp 1644511149
transform 1 0 29072 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_312 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 29808 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_324
timestamp 1644511149
transform 1 0 30912 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_329
timestamp 1644511149
transform 1 0 31372 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_335
timestamp 1644511149
transform 1 0 31924 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_358
timestamp 1644511149
transform 1 0 34040 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_386
timestamp 1644511149
transform 1 0 36616 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_414
timestamp 1644511149
transform 1 0 39192 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_421
timestamp 1644511149
transform 1 0 39836 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_443
timestamp 1644511149
transform 1 0 41860 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_447
timestamp 1644511149
transform 1 0 42228 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_449
timestamp 1644511149
transform 1 0 42412 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_472
timestamp 1644511149
transform 1 0 44528 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_477
timestamp 1644511149
transform 1 0 44988 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_500
timestamp 1644511149
transform 1 0 47104 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_508
timestamp 1644511149
transform 1 0 47840 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_3
timestamp 1644511149
transform 1 0 1380 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_7
timestamp 1644511149
transform 1 0 1748 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_32
timestamp 1644511149
transform 1 0 4048 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_39
timestamp 1644511149
transform 1 0 4692 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_47
timestamp 1644511149
transform 1 0 5428 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_52
timestamp 1644511149
transform 1 0 5888 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_57
timestamp 1644511149
transform 1 0 6348 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_64
timestamp 1644511149
transform 1 0 6992 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_73
timestamp 1644511149
transform 1 0 7820 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_80
timestamp 1644511149
transform 1 0 8464 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_105
timestamp 1644511149
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 1644511149
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_113
timestamp 1644511149
transform 1 0 11500 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_118
timestamp 1644511149
transform 1 0 11960 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_122
timestamp 1644511149
transform 1 0 12328 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_126
timestamp 1644511149
transform 1 0 12696 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_134
timestamp 1644511149
transform 1 0 13432 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_157
timestamp 1644511149
transform 1 0 15548 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_164
timestamp 1644511149
transform 1 0 16192 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_172
timestamp 1644511149
transform 1 0 16928 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_181
timestamp 1644511149
transform 1 0 17756 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_206
timestamp 1644511149
transform 1 0 20056 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_213
timestamp 1644511149
transform 1 0 20700 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_220
timestamp 1644511149
transform 1 0 21344 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_225
timestamp 1644511149
transform 1 0 21804 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_234
timestamp 1644511149
transform 1 0 22632 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_241
timestamp 1644511149
transform 1 0 23276 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_247
timestamp 1644511149
transform 1 0 23828 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_269
timestamp 1644511149
transform 1 0 25852 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_276
timestamp 1644511149
transform 1 0 26496 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_284
timestamp 1644511149
transform 1 0 27232 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_292
timestamp 1644511149
transform 1 0 27968 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_297
timestamp 1644511149
transform 1 0 28428 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_322
timestamp 1644511149
transform 1 0 30728 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_328
timestamp 1644511149
transform 1 0 31280 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_332
timestamp 1644511149
transform 1 0 31648 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_358
timestamp 1644511149
transform 1 0 34040 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_366
timestamp 1644511149
transform 1 0 34776 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_388
timestamp 1644511149
transform 1 0 36800 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_396
timestamp 1644511149
transform 1 0 37536 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_404
timestamp 1644511149
transform 1 0 38272 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_409
timestamp 1644511149
transform 1 0 38732 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_434
timestamp 1644511149
transform 1 0 41032 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_444
timestamp 1644511149
transform 1 0 41952 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_449
timestamp 1644511149
transform 1 0 42412 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_453
timestamp 1644511149
transform 1 0 42780 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_478
timestamp 1644511149
transform 1 0 45080 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_485
timestamp 1644511149
transform 1 0 45724 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_493
timestamp 1644511149
transform 1 0 46460 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_497
timestamp 1644511149
transform 1 0 46828 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_503
timestamp 1644511149
transform 1 0 47380 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_508
timestamp 1644511149
transform 1 0 47840 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_2_24
timestamp 1644511149
transform 1 0 3312 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_32
timestamp 1644511149
transform 1 0 4048 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_39
timestamp 1644511149
transform 1 0 4692 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_46
timestamp 1644511149
transform 1 0 5336 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_71
timestamp 1644511149
transform 1 0 7636 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_80
timestamp 1644511149
transform 1 0 8464 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_85
timestamp 1644511149
transform 1 0 8924 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_2_108
timestamp 1644511149
transform 1 0 11040 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_135
timestamp 1644511149
transform 1 0 13524 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 1644511149
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_141
timestamp 1644511149
transform 1 0 14076 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_146
timestamp 1644511149
transform 1 0 14536 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_153
timestamp 1644511149
transform 1 0 15180 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_180
timestamp 1644511149
transform 1 0 17664 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_184
timestamp 1644511149
transform 1 0 18032 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_188
timestamp 1644511149
transform 1 0 18400 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_2_200
timestamp 1644511149
transform 1 0 19504 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_207
timestamp 1644511149
transform 1 0 20148 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_219
timestamp 1644511149
transform 1 0 21252 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_231
timestamp 1644511149
transform 1 0 22356 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_2_243
timestamp 1644511149
transform 1 0 23460 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_248
timestamp 1644511149
transform 1 0 23920 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_2_253
timestamp 1644511149
transform 1 0 24380 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_259
timestamp 1644511149
transform 1 0 24932 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_266
timestamp 1644511149
transform 1 0 25576 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_272
timestamp 1644511149
transform 1 0 26128 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_276
timestamp 1644511149
transform 1 0 26496 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_301
timestamp 1644511149
transform 1 0 28796 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_307
timestamp 1644511149
transform 1 0 29348 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_312
timestamp 1644511149
transform 1 0 29808 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_2_324
timestamp 1644511149
transform 1 0 30912 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_2_329
timestamp 1644511149
transform 1 0 31372 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_335
timestamp 1644511149
transform 1 0 31924 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_357
timestamp 1644511149
transform 1 0 33948 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_363
timestamp 1644511149
transform 1 0 34500 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_368
timestamp 1644511149
transform 1 0 34960 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_376
timestamp 1644511149
transform 1 0 35696 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_399
timestamp 1644511149
transform 1 0 37812 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_406
timestamp 1644511149
transform 1 0 38456 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_412
timestamp 1644511149
transform 1 0 39008 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_416
timestamp 1644511149
transform 1 0 39376 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_424
timestamp 1644511149
transform 1 0 40112 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_428
timestamp 1644511149
transform 1 0 40480 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_445
timestamp 1644511149
transform 1 0 42044 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_470
timestamp 1644511149
transform 1 0 44344 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_480
timestamp 1644511149
transform 1 0 45264 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_487
timestamp 1644511149
transform 1 0 45908 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_512
timestamp 1644511149
transform 1 0 48208 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_3
timestamp 1644511149
transform 1 0 1380 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_9
timestamp 1644511149
transform 1 0 1932 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_13
timestamp 1644511149
transform 1 0 2300 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_38
timestamp 1644511149
transform 1 0 4600 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_45
timestamp 1644511149
transform 1 0 5244 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_52
timestamp 1644511149
transform 1 0 5888 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_78
timestamp 1644511149
transform 1 0 8280 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_86
timestamp 1644511149
transform 1 0 9016 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_91
timestamp 1644511149
transform 1 0 9476 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_98
timestamp 1644511149
transform 1 0 10120 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_110
timestamp 1644511149
transform 1 0 11224 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_113
timestamp 1644511149
transform 1 0 11500 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_118
timestamp 1644511149
transform 1 0 11960 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_125
timestamp 1644511149
transform 1 0 12604 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_3_133
timestamp 1644511149
transform 1 0 13340 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_139
timestamp 1644511149
transform 1 0 13892 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_146
timestamp 1644511149
transform 1 0 14536 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_158
timestamp 1644511149
transform 1 0 15640 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_163
timestamp 1644511149
transform 1 0 16100 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1644511149
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_169
timestamp 1644511149
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_181
timestamp 1644511149
transform 1 0 17756 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_185
timestamp 1644511149
transform 1 0 18124 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_207
timestamp 1644511149
transform 1 0 20148 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_219
timestamp 1644511149
transform 1 0 21252 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_223
timestamp 1644511149
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_225
timestamp 1644511149
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_237
timestamp 1644511149
transform 1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_249
timestamp 1644511149
transform 1 0 24012 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_261
timestamp 1644511149
transform 1 0 25116 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_273
timestamp 1644511149
transform 1 0 26220 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_279
timestamp 1644511149
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_287
timestamp 1644511149
transform 1 0 27508 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_312
timestamp 1644511149
transform 1 0 29808 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_324
timestamp 1644511149
transform 1 0 30912 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_328
timestamp 1644511149
transform 1 0 31280 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_332
timestamp 1644511149
transform 1 0 31648 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_340
timestamp 1644511149
transform 1 0 32384 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_367
timestamp 1644511149
transform 1 0 34868 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_374
timestamp 1644511149
transform 1 0 35512 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_381
timestamp 1644511149
transform 1 0 36156 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_388
timestamp 1644511149
transform 1 0 36800 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_414
timestamp 1644511149
transform 1 0 39192 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_3_425
timestamp 1644511149
transform 1 0 40204 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_437
timestamp 1644511149
transform 1 0 41308 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_444
timestamp 1644511149
transform 1 0 41952 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_470
timestamp 1644511149
transform 1 0 44344 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_495
timestamp 1644511149
transform 1 0 46644 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_503
timestamp 1644511149
transform 1 0 47380 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_508
timestamp 1644511149
transform 1 0 47840 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_4_24
timestamp 1644511149
transform 1 0 3312 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_32
timestamp 1644511149
transform 1 0 4048 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_40
timestamp 1644511149
transform 1 0 4784 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_63
timestamp 1644511149
transform 1 0 6900 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_71
timestamp 1644511149
transform 1 0 7636 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_78
timestamp 1644511149
transform 1 0 8280 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_4_88
timestamp 1644511149
transform 1 0 9200 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_100
timestamp 1644511149
transform 1 0 10304 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_112
timestamp 1644511149
transform 1 0 11408 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_124
timestamp 1644511149
transform 1 0 12512 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_136
timestamp 1644511149
transform 1 0 13616 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_141
timestamp 1644511149
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_153
timestamp 1644511149
transform 1 0 15180 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_4_162
timestamp 1644511149
transform 1 0 16008 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_174
timestamp 1644511149
transform 1 0 17112 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_186
timestamp 1644511149
transform 1 0 18216 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_194
timestamp 1644511149
transform 1 0 18952 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_4_197
timestamp 1644511149
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_209
timestamp 1644511149
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_221
timestamp 1644511149
transform 1 0 21436 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_233
timestamp 1644511149
transform 1 0 22540 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_245
timestamp 1644511149
transform 1 0 23644 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_251
timestamp 1644511149
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_253
timestamp 1644511149
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_265
timestamp 1644511149
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_277
timestamp 1644511149
transform 1 0 26588 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_289
timestamp 1644511149
transform 1 0 27692 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_294
timestamp 1644511149
transform 1 0 28152 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_301
timestamp 1644511149
transform 1 0 28796 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_307
timestamp 1644511149
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_309
timestamp 1644511149
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_321
timestamp 1644511149
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_333
timestamp 1644511149
transform 1 0 31740 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_4_339
timestamp 1644511149
transform 1 0 32292 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_4_350
timestamp 1644511149
transform 1 0 33304 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_356
timestamp 1644511149
transform 1 0 33856 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_360
timestamp 1644511149
transform 1 0 34224 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_368
timestamp 1644511149
transform 1 0 34960 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_376
timestamp 1644511149
transform 1 0 35696 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_381
timestamp 1644511149
transform 1 0 36156 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_389
timestamp 1644511149
transform 1 0 36892 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_393
timestamp 1644511149
transform 1 0 37260 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_405
timestamp 1644511149
transform 1 0 38364 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_417
timestamp 1644511149
transform 1 0 39468 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_421
timestamp 1644511149
transform 1 0 39836 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_433
timestamp 1644511149
transform 1 0 40940 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_445
timestamp 1644511149
transform 1 0 42044 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_451
timestamp 1644511149
transform 1 0 42596 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_455
timestamp 1644511149
transform 1 0 42964 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_459
timestamp 1644511149
transform 1 0 43332 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_466
timestamp 1644511149
transform 1 0 43976 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_474
timestamp 1644511149
transform 1 0 44712 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_477
timestamp 1644511149
transform 1 0 44988 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_482
timestamp 1644511149
transform 1 0 45448 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_490
timestamp 1644511149
transform 1 0 46184 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_512
timestamp 1644511149
transform 1 0 48208 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_3
timestamp 1644511149
transform 1 0 1380 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_7
timestamp 1644511149
transform 1 0 1748 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_5_32
timestamp 1644511149
transform 1 0 4048 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_5_44
timestamp 1644511149
transform 1 0 5152 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_5_50
timestamp 1644511149
transform 1 0 5704 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_5_57
timestamp 1644511149
transform 1 0 6348 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_5_64
timestamp 1644511149
transform 1 0 6992 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_76
timestamp 1644511149
transform 1 0 8096 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_88
timestamp 1644511149
transform 1 0 9200 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_100
timestamp 1644511149
transform 1 0 10304 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_113
timestamp 1644511149
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_125
timestamp 1644511149
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_137
timestamp 1644511149
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_149
timestamp 1644511149
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp 1644511149
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1644511149
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_169
timestamp 1644511149
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_181
timestamp 1644511149
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_193
timestamp 1644511149
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_205
timestamp 1644511149
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_217
timestamp 1644511149
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_223
timestamp 1644511149
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_225
timestamp 1644511149
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_237
timestamp 1644511149
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_249
timestamp 1644511149
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_261
timestamp 1644511149
transform 1 0 25116 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_273
timestamp 1644511149
transform 1 0 26220 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_279
timestamp 1644511149
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_281
timestamp 1644511149
transform 1 0 26956 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_289
timestamp 1644511149
transform 1 0 27692 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_295
timestamp 1644511149
transform 1 0 28244 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_307
timestamp 1644511149
transform 1 0 29348 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_319
timestamp 1644511149
transform 1 0 30452 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_331
timestamp 1644511149
transform 1 0 31556 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_335
timestamp 1644511149
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_337
timestamp 1644511149
transform 1 0 32108 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_345
timestamp 1644511149
transform 1 0 32844 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_350
timestamp 1644511149
transform 1 0 33304 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_362
timestamp 1644511149
transform 1 0 34408 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_374
timestamp 1644511149
transform 1 0 35512 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_386
timestamp 1644511149
transform 1 0 36616 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_5_393
timestamp 1644511149
transform 1 0 37260 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_405
timestamp 1644511149
transform 1 0 38364 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_417
timestamp 1644511149
transform 1 0 39468 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_429
timestamp 1644511149
transform 1 0 40572 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_441
timestamp 1644511149
transform 1 0 41676 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_447
timestamp 1644511149
transform 1 0 42228 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_449
timestamp 1644511149
transform 1 0 42412 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_461
timestamp 1644511149
transform 1 0 43516 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_468
timestamp 1644511149
transform 1 0 44160 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_475
timestamp 1644511149
transform 1 0 44804 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_500
timestamp 1644511149
transform 1 0 47104 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_508
timestamp 1644511149
transform 1 0 47840 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_6_3
timestamp 1644511149
transform 1 0 1380 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_10
timestamp 1644511149
transform 1 0 2024 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_17
timestamp 1644511149
transform 1 0 2668 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_24
timestamp 1644511149
transform 1 0 3312 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_29
timestamp 1644511149
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_41
timestamp 1644511149
transform 1 0 4876 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_49
timestamp 1644511149
transform 1 0 5612 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_53
timestamp 1644511149
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_65
timestamp 1644511149
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 1644511149
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1644511149
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_85
timestamp 1644511149
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_97
timestamp 1644511149
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_109
timestamp 1644511149
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_121
timestamp 1644511149
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1644511149
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1644511149
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_141
timestamp 1644511149
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_153
timestamp 1644511149
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_165
timestamp 1644511149
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_177
timestamp 1644511149
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_189
timestamp 1644511149
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1644511149
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_197
timestamp 1644511149
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_209
timestamp 1644511149
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_221
timestamp 1644511149
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_233
timestamp 1644511149
transform 1 0 22540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_245
timestamp 1644511149
transform 1 0 23644 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp 1644511149
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_253
timestamp 1644511149
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_265
timestamp 1644511149
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_277
timestamp 1644511149
transform 1 0 26588 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_289
timestamp 1644511149
transform 1 0 27692 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_301
timestamp 1644511149
transform 1 0 28796 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_307
timestamp 1644511149
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_309
timestamp 1644511149
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_321
timestamp 1644511149
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_333
timestamp 1644511149
transform 1 0 31740 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_345
timestamp 1644511149
transform 1 0 32844 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_357
timestamp 1644511149
transform 1 0 33948 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_363
timestamp 1644511149
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_365
timestamp 1644511149
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_377
timestamp 1644511149
transform 1 0 35788 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_389
timestamp 1644511149
transform 1 0 36892 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_401
timestamp 1644511149
transform 1 0 37996 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_413
timestamp 1644511149
transform 1 0 39100 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_419
timestamp 1644511149
transform 1 0 39652 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_421
timestamp 1644511149
transform 1 0 39836 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_433
timestamp 1644511149
transform 1 0 40940 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_445
timestamp 1644511149
transform 1 0 42044 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_457
timestamp 1644511149
transform 1 0 43148 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_469
timestamp 1644511149
transform 1 0 44252 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_475
timestamp 1644511149
transform 1 0 44804 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_480
timestamp 1644511149
transform 1 0 45264 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_487
timestamp 1644511149
transform 1 0 45908 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_512
timestamp 1644511149
transform 1 0 48208 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_3
timestamp 1644511149
transform 1 0 1380 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_7_32
timestamp 1644511149
transform 1 0 4048 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_44
timestamp 1644511149
transform 1 0 5152 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_57
timestamp 1644511149
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_69
timestamp 1644511149
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_81
timestamp 1644511149
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_93
timestamp 1644511149
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 1644511149
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1644511149
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_113
timestamp 1644511149
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_125
timestamp 1644511149
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_137
timestamp 1644511149
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_149
timestamp 1644511149
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_161
timestamp 1644511149
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1644511149
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_169
timestamp 1644511149
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_181
timestamp 1644511149
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_193
timestamp 1644511149
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_205
timestamp 1644511149
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_217
timestamp 1644511149
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp 1644511149
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_225
timestamp 1644511149
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_237
timestamp 1644511149
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_249
timestamp 1644511149
transform 1 0 24012 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_261
timestamp 1644511149
transform 1 0 25116 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_273
timestamp 1644511149
transform 1 0 26220 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_279
timestamp 1644511149
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_281
timestamp 1644511149
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_293
timestamp 1644511149
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_305
timestamp 1644511149
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_317
timestamp 1644511149
transform 1 0 30268 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_329
timestamp 1644511149
transform 1 0 31372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_335
timestamp 1644511149
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_337
timestamp 1644511149
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_349
timestamp 1644511149
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_361
timestamp 1644511149
transform 1 0 34316 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_373
timestamp 1644511149
transform 1 0 35420 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_385
timestamp 1644511149
transform 1 0 36524 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_391
timestamp 1644511149
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_393
timestamp 1644511149
transform 1 0 37260 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_405
timestamp 1644511149
transform 1 0 38364 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_417
timestamp 1644511149
transform 1 0 39468 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_429
timestamp 1644511149
transform 1 0 40572 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_441
timestamp 1644511149
transform 1 0 41676 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_447
timestamp 1644511149
transform 1 0 42228 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_449
timestamp 1644511149
transform 1 0 42412 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_461
timestamp 1644511149
transform 1 0 43516 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_473
timestamp 1644511149
transform 1 0 44620 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_7_500
timestamp 1644511149
transform 1 0 47104 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_508
timestamp 1644511149
transform 1 0 47840 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_8_3
timestamp 1644511149
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_18
timestamp 1644511149
transform 1 0 2760 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_26
timestamp 1644511149
transform 1 0 3496 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_8_29
timestamp 1644511149
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_41
timestamp 1644511149
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_53
timestamp 1644511149
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_65
timestamp 1644511149
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1644511149
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1644511149
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_85
timestamp 1644511149
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_97
timestamp 1644511149
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_109
timestamp 1644511149
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_121
timestamp 1644511149
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_133
timestamp 1644511149
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1644511149
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_141
timestamp 1644511149
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_153
timestamp 1644511149
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_165
timestamp 1644511149
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_177
timestamp 1644511149
transform 1 0 17388 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_8_188
timestamp 1644511149
transform 1 0 18400 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_8_197
timestamp 1644511149
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_209
timestamp 1644511149
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_221
timestamp 1644511149
transform 1 0 21436 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_233
timestamp 1644511149
transform 1 0 22540 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_245
timestamp 1644511149
transform 1 0 23644 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_251
timestamp 1644511149
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_253
timestamp 1644511149
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_265
timestamp 1644511149
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_277
timestamp 1644511149
transform 1 0 26588 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_289
timestamp 1644511149
transform 1 0 27692 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_301
timestamp 1644511149
transform 1 0 28796 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_307
timestamp 1644511149
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_309
timestamp 1644511149
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_321
timestamp 1644511149
transform 1 0 30636 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_333
timestamp 1644511149
transform 1 0 31740 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_345
timestamp 1644511149
transform 1 0 32844 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_353
timestamp 1644511149
transform 1 0 33580 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_357
timestamp 1644511149
transform 1 0 33948 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_363
timestamp 1644511149
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_365
timestamp 1644511149
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_377
timestamp 1644511149
transform 1 0 35788 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_389
timestamp 1644511149
transform 1 0 36892 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_401
timestamp 1644511149
transform 1 0 37996 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_413
timestamp 1644511149
transform 1 0 39100 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_419
timestamp 1644511149
transform 1 0 39652 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_421
timestamp 1644511149
transform 1 0 39836 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_433
timestamp 1644511149
transform 1 0 40940 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_445
timestamp 1644511149
transform 1 0 42044 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_457
timestamp 1644511149
transform 1 0 43148 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_469
timestamp 1644511149
transform 1 0 44252 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_475
timestamp 1644511149
transform 1 0 44804 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_477
timestamp 1644511149
transform 1 0 44988 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_489
timestamp 1644511149
transform 1 0 46092 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_495
timestamp 1644511149
transform 1 0 46644 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_499
timestamp 1644511149
transform 1 0 47012 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_503
timestamp 1644511149
transform 1 0 47380 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_507
timestamp 1644511149
transform 1 0 47748 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_515
timestamp 1644511149
transform 1 0 48484 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_3
timestamp 1644511149
transform 1 0 1380 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_11
timestamp 1644511149
transform 1 0 2116 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_15
timestamp 1644511149
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_27
timestamp 1644511149
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_39
timestamp 1644511149
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_51
timestamp 1644511149
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1644511149
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_57
timestamp 1644511149
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_69
timestamp 1644511149
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_81
timestamp 1644511149
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_93
timestamp 1644511149
transform 1 0 9660 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_9_104
timestamp 1644511149
transform 1 0 10672 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_9_113
timestamp 1644511149
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_125
timestamp 1644511149
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_137
timestamp 1644511149
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_149
timestamp 1644511149
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_161
timestamp 1644511149
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1644511149
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_169
timestamp 1644511149
transform 1 0 16652 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_177
timestamp 1644511149
transform 1 0 17388 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_201
timestamp 1644511149
transform 1 0 19596 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_213
timestamp 1644511149
transform 1 0 20700 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_221
timestamp 1644511149
transform 1 0 21436 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_225
timestamp 1644511149
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_237
timestamp 1644511149
transform 1 0 22908 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_249
timestamp 1644511149
transform 1 0 24012 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_261
timestamp 1644511149
transform 1 0 25116 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_273
timestamp 1644511149
transform 1 0 26220 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_279
timestamp 1644511149
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_281
timestamp 1644511149
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_293
timestamp 1644511149
transform 1 0 28060 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_301
timestamp 1644511149
transform 1 0 28796 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_307
timestamp 1644511149
transform 1 0 29348 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_332
timestamp 1644511149
transform 1 0 31648 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_9_337
timestamp 1644511149
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_349
timestamp 1644511149
transform 1 0 33212 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_353
timestamp 1644511149
transform 1 0 33580 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_375
timestamp 1644511149
transform 1 0 35604 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_387
timestamp 1644511149
transform 1 0 36708 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_391
timestamp 1644511149
transform 1 0 37076 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_393
timestamp 1644511149
transform 1 0 37260 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_405
timestamp 1644511149
transform 1 0 38364 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_417
timestamp 1644511149
transform 1 0 39468 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_429
timestamp 1644511149
transform 1 0 40572 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_441
timestamp 1644511149
transform 1 0 41676 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_447
timestamp 1644511149
transform 1 0 42228 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_449
timestamp 1644511149
transform 1 0 42412 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_461
timestamp 1644511149
transform 1 0 43516 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_473
timestamp 1644511149
transform 1 0 44620 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_485
timestamp 1644511149
transform 1 0 45724 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_497
timestamp 1644511149
transform 1 0 46828 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_503
timestamp 1644511149
transform 1 0 47380 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_505
timestamp 1644511149
transform 1 0 47564 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_513
timestamp 1644511149
transform 1 0 48300 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_10_3
timestamp 1644511149
transform 1 0 1380 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_11
timestamp 1644511149
transform 1 0 2116 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_15
timestamp 1644511149
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1644511149
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_29
timestamp 1644511149
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_41
timestamp 1644511149
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_53
timestamp 1644511149
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_65
timestamp 1644511149
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp 1644511149
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1644511149
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_85
timestamp 1644511149
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_10_97
timestamp 1644511149
transform 1 0 10028 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_121
timestamp 1644511149
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_133
timestamp 1644511149
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1644511149
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_141
timestamp 1644511149
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_153
timestamp 1644511149
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_165
timestamp 1644511149
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_10_177
timestamp 1644511149
transform 1 0 17388 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_183
timestamp 1644511149
transform 1 0 17940 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_195
timestamp 1644511149
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_197
timestamp 1644511149
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_209
timestamp 1644511149
transform 1 0 20332 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_221
timestamp 1644511149
transform 1 0 21436 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_233
timestamp 1644511149
transform 1 0 22540 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_245
timestamp 1644511149
transform 1 0 23644 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_251
timestamp 1644511149
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_253
timestamp 1644511149
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_265
timestamp 1644511149
transform 1 0 25484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_277
timestamp 1644511149
transform 1 0 26588 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_289
timestamp 1644511149
transform 1 0 27692 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_301
timestamp 1644511149
transform 1 0 28796 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_307
timestamp 1644511149
transform 1 0 29348 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_309
timestamp 1644511149
transform 1 0 29532 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_315
timestamp 1644511149
transform 1 0 30084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_327
timestamp 1644511149
transform 1 0 31188 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_339
timestamp 1644511149
transform 1 0 32292 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_347
timestamp 1644511149
transform 1 0 33028 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_10_352
timestamp 1644511149
transform 1 0 33488 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_365
timestamp 1644511149
transform 1 0 34684 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_377
timestamp 1644511149
transform 1 0 35788 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_389
timestamp 1644511149
transform 1 0 36892 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_401
timestamp 1644511149
transform 1 0 37996 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_413
timestamp 1644511149
transform 1 0 39100 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_419
timestamp 1644511149
transform 1 0 39652 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_421
timestamp 1644511149
transform 1 0 39836 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_433
timestamp 1644511149
transform 1 0 40940 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_445
timestamp 1644511149
transform 1 0 42044 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_457
timestamp 1644511149
transform 1 0 43148 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_469
timestamp 1644511149
transform 1 0 44252 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_475
timestamp 1644511149
transform 1 0 44804 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_477
timestamp 1644511149
transform 1 0 44988 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_489
timestamp 1644511149
transform 1 0 46092 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_501
timestamp 1644511149
transform 1 0 47196 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_10_513
timestamp 1644511149
transform 1 0 48300 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_11_3
timestamp 1644511149
transform 1 0 1380 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_9
timestamp 1644511149
transform 1 0 1932 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_31
timestamp 1644511149
transform 1 0 3956 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_43
timestamp 1644511149
transform 1 0 5060 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1644511149
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_57
timestamp 1644511149
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_69
timestamp 1644511149
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_81
timestamp 1644511149
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_93
timestamp 1644511149
transform 1 0 9660 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_11_104
timestamp 1644511149
transform 1 0 10672 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_11_113
timestamp 1644511149
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_125
timestamp 1644511149
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_137
timestamp 1644511149
transform 1 0 13708 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_149
timestamp 1644511149
transform 1 0 14812 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_161
timestamp 1644511149
transform 1 0 15916 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp 1644511149
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_169
timestamp 1644511149
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_181
timestamp 1644511149
transform 1 0 17756 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_193
timestamp 1644511149
transform 1 0 18860 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_205
timestamp 1644511149
transform 1 0 19964 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_217
timestamp 1644511149
transform 1 0 21068 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_223
timestamp 1644511149
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_225
timestamp 1644511149
transform 1 0 21804 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_237
timestamp 1644511149
transform 1 0 22908 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_249
timestamp 1644511149
transform 1 0 24012 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_261
timestamp 1644511149
transform 1 0 25116 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_273
timestamp 1644511149
transform 1 0 26220 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_279
timestamp 1644511149
transform 1 0 26772 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_281
timestamp 1644511149
transform 1 0 26956 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_293
timestamp 1644511149
transform 1 0 28060 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_305
timestamp 1644511149
transform 1 0 29164 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_317
timestamp 1644511149
transform 1 0 30268 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_329
timestamp 1644511149
transform 1 0 31372 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_335
timestamp 1644511149
transform 1 0 31924 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_337
timestamp 1644511149
transform 1 0 32108 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_349
timestamp 1644511149
transform 1 0 33212 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_361
timestamp 1644511149
transform 1 0 34316 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_373
timestamp 1644511149
transform 1 0 35420 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_385
timestamp 1644511149
transform 1 0 36524 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_391
timestamp 1644511149
transform 1 0 37076 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_393
timestamp 1644511149
transform 1 0 37260 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_405
timestamp 1644511149
transform 1 0 38364 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_417
timestamp 1644511149
transform 1 0 39468 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_429
timestamp 1644511149
transform 1 0 40572 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_441
timestamp 1644511149
transform 1 0 41676 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_447
timestamp 1644511149
transform 1 0 42228 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_449
timestamp 1644511149
transform 1 0 42412 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_461
timestamp 1644511149
transform 1 0 43516 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_473
timestamp 1644511149
transform 1 0 44620 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_485
timestamp 1644511149
transform 1 0 45724 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_497
timestamp 1644511149
transform 1 0 46828 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_503
timestamp 1644511149
transform 1 0 47380 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_505
timestamp 1644511149
transform 1 0 47564 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_513
timestamp 1644511149
transform 1 0 48300 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_12_3
timestamp 1644511149
transform 1 0 1380 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_9
timestamp 1644511149
transform 1 0 1932 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_13
timestamp 1644511149
transform 1 0 2300 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_12_25
timestamp 1644511149
transform 1 0 3404 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_29
timestamp 1644511149
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_41
timestamp 1644511149
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_53
timestamp 1644511149
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_65
timestamp 1644511149
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 1644511149
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1644511149
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_85
timestamp 1644511149
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_97
timestamp 1644511149
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_109
timestamp 1644511149
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_121
timestamp 1644511149
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_133
timestamp 1644511149
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1644511149
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_141
timestamp 1644511149
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_153
timestamp 1644511149
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_165
timestamp 1644511149
transform 1 0 16284 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_177
timestamp 1644511149
transform 1 0 17388 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_189
timestamp 1644511149
transform 1 0 18492 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_195
timestamp 1644511149
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_197
timestamp 1644511149
transform 1 0 19228 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_209
timestamp 1644511149
transform 1 0 20332 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_221
timestamp 1644511149
transform 1 0 21436 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_233
timestamp 1644511149
transform 1 0 22540 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_245
timestamp 1644511149
transform 1 0 23644 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_251
timestamp 1644511149
transform 1 0 24196 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_253
timestamp 1644511149
transform 1 0 24380 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_265
timestamp 1644511149
transform 1 0 25484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_277
timestamp 1644511149
transform 1 0 26588 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_289
timestamp 1644511149
transform 1 0 27692 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_301
timestamp 1644511149
transform 1 0 28796 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_307
timestamp 1644511149
transform 1 0 29348 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_309
timestamp 1644511149
transform 1 0 29532 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_321
timestamp 1644511149
transform 1 0 30636 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_333
timestamp 1644511149
transform 1 0 31740 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_345
timestamp 1644511149
transform 1 0 32844 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_357
timestamp 1644511149
transform 1 0 33948 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_363
timestamp 1644511149
transform 1 0 34500 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_365
timestamp 1644511149
transform 1 0 34684 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_377
timestamp 1644511149
transform 1 0 35788 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_389
timestamp 1644511149
transform 1 0 36892 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_401
timestamp 1644511149
transform 1 0 37996 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_413
timestamp 1644511149
transform 1 0 39100 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_419
timestamp 1644511149
transform 1 0 39652 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_421
timestamp 1644511149
transform 1 0 39836 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_12_426
timestamp 1644511149
transform 1 0 40296 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_438
timestamp 1644511149
transform 1 0 41400 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_450
timestamp 1644511149
transform 1 0 42504 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_462
timestamp 1644511149
transform 1 0 43608 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_474
timestamp 1644511149
transform 1 0 44712 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_12_477
timestamp 1644511149
transform 1 0 44988 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_489
timestamp 1644511149
transform 1 0 46092 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_501
timestamp 1644511149
transform 1 0 47196 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_12_513
timestamp 1644511149
transform 1 0 48300 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_13_3
timestamp 1644511149
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_15
timestamp 1644511149
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_27
timestamp 1644511149
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_39
timestamp 1644511149
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_51
timestamp 1644511149
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1644511149
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_57
timestamp 1644511149
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_69
timestamp 1644511149
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_81
timestamp 1644511149
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_93
timestamp 1644511149
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_105
timestamp 1644511149
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1644511149
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_116
timestamp 1644511149
transform 1 0 11776 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_13_128
timestamp 1644511149
transform 1 0 12880 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_150
timestamp 1644511149
transform 1 0 14904 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_162
timestamp 1644511149
transform 1 0 16008 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_13_169
timestamp 1644511149
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_181
timestamp 1644511149
transform 1 0 17756 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_193
timestamp 1644511149
transform 1 0 18860 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_205
timestamp 1644511149
transform 1 0 19964 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_217
timestamp 1644511149
transform 1 0 21068 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_223
timestamp 1644511149
transform 1 0 21620 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_225
timestamp 1644511149
transform 1 0 21804 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_237
timestamp 1644511149
transform 1 0 22908 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_249
timestamp 1644511149
transform 1 0 24012 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_261
timestamp 1644511149
transform 1 0 25116 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_273
timestamp 1644511149
transform 1 0 26220 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_279
timestamp 1644511149
transform 1 0 26772 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_281
timestamp 1644511149
transform 1 0 26956 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_293
timestamp 1644511149
transform 1 0 28060 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_305
timestamp 1644511149
transform 1 0 29164 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_317
timestamp 1644511149
transform 1 0 30268 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_329
timestamp 1644511149
transform 1 0 31372 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_335
timestamp 1644511149
transform 1 0 31924 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_337
timestamp 1644511149
transform 1 0 32108 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_349
timestamp 1644511149
transform 1 0 33212 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_361
timestamp 1644511149
transform 1 0 34316 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_373
timestamp 1644511149
transform 1 0 35420 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_385
timestamp 1644511149
transform 1 0 36524 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_391
timestamp 1644511149
transform 1 0 37076 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_393
timestamp 1644511149
transform 1 0 37260 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_405
timestamp 1644511149
transform 1 0 38364 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_417
timestamp 1644511149
transform 1 0 39468 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_13_444
timestamp 1644511149
transform 1 0 41952 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_13_449
timestamp 1644511149
transform 1 0 42412 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_461
timestamp 1644511149
transform 1 0 43516 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_473
timestamp 1644511149
transform 1 0 44620 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_485
timestamp 1644511149
transform 1 0 45724 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_497
timestamp 1644511149
transform 1 0 46828 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_503
timestamp 1644511149
transform 1 0 47380 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_508
timestamp 1644511149
transform 1 0 47840 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_14_3
timestamp 1644511149
transform 1 0 1380 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_11
timestamp 1644511149
transform 1 0 2116 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_14_17
timestamp 1644511149
transform 1 0 2668 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_25
timestamp 1644511149
transform 1 0 3404 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_14_29
timestamp 1644511149
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_41
timestamp 1644511149
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_53
timestamp 1644511149
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_65
timestamp 1644511149
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp 1644511149
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1644511149
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_85
timestamp 1644511149
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_97
timestamp 1644511149
transform 1 0 10028 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_105
timestamp 1644511149
transform 1 0 10764 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_129
timestamp 1644511149
transform 1 0 12972 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_136
timestamp 1644511149
transform 1 0 13616 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_14_141
timestamp 1644511149
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_153
timestamp 1644511149
transform 1 0 15180 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_165
timestamp 1644511149
transform 1 0 16284 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_177
timestamp 1644511149
transform 1 0 17388 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_189
timestamp 1644511149
transform 1 0 18492 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_195
timestamp 1644511149
transform 1 0 19044 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_197
timestamp 1644511149
transform 1 0 19228 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_209
timestamp 1644511149
transform 1 0 20332 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_221
timestamp 1644511149
transform 1 0 21436 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_233
timestamp 1644511149
transform 1 0 22540 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_245
timestamp 1644511149
transform 1 0 23644 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_251
timestamp 1644511149
transform 1 0 24196 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_253
timestamp 1644511149
transform 1 0 24380 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_265
timestamp 1644511149
transform 1 0 25484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_277
timestamp 1644511149
transform 1 0 26588 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_289
timestamp 1644511149
transform 1 0 27692 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_301
timestamp 1644511149
transform 1 0 28796 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_307
timestamp 1644511149
transform 1 0 29348 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_309
timestamp 1644511149
transform 1 0 29532 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_321
timestamp 1644511149
transform 1 0 30636 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_333
timestamp 1644511149
transform 1 0 31740 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_345
timestamp 1644511149
transform 1 0 32844 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_357
timestamp 1644511149
transform 1 0 33948 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_363
timestamp 1644511149
transform 1 0 34500 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_365
timestamp 1644511149
transform 1 0 34684 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_377
timestamp 1644511149
transform 1 0 35788 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_389
timestamp 1644511149
transform 1 0 36892 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_401
timestamp 1644511149
transform 1 0 37996 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_413
timestamp 1644511149
transform 1 0 39100 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_419
timestamp 1644511149
transform 1 0 39652 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_421
timestamp 1644511149
transform 1 0 39836 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_14_426
timestamp 1644511149
transform 1 0 40296 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_438
timestamp 1644511149
transform 1 0 41400 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_450
timestamp 1644511149
transform 1 0 42504 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_462
timestamp 1644511149
transform 1 0 43608 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_474
timestamp 1644511149
transform 1 0 44712 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_14_477
timestamp 1644511149
transform 1 0 44988 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_489
timestamp 1644511149
transform 1 0 46092 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_512
timestamp 1644511149
transform 1 0 48208 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_3
timestamp 1644511149
transform 1 0 1380 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_9
timestamp 1644511149
transform 1 0 1932 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_31
timestamp 1644511149
transform 1 0 3956 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_43
timestamp 1644511149
transform 1 0 5060 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1644511149
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_57
timestamp 1644511149
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_69
timestamp 1644511149
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_81
timestamp 1644511149
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_93
timestamp 1644511149
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_105
timestamp 1644511149
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1644511149
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_116
timestamp 1644511149
transform 1 0 11776 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_128
timestamp 1644511149
transform 1 0 12880 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_132
timestamp 1644511149
transform 1 0 13248 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_144
timestamp 1644511149
transform 1 0 14352 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_156
timestamp 1644511149
transform 1 0 15456 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_169
timestamp 1644511149
transform 1 0 16652 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_181
timestamp 1644511149
transform 1 0 17756 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_193
timestamp 1644511149
transform 1 0 18860 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_205
timestamp 1644511149
transform 1 0 19964 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_217
timestamp 1644511149
transform 1 0 21068 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_223
timestamp 1644511149
transform 1 0 21620 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_225
timestamp 1644511149
transform 1 0 21804 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_237
timestamp 1644511149
transform 1 0 22908 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_249
timestamp 1644511149
transform 1 0 24012 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_261
timestamp 1644511149
transform 1 0 25116 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_273
timestamp 1644511149
transform 1 0 26220 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_279
timestamp 1644511149
transform 1 0 26772 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_281
timestamp 1644511149
transform 1 0 26956 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_293
timestamp 1644511149
transform 1 0 28060 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_305
timestamp 1644511149
transform 1 0 29164 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_317
timestamp 1644511149
transform 1 0 30268 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_329
timestamp 1644511149
transform 1 0 31372 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_335
timestamp 1644511149
transform 1 0 31924 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_337
timestamp 1644511149
transform 1 0 32108 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_349
timestamp 1644511149
transform 1 0 33212 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_361
timestamp 1644511149
transform 1 0 34316 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_373
timestamp 1644511149
transform 1 0 35420 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_385
timestamp 1644511149
transform 1 0 36524 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_391
timestamp 1644511149
transform 1 0 37076 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_393
timestamp 1644511149
transform 1 0 37260 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_405
timestamp 1644511149
transform 1 0 38364 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_417
timestamp 1644511149
transform 1 0 39468 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_429
timestamp 1644511149
transform 1 0 40572 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_441
timestamp 1644511149
transform 1 0 41676 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_447
timestamp 1644511149
transform 1 0 42228 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_449
timestamp 1644511149
transform 1 0 42412 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_461
timestamp 1644511149
transform 1 0 43516 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_473
timestamp 1644511149
transform 1 0 44620 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_485
timestamp 1644511149
transform 1 0 45724 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_489
timestamp 1644511149
transform 1 0 46092 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_496
timestamp 1644511149
transform 1 0 46736 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_15_508
timestamp 1644511149
transform 1 0 47840 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_16_3
timestamp 1644511149
transform 1 0 1380 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_16_14
timestamp 1644511149
transform 1 0 2392 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_26
timestamp 1644511149
transform 1 0 3496 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_16_29
timestamp 1644511149
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_41
timestamp 1644511149
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_53
timestamp 1644511149
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_65
timestamp 1644511149
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp 1644511149
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1644511149
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_85
timestamp 1644511149
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_97
timestamp 1644511149
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_109
timestamp 1644511149
transform 1 0 11132 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_121
timestamp 1644511149
transform 1 0 12236 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_133
timestamp 1644511149
transform 1 0 13340 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 1644511149
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_141
timestamp 1644511149
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_153
timestamp 1644511149
transform 1 0 15180 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_165
timestamp 1644511149
transform 1 0 16284 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_177
timestamp 1644511149
transform 1 0 17388 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_189
timestamp 1644511149
transform 1 0 18492 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_195
timestamp 1644511149
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_197
timestamp 1644511149
transform 1 0 19228 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_209
timestamp 1644511149
transform 1 0 20332 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_221
timestamp 1644511149
transform 1 0 21436 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_233
timestamp 1644511149
transform 1 0 22540 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_245
timestamp 1644511149
transform 1 0 23644 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_251
timestamp 1644511149
transform 1 0 24196 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_253
timestamp 1644511149
transform 1 0 24380 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_265
timestamp 1644511149
transform 1 0 25484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_277
timestamp 1644511149
transform 1 0 26588 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_289
timestamp 1644511149
transform 1 0 27692 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_301
timestamp 1644511149
transform 1 0 28796 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_307
timestamp 1644511149
transform 1 0 29348 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_309
timestamp 1644511149
transform 1 0 29532 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_321
timestamp 1644511149
transform 1 0 30636 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_333
timestamp 1644511149
transform 1 0 31740 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_345
timestamp 1644511149
transform 1 0 32844 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_357
timestamp 1644511149
transform 1 0 33948 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_363
timestamp 1644511149
transform 1 0 34500 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_365
timestamp 1644511149
transform 1 0 34684 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_377
timestamp 1644511149
transform 1 0 35788 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_389
timestamp 1644511149
transform 1 0 36892 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_401
timestamp 1644511149
transform 1 0 37996 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_413
timestamp 1644511149
transform 1 0 39100 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_419
timestamp 1644511149
transform 1 0 39652 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_421
timestamp 1644511149
transform 1 0 39836 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_433
timestamp 1644511149
transform 1 0 40940 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_445
timestamp 1644511149
transform 1 0 42044 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_457
timestamp 1644511149
transform 1 0 43148 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_469
timestamp 1644511149
transform 1 0 44252 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_475
timestamp 1644511149
transform 1 0 44804 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_477
timestamp 1644511149
transform 1 0 44988 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_483
timestamp 1644511149
transform 1 0 45540 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_487
timestamp 1644511149
transform 1 0 45908 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_512
timestamp 1644511149
transform 1 0 48208 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_17_3
timestamp 1644511149
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_15
timestamp 1644511149
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_27
timestamp 1644511149
transform 1 0 3588 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_32
timestamp 1644511149
transform 1 0 4048 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_44
timestamp 1644511149
transform 1 0 5152 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_57
timestamp 1644511149
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_69
timestamp 1644511149
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_81
timestamp 1644511149
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_93
timestamp 1644511149
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_105
timestamp 1644511149
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1644511149
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_113
timestamp 1644511149
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_125
timestamp 1644511149
transform 1 0 12604 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_137
timestamp 1644511149
transform 1 0 13708 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_149
timestamp 1644511149
transform 1 0 14812 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_161
timestamp 1644511149
transform 1 0 15916 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_167
timestamp 1644511149
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_169
timestamp 1644511149
transform 1 0 16652 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_181
timestamp 1644511149
transform 1 0 17756 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_193
timestamp 1644511149
transform 1 0 18860 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_205
timestamp 1644511149
transform 1 0 19964 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_217
timestamp 1644511149
transform 1 0 21068 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_223
timestamp 1644511149
transform 1 0 21620 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_225
timestamp 1644511149
transform 1 0 21804 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_237
timestamp 1644511149
transform 1 0 22908 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_249
timestamp 1644511149
transform 1 0 24012 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_261
timestamp 1644511149
transform 1 0 25116 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_273
timestamp 1644511149
transform 1 0 26220 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_279
timestamp 1644511149
transform 1 0 26772 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_281
timestamp 1644511149
transform 1 0 26956 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_293
timestamp 1644511149
transform 1 0 28060 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_305
timestamp 1644511149
transform 1 0 29164 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_317
timestamp 1644511149
transform 1 0 30268 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_329
timestamp 1644511149
transform 1 0 31372 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_335
timestamp 1644511149
transform 1 0 31924 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_337
timestamp 1644511149
transform 1 0 32108 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_349
timestamp 1644511149
transform 1 0 33212 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_361
timestamp 1644511149
transform 1 0 34316 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_373
timestamp 1644511149
transform 1 0 35420 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_385
timestamp 1644511149
transform 1 0 36524 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_391
timestamp 1644511149
transform 1 0 37076 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_393
timestamp 1644511149
transform 1 0 37260 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_405
timestamp 1644511149
transform 1 0 38364 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_417
timestamp 1644511149
transform 1 0 39468 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_429
timestamp 1644511149
transform 1 0 40572 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_441
timestamp 1644511149
transform 1 0 41676 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_447
timestamp 1644511149
transform 1 0 42228 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_449
timestamp 1644511149
transform 1 0 42412 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_461
timestamp 1644511149
transform 1 0 43516 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_469
timestamp 1644511149
transform 1 0 44252 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_475
timestamp 1644511149
transform 1 0 44804 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_500
timestamp 1644511149
transform 1 0 47104 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_508
timestamp 1644511149
transform 1 0 47840 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_18_3
timestamp 1644511149
transform 1 0 1380 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_11
timestamp 1644511149
transform 1 0 2116 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_18_17
timestamp 1644511149
transform 1 0 2668 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_25
timestamp 1644511149
transform 1 0 3404 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_50
timestamp 1644511149
transform 1 0 5704 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_62
timestamp 1644511149
transform 1 0 6808 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_74
timestamp 1644511149
transform 1 0 7912 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_82
timestamp 1644511149
transform 1 0 8648 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_18_85
timestamp 1644511149
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_97
timestamp 1644511149
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_109
timestamp 1644511149
transform 1 0 11132 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_121
timestamp 1644511149
transform 1 0 12236 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_133
timestamp 1644511149
transform 1 0 13340 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_139
timestamp 1644511149
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_141
timestamp 1644511149
transform 1 0 14076 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_153
timestamp 1644511149
transform 1 0 15180 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_165
timestamp 1644511149
transform 1 0 16284 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_177
timestamp 1644511149
transform 1 0 17388 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_189
timestamp 1644511149
transform 1 0 18492 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_195
timestamp 1644511149
transform 1 0 19044 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_197
timestamp 1644511149
transform 1 0 19228 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_209
timestamp 1644511149
transform 1 0 20332 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_221
timestamp 1644511149
transform 1 0 21436 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_233
timestamp 1644511149
transform 1 0 22540 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_245
timestamp 1644511149
transform 1 0 23644 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_251
timestamp 1644511149
transform 1 0 24196 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_253
timestamp 1644511149
transform 1 0 24380 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_265
timestamp 1644511149
transform 1 0 25484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_277
timestamp 1644511149
transform 1 0 26588 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_289
timestamp 1644511149
transform 1 0 27692 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_301
timestamp 1644511149
transform 1 0 28796 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_307
timestamp 1644511149
transform 1 0 29348 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_309
timestamp 1644511149
transform 1 0 29532 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_321
timestamp 1644511149
transform 1 0 30636 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_333
timestamp 1644511149
transform 1 0 31740 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_345
timestamp 1644511149
transform 1 0 32844 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_357
timestamp 1644511149
transform 1 0 33948 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_363
timestamp 1644511149
transform 1 0 34500 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_365
timestamp 1644511149
transform 1 0 34684 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_377
timestamp 1644511149
transform 1 0 35788 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_389
timestamp 1644511149
transform 1 0 36892 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_401
timestamp 1644511149
transform 1 0 37996 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_413
timestamp 1644511149
transform 1 0 39100 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_419
timestamp 1644511149
transform 1 0 39652 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_421
timestamp 1644511149
transform 1 0 39836 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_433
timestamp 1644511149
transform 1 0 40940 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_445
timestamp 1644511149
transform 1 0 42044 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_457
timestamp 1644511149
transform 1 0 43148 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_472
timestamp 1644511149
transform 1 0 44528 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_18_477
timestamp 1644511149
transform 1 0 44988 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_483
timestamp 1644511149
transform 1 0 45540 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_508
timestamp 1644511149
transform 1 0 47840 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_19_3
timestamp 1644511149
transform 1 0 1380 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_9
timestamp 1644511149
transform 1 0 1932 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_31
timestamp 1644511149
transform 1 0 3956 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_43
timestamp 1644511149
transform 1 0 5060 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1644511149
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_57
timestamp 1644511149
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_69
timestamp 1644511149
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_81
timestamp 1644511149
transform 1 0 8556 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_93
timestamp 1644511149
transform 1 0 9660 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_105
timestamp 1644511149
transform 1 0 10764 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1644511149
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_113
timestamp 1644511149
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_125
timestamp 1644511149
transform 1 0 12604 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_137
timestamp 1644511149
transform 1 0 13708 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_149
timestamp 1644511149
transform 1 0 14812 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_161
timestamp 1644511149
transform 1 0 15916 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_167
timestamp 1644511149
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_169
timestamp 1644511149
transform 1 0 16652 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_181
timestamp 1644511149
transform 1 0 17756 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_193
timestamp 1644511149
transform 1 0 18860 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_205
timestamp 1644511149
transform 1 0 19964 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_217
timestamp 1644511149
transform 1 0 21068 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_223
timestamp 1644511149
transform 1 0 21620 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_225
timestamp 1644511149
transform 1 0 21804 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_237
timestamp 1644511149
transform 1 0 22908 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_249
timestamp 1644511149
transform 1 0 24012 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_261
timestamp 1644511149
transform 1 0 25116 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_273
timestamp 1644511149
transform 1 0 26220 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_279
timestamp 1644511149
transform 1 0 26772 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_290
timestamp 1644511149
transform 1 0 27784 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_302
timestamp 1644511149
transform 1 0 28888 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_314
timestamp 1644511149
transform 1 0 29992 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_326
timestamp 1644511149
transform 1 0 31096 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_334
timestamp 1644511149
transform 1 0 31832 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_19_337
timestamp 1644511149
transform 1 0 32108 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_349
timestamp 1644511149
transform 1 0 33212 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_361
timestamp 1644511149
transform 1 0 34316 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_373
timestamp 1644511149
transform 1 0 35420 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_385
timestamp 1644511149
transform 1 0 36524 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_391
timestamp 1644511149
transform 1 0 37076 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_393
timestamp 1644511149
transform 1 0 37260 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_405
timestamp 1644511149
transform 1 0 38364 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_417
timestamp 1644511149
transform 1 0 39468 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_429
timestamp 1644511149
transform 1 0 40572 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_441
timestamp 1644511149
transform 1 0 41676 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_447
timestamp 1644511149
transform 1 0 42228 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_449
timestamp 1644511149
transform 1 0 42412 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_461
timestamp 1644511149
transform 1 0 43516 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_473
timestamp 1644511149
transform 1 0 44620 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_19_500
timestamp 1644511149
transform 1 0 47104 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_508
timestamp 1644511149
transform 1 0 47840 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_20_3
timestamp 1644511149
transform 1 0 1380 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_20_14
timestamp 1644511149
transform 1 0 2392 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_26
timestamp 1644511149
transform 1 0 3496 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_20_32
timestamp 1644511149
transform 1 0 4048 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_44
timestamp 1644511149
transform 1 0 5152 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_56
timestamp 1644511149
transform 1 0 6256 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_68
timestamp 1644511149
transform 1 0 7360 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_80
timestamp 1644511149
transform 1 0 8464 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_20_85
timestamp 1644511149
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_97
timestamp 1644511149
transform 1 0 10028 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_109
timestamp 1644511149
transform 1 0 11132 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_121
timestamp 1644511149
transform 1 0 12236 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_133
timestamp 1644511149
transform 1 0 13340 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_139
timestamp 1644511149
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_141
timestamp 1644511149
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_153
timestamp 1644511149
transform 1 0 15180 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_165
timestamp 1644511149
transform 1 0 16284 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_177
timestamp 1644511149
transform 1 0 17388 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_189
timestamp 1644511149
transform 1 0 18492 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_195
timestamp 1644511149
transform 1 0 19044 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_197
timestamp 1644511149
transform 1 0 19228 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_209
timestamp 1644511149
transform 1 0 20332 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_221
timestamp 1644511149
transform 1 0 21436 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_233
timestamp 1644511149
transform 1 0 22540 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_245
timestamp 1644511149
transform 1 0 23644 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_251
timestamp 1644511149
transform 1 0 24196 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_253
timestamp 1644511149
transform 1 0 24380 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_265
timestamp 1644511149
transform 1 0 25484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_277
timestamp 1644511149
transform 1 0 26588 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_20_288
timestamp 1644511149
transform 1 0 27600 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_300
timestamp 1644511149
transform 1 0 28704 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_20_309
timestamp 1644511149
transform 1 0 29532 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_321
timestamp 1644511149
transform 1 0 30636 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_333
timestamp 1644511149
transform 1 0 31740 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_345
timestamp 1644511149
transform 1 0 32844 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_357
timestamp 1644511149
transform 1 0 33948 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_363
timestamp 1644511149
transform 1 0 34500 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_365
timestamp 1644511149
transform 1 0 34684 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_377
timestamp 1644511149
transform 1 0 35788 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_389
timestamp 1644511149
transform 1 0 36892 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_401
timestamp 1644511149
transform 1 0 37996 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_413
timestamp 1644511149
transform 1 0 39100 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_419
timestamp 1644511149
transform 1 0 39652 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_421
timestamp 1644511149
transform 1 0 39836 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_433
timestamp 1644511149
transform 1 0 40940 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_445
timestamp 1644511149
transform 1 0 42044 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_457
timestamp 1644511149
transform 1 0 43148 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_469
timestamp 1644511149
transform 1 0 44252 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_475
timestamp 1644511149
transform 1 0 44804 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_480
timestamp 1644511149
transform 1 0 45264 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_487
timestamp 1644511149
transform 1 0 45908 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_512
timestamp 1644511149
transform 1 0 48208 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_3
timestamp 1644511149
transform 1 0 1380 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_9
timestamp 1644511149
transform 1 0 1932 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_31
timestamp 1644511149
transform 1 0 3956 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_43
timestamp 1644511149
transform 1 0 5060 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1644511149
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_57
timestamp 1644511149
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_69
timestamp 1644511149
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_81
timestamp 1644511149
transform 1 0 8556 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_93
timestamp 1644511149
transform 1 0 9660 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_105
timestamp 1644511149
transform 1 0 10764 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 1644511149
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_113
timestamp 1644511149
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_125
timestamp 1644511149
transform 1 0 12604 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_137
timestamp 1644511149
transform 1 0 13708 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_149
timestamp 1644511149
transform 1 0 14812 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_161
timestamp 1644511149
transform 1 0 15916 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_167
timestamp 1644511149
transform 1 0 16468 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_169
timestamp 1644511149
transform 1 0 16652 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_181
timestamp 1644511149
transform 1 0 17756 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_193
timestamp 1644511149
transform 1 0 18860 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_205
timestamp 1644511149
transform 1 0 19964 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_217
timestamp 1644511149
transform 1 0 21068 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_223
timestamp 1644511149
transform 1 0 21620 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_225
timestamp 1644511149
transform 1 0 21804 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_237
timestamp 1644511149
transform 1 0 22908 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_249
timestamp 1644511149
transform 1 0 24012 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_270
timestamp 1644511149
transform 1 0 25944 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_278
timestamp 1644511149
transform 1 0 26680 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_281
timestamp 1644511149
transform 1 0 26956 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_296
timestamp 1644511149
transform 1 0 28336 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_21_306
timestamp 1644511149
transform 1 0 29256 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_318
timestamp 1644511149
transform 1 0 30360 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_330
timestamp 1644511149
transform 1 0 31464 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_21_337
timestamp 1644511149
transform 1 0 32108 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_349
timestamp 1644511149
transform 1 0 33212 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_361
timestamp 1644511149
transform 1 0 34316 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_373
timestamp 1644511149
transform 1 0 35420 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_385
timestamp 1644511149
transform 1 0 36524 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_391
timestamp 1644511149
transform 1 0 37076 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_393
timestamp 1644511149
transform 1 0 37260 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_405
timestamp 1644511149
transform 1 0 38364 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_417
timestamp 1644511149
transform 1 0 39468 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_429
timestamp 1644511149
transform 1 0 40572 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_441
timestamp 1644511149
transform 1 0 41676 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_447
timestamp 1644511149
transform 1 0 42228 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_449
timestamp 1644511149
transform 1 0 42412 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_461
timestamp 1644511149
transform 1 0 43516 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_473
timestamp 1644511149
transform 1 0 44620 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_21_500
timestamp 1644511149
transform 1 0 47104 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_508
timestamp 1644511149
transform 1 0 47840 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_22_3
timestamp 1644511149
transform 1 0 1380 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_10
timestamp 1644511149
transform 1 0 2024 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_17
timestamp 1644511149
transform 1 0 2668 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_25
timestamp 1644511149
transform 1 0 3404 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_29
timestamp 1644511149
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_41
timestamp 1644511149
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_53
timestamp 1644511149
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_65
timestamp 1644511149
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_77
timestamp 1644511149
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1644511149
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_85
timestamp 1644511149
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_97
timestamp 1644511149
transform 1 0 10028 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_109
timestamp 1644511149
transform 1 0 11132 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_121
timestamp 1644511149
transform 1 0 12236 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_133
timestamp 1644511149
transform 1 0 13340 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_139
timestamp 1644511149
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_141
timestamp 1644511149
transform 1 0 14076 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_153
timestamp 1644511149
transform 1 0 15180 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_165
timestamp 1644511149
transform 1 0 16284 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_177
timestamp 1644511149
transform 1 0 17388 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_185
timestamp 1644511149
transform 1 0 18124 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_192
timestamp 1644511149
transform 1 0 18768 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_206
timestamp 1644511149
transform 1 0 20056 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_218
timestamp 1644511149
transform 1 0 21160 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_230
timestamp 1644511149
transform 1 0 22264 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_242
timestamp 1644511149
transform 1 0 23368 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_250
timestamp 1644511149
transform 1 0 24104 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_22_253
timestamp 1644511149
transform 1 0 24380 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_22_270
timestamp 1644511149
transform 1 0 25944 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_278
timestamp 1644511149
transform 1 0 26680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_285
timestamp 1644511149
transform 1 0 27324 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_293
timestamp 1644511149
transform 1 0 28060 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_22_305
timestamp 1644511149
transform 1 0 29164 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_309
timestamp 1644511149
transform 1 0 29532 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_321
timestamp 1644511149
transform 1 0 30636 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_22_333
timestamp 1644511149
transform 1 0 31740 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_345
timestamp 1644511149
transform 1 0 32844 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_357
timestamp 1644511149
transform 1 0 33948 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_363
timestamp 1644511149
transform 1 0 34500 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_365
timestamp 1644511149
transform 1 0 34684 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_377
timestamp 1644511149
transform 1 0 35788 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_389
timestamp 1644511149
transform 1 0 36892 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_401
timestamp 1644511149
transform 1 0 37996 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_413
timestamp 1644511149
transform 1 0 39100 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_419
timestamp 1644511149
transform 1 0 39652 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_421
timestamp 1644511149
transform 1 0 39836 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_433
timestamp 1644511149
transform 1 0 40940 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_445
timestamp 1644511149
transform 1 0 42044 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_457
timestamp 1644511149
transform 1 0 43148 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_469
timestamp 1644511149
transform 1 0 44252 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_475
timestamp 1644511149
transform 1 0 44804 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_477
timestamp 1644511149
transform 1 0 44988 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_483
timestamp 1644511149
transform 1 0 45540 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_487
timestamp 1644511149
transform 1 0 45908 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_512
timestamp 1644511149
transform 1 0 48208 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_3
timestamp 1644511149
transform 1 0 1380 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_9
timestamp 1644511149
transform 1 0 1932 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_31
timestamp 1644511149
transform 1 0 3956 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_43
timestamp 1644511149
transform 1 0 5060 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1644511149
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_57
timestamp 1644511149
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_69
timestamp 1644511149
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_81
timestamp 1644511149
transform 1 0 8556 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_93
timestamp 1644511149
transform 1 0 9660 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_105
timestamp 1644511149
transform 1 0 10764 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp 1644511149
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_23_113
timestamp 1644511149
transform 1 0 11500 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_119
timestamp 1644511149
transform 1 0 12052 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_126
timestamp 1644511149
transform 1 0 12696 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_138
timestamp 1644511149
transform 1 0 13800 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_150
timestamp 1644511149
transform 1 0 14904 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_162
timestamp 1644511149
transform 1 0 16008 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_23_169
timestamp 1644511149
transform 1 0 16652 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_23_181
timestamp 1644511149
transform 1 0 17756 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_190
timestamp 1644511149
transform 1 0 18584 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_205
timestamp 1644511149
transform 1 0 19964 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_215
timestamp 1644511149
transform 1 0 20884 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_223
timestamp 1644511149
transform 1 0 21620 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_225
timestamp 1644511149
transform 1 0 21804 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_237
timestamp 1644511149
transform 1 0 22908 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_249
timestamp 1644511149
transform 1 0 24012 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_257
timestamp 1644511149
transform 1 0 24748 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_272
timestamp 1644511149
transform 1 0 26128 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_23_285
timestamp 1644511149
transform 1 0 27324 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_289
timestamp 1644511149
transform 1 0 27692 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_296
timestamp 1644511149
transform 1 0 28336 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_306
timestamp 1644511149
transform 1 0 29256 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_318
timestamp 1644511149
transform 1 0 30360 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_322
timestamp 1644511149
transform 1 0 30728 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_332
timestamp 1644511149
transform 1 0 31648 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_343
timestamp 1644511149
transform 1 0 32660 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_355
timestamp 1644511149
transform 1 0 33764 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_367
timestamp 1644511149
transform 1 0 34868 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_375
timestamp 1644511149
transform 1 0 35604 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_23_380
timestamp 1644511149
transform 1 0 36064 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_393
timestamp 1644511149
transform 1 0 37260 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_405
timestamp 1644511149
transform 1 0 38364 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_417
timestamp 1644511149
transform 1 0 39468 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_429
timestamp 1644511149
transform 1 0 40572 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_441
timestamp 1644511149
transform 1 0 41676 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_447
timestamp 1644511149
transform 1 0 42228 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_449
timestamp 1644511149
transform 1 0 42412 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_461
timestamp 1644511149
transform 1 0 43516 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_473
timestamp 1644511149
transform 1 0 44620 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_481
timestamp 1644511149
transform 1 0 45356 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_486
timestamp 1644511149
transform 1 0 45816 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_493
timestamp 1644511149
transform 1 0 46460 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_500
timestamp 1644511149
transform 1 0 47104 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_508
timestamp 1644511149
transform 1 0 47840 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_24_3
timestamp 1644511149
transform 1 0 1380 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_11
timestamp 1644511149
transform 1 0 2116 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_24_16
timestamp 1644511149
transform 1 0 2576 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_29
timestamp 1644511149
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_41
timestamp 1644511149
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_53
timestamp 1644511149
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_65
timestamp 1644511149
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_77
timestamp 1644511149
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1644511149
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_85
timestamp 1644511149
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_97
timestamp 1644511149
transform 1 0 10028 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_109
timestamp 1644511149
transform 1 0 11132 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_24_136
timestamp 1644511149
transform 1 0 13616 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_141
timestamp 1644511149
transform 1 0 14076 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_24_153
timestamp 1644511149
transform 1 0 15180 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_159
timestamp 1644511149
transform 1 0 15732 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_184
timestamp 1644511149
transform 1 0 18032 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_191
timestamp 1644511149
transform 1 0 18676 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_195
timestamp 1644511149
transform 1 0 19044 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_206
timestamp 1644511149
transform 1 0 20056 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_218
timestamp 1644511149
transform 1 0 21160 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_230
timestamp 1644511149
transform 1 0 22264 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_242
timestamp 1644511149
transform 1 0 23368 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_250
timestamp 1644511149
transform 1 0 24104 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_253
timestamp 1644511149
transform 1 0 24380 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_258
timestamp 1644511149
transform 1 0 24840 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_283
timestamp 1644511149
transform 1 0 27140 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_295
timestamp 1644511149
transform 1 0 28244 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_299
timestamp 1644511149
transform 1 0 28612 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_307
timestamp 1644511149
transform 1 0 29348 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_309
timestamp 1644511149
transform 1 0 29532 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_321
timestamp 1644511149
transform 1 0 30636 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_333
timestamp 1644511149
transform 1 0 31740 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_345
timestamp 1644511149
transform 1 0 32844 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_357
timestamp 1644511149
transform 1 0 33948 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_363
timestamp 1644511149
transform 1 0 34500 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_365
timestamp 1644511149
transform 1 0 34684 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_373
timestamp 1644511149
transform 1 0 35420 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_24_396
timestamp 1644511149
transform 1 0 37536 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_408
timestamp 1644511149
transform 1 0 38640 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_421
timestamp 1644511149
transform 1 0 39836 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_428
timestamp 1644511149
transform 1 0 40480 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_453
timestamp 1644511149
transform 1 0 42780 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_457
timestamp 1644511149
transform 1 0 43148 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_461
timestamp 1644511149
transform 1 0 43516 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_24_473
timestamp 1644511149
transform 1 0 44620 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_477
timestamp 1644511149
transform 1 0 44988 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_482
timestamp 1644511149
transform 1 0 45448 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_490
timestamp 1644511149
transform 1 0 46184 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_512
timestamp 1644511149
transform 1 0 48208 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_3
timestamp 1644511149
transform 1 0 1380 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_9
timestamp 1644511149
transform 1 0 1932 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_13
timestamp 1644511149
transform 1 0 2300 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_25
timestamp 1644511149
transform 1 0 3404 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_37
timestamp 1644511149
transform 1 0 4508 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_49
timestamp 1644511149
transform 1 0 5612 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_55
timestamp 1644511149
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_57
timestamp 1644511149
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_69
timestamp 1644511149
transform 1 0 7452 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_25_76
timestamp 1644511149
transform 1 0 8096 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_88
timestamp 1644511149
transform 1 0 9200 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_96
timestamp 1644511149
transform 1 0 9936 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_25_102
timestamp 1644511149
transform 1 0 10488 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_110
timestamp 1644511149
transform 1 0 11224 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_113
timestamp 1644511149
transform 1 0 11500 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_118
timestamp 1644511149
transform 1 0 11960 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_25_143
timestamp 1644511149
transform 1 0 14260 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_25_155
timestamp 1644511149
transform 1 0 15364 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_25_161
timestamp 1644511149
transform 1 0 15916 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_167
timestamp 1644511149
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_172
timestamp 1644511149
transform 1 0 16928 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_184
timestamp 1644511149
transform 1 0 18032 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_25_207
timestamp 1644511149
transform 1 0 20148 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_219
timestamp 1644511149
transform 1 0 21252 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_223
timestamp 1644511149
transform 1 0 21620 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_225
timestamp 1644511149
transform 1 0 21804 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_237
timestamp 1644511149
transform 1 0 22908 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_245
timestamp 1644511149
transform 1 0 23644 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_250
timestamp 1644511149
transform 1 0 24104 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_257
timestamp 1644511149
transform 1 0 24748 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_267
timestamp 1644511149
transform 1 0 25668 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_274
timestamp 1644511149
transform 1 0 26312 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_25_284
timestamp 1644511149
transform 1 0 27232 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_296
timestamp 1644511149
transform 1 0 28336 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_300
timestamp 1644511149
transform 1 0 28704 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_25_322
timestamp 1644511149
transform 1 0 30728 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_328
timestamp 1644511149
transform 1 0 31280 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_332
timestamp 1644511149
transform 1 0 31648 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_337
timestamp 1644511149
transform 1 0 32108 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_342
timestamp 1644511149
transform 1 0 32568 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_349
timestamp 1644511149
transform 1 0 33212 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_25_358
timestamp 1644511149
transform 1 0 34040 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_365
timestamp 1644511149
transform 1 0 34684 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_369
timestamp 1644511149
transform 1 0 35052 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_373
timestamp 1644511149
transform 1 0 35420 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_380
timestamp 1644511149
transform 1 0 36064 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_387
timestamp 1644511149
transform 1 0 36708 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_391
timestamp 1644511149
transform 1 0 37076 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_396
timestamp 1644511149
transform 1 0 37536 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_25_408
timestamp 1644511149
transform 1 0 38640 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_432
timestamp 1644511149
transform 1 0 40848 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_439
timestamp 1644511149
transform 1 0 41492 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_447
timestamp 1644511149
transform 1 0 42228 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_25_449
timestamp 1644511149
transform 1 0 42412 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_25_453
timestamp 1644511149
transform 1 0 42780 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_25_462
timestamp 1644511149
transform 1 0 43608 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_470
timestamp 1644511149
transform 1 0 44344 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_475
timestamp 1644511149
transform 1 0 44804 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_500
timestamp 1644511149
transform 1 0 47104 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_508
timestamp 1644511149
transform 1 0 47840 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_26_3
timestamp 1644511149
transform 1 0 1380 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_11
timestamp 1644511149
transform 1 0 2116 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_15
timestamp 1644511149
transform 1 0 2484 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_22
timestamp 1644511149
transform 1 0 3128 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_26_29
timestamp 1644511149
transform 1 0 3772 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_26_38
timestamp 1644511149
transform 1 0 4600 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_45
timestamp 1644511149
transform 1 0 5244 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_26_57
timestamp 1644511149
transform 1 0 6348 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_62
timestamp 1644511149
transform 1 0 6808 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_69
timestamp 1644511149
transform 1 0 7452 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_76
timestamp 1644511149
transform 1 0 8096 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_26_85
timestamp 1644511149
transform 1 0 8924 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_26_94
timestamp 1644511149
transform 1 0 9752 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_119
timestamp 1644511149
transform 1 0 12052 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_126
timestamp 1644511149
transform 1 0 12696 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_132
timestamp 1644511149
transform 1 0 13248 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_136
timestamp 1644511149
transform 1 0 13616 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_141
timestamp 1644511149
transform 1 0 14076 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_149
timestamp 1644511149
transform 1 0 14812 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_153
timestamp 1644511149
transform 1 0 15180 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_178
timestamp 1644511149
transform 1 0 17480 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_185
timestamp 1644511149
transform 1 0 18124 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_192
timestamp 1644511149
transform 1 0 18768 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_197
timestamp 1644511149
transform 1 0 19228 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_201
timestamp 1644511149
transform 1 0 19596 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_226
timestamp 1644511149
transform 1 0 21896 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_233
timestamp 1644511149
transform 1 0 22540 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_248
timestamp 1644511149
transform 1 0 23920 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_256
timestamp 1644511149
transform 1 0 24656 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_26_283
timestamp 1644511149
transform 1 0 27140 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_290
timestamp 1644511149
transform 1 0 27784 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_297
timestamp 1644511149
transform 1 0 28428 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_304
timestamp 1644511149
transform 1 0 29072 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_309
timestamp 1644511149
transform 1 0 29532 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_316
timestamp 1644511149
transform 1 0 30176 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_323
timestamp 1644511149
transform 1 0 30820 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_26_334
timestamp 1644511149
transform 1 0 31832 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_359
timestamp 1644511149
transform 1 0 34132 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_363
timestamp 1644511149
transform 1 0 34500 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_365
timestamp 1644511149
transform 1 0 34684 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_390
timestamp 1644511149
transform 1 0 36984 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_397
timestamp 1644511149
transform 1 0 37628 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_405
timestamp 1644511149
transform 1 0 38364 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_409
timestamp 1644511149
transform 1 0 38732 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_416
timestamp 1644511149
transform 1 0 39376 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_424
timestamp 1644511149
transform 1 0 40112 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_431
timestamp 1644511149
transform 1 0 40756 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_443
timestamp 1644511149
transform 1 0 41860 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_447
timestamp 1644511149
transform 1 0 42228 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_472
timestamp 1644511149
transform 1 0 44528 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_480
timestamp 1644511149
transform 1 0 45264 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_487
timestamp 1644511149
transform 1 0 45908 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_512
timestamp 1644511149
transform 1 0 48208 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_24
timestamp 1644511149
transform 1 0 3312 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_29
timestamp 1644511149
transform 1 0 3772 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_52
timestamp 1644511149
transform 1 0 5888 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_57
timestamp 1644511149
transform 1 0 6348 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_80
timestamp 1644511149
transform 1 0 8464 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_27_106
timestamp 1644511149
transform 1 0 10856 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_27_113
timestamp 1644511149
transform 1 0 11500 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_27_121
timestamp 1644511149
transform 1 0 12236 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_27_130
timestamp 1644511149
transform 1 0 13064 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_138
timestamp 1644511149
transform 1 0 13800 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_27_162
timestamp 1644511149
transform 1 0 16008 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_27_169
timestamp 1644511149
transform 1 0 16652 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_192
timestamp 1644511149
transform 1 0 18768 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_200
timestamp 1644511149
transform 1 0 19504 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_204
timestamp 1644511149
transform 1 0 19872 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_208
timestamp 1644511149
transform 1 0 20240 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_216
timestamp 1644511149
transform 1 0 20976 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_220
timestamp 1644511149
transform 1 0 21344 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_225
timestamp 1644511149
transform 1 0 21804 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_248
timestamp 1644511149
transform 1 0 23920 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_27_274
timestamp 1644511149
transform 1 0 26312 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_27_281
timestamp 1644511149
transform 1 0 26956 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_304
timestamp 1644511149
transform 1 0 29072 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_309
timestamp 1644511149
transform 1 0 29532 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_332
timestamp 1644511149
transform 1 0 31648 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_27_358
timestamp 1644511149
transform 1 0 34040 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_27_386
timestamp 1644511149
transform 1 0 36616 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_27_414
timestamp 1644511149
transform 1 0 39192 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_421
timestamp 1644511149
transform 1 0 39836 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_443
timestamp 1644511149
transform 1 0 41860 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_447
timestamp 1644511149
transform 1 0 42228 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_449
timestamp 1644511149
transform 1 0 42412 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_471
timestamp 1644511149
transform 1 0 44436 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_475
timestamp 1644511149
transform 1 0 44804 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_477
timestamp 1644511149
transform 1 0 44988 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_500
timestamp 1644511149
transform 1 0 47104 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_508
timestamp 1644511149
transform 1 0 47840 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1644511149
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1644511149
transform -1 0 48852 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1644511149
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1644511149
transform -1 0 48852 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1644511149
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1644511149
transform -1 0 48852 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1644511149
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1644511149
transform -1 0 48852 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1644511149
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1644511149
transform -1 0 48852 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1644511149
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1644511149
transform -1 0 48852 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1644511149
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1644511149
transform -1 0 48852 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1644511149
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1644511149
transform -1 0 48852 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1644511149
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1644511149
transform -1 0 48852 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1644511149
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1644511149
transform -1 0 48852 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1644511149
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1644511149
transform -1 0 48852 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1644511149
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1644511149
transform -1 0 48852 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1644511149
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1644511149
transform -1 0 48852 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1644511149
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1644511149
transform -1 0 48852 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1644511149
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1644511149
transform -1 0 48852 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1644511149
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1644511149
transform -1 0 48852 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1644511149
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1644511149
transform -1 0 48852 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1644511149
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1644511149
transform -1 0 48852 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1644511149
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1644511149
transform -1 0 48852 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1644511149
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1644511149
transform -1 0 48852 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1644511149
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1644511149
transform -1 0 48852 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1644511149
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1644511149
transform -1 0 48852 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1644511149
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1644511149
transform -1 0 48852 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1644511149
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1644511149
transform -1 0 48852 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1644511149
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1644511149
transform -1 0 48852 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1644511149
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1644511149
transform -1 0 48852 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1644511149
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1644511149
transform -1 0 48852 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1644511149
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1644511149
transform -1 0 48852 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_56 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_57
timestamp 1644511149
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_58
timestamp 1644511149
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_59
timestamp 1644511149
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_60
timestamp 1644511149
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_61
timestamp 1644511149
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_62
timestamp 1644511149
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_63
timestamp 1644511149
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_64
timestamp 1644511149
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_65
timestamp 1644511149
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_66
timestamp 1644511149
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_67
timestamp 1644511149
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_68
timestamp 1644511149
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_69
timestamp 1644511149
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_70
timestamp 1644511149
transform 1 0 39744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_71
timestamp 1644511149
transform 1 0 42320 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72
timestamp 1644511149
transform 1 0 44896 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 1644511149
transform 1 0 47472 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74
timestamp 1644511149
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 1644511149
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 1644511149
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 1644511149
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 1644511149
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 1644511149
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 1644511149
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1644511149
transform 1 0 42320 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1644511149
transform 1 0 47472 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1644511149
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1644511149
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1644511149
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1644511149
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1644511149
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1644511149
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1644511149
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1644511149
transform 1 0 39744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1644511149
transform 1 0 44896 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1644511149
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1644511149
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1644511149
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1644511149
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1644511149
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1644511149
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1644511149
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1644511149
transform 1 0 42320 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1644511149
transform 1 0 47472 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1644511149
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1644511149
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1644511149
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1644511149
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1644511149
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1644511149
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1644511149
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1644511149
transform 1 0 39744 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1644511149
transform 1 0 44896 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1644511149
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1644511149
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1644511149
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1644511149
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1644511149
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1644511149
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1644511149
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1644511149
transform 1 0 42320 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1644511149
transform 1 0 47472 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1644511149
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1644511149
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1644511149
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1644511149
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1644511149
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1644511149
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1644511149
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1644511149
transform 1 0 39744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1644511149
transform 1 0 44896 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1644511149
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1644511149
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1644511149
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1644511149
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1644511149
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1644511149
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1644511149
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1644511149
transform 1 0 42320 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1644511149
transform 1 0 47472 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1644511149
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1644511149
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1644511149
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1644511149
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1644511149
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1644511149
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1644511149
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1644511149
transform 1 0 39744 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1644511149
transform 1 0 44896 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1644511149
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1644511149
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1644511149
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1644511149
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1644511149
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1644511149
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1644511149
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1644511149
transform 1 0 42320 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1644511149
transform 1 0 47472 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1644511149
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1644511149
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1644511149
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1644511149
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1644511149
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1644511149
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1644511149
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1644511149
transform 1 0 39744 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1644511149
transform 1 0 44896 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1644511149
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1644511149
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1644511149
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1644511149
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1644511149
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1644511149
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1644511149
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1644511149
transform 1 0 42320 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1644511149
transform 1 0 47472 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1644511149
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1644511149
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1644511149
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1644511149
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1644511149
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1644511149
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1644511149
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1644511149
transform 1 0 39744 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1644511149
transform 1 0 44896 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1644511149
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1644511149
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1644511149
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1644511149
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1644511149
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1644511149
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1644511149
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1644511149
transform 1 0 42320 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1644511149
transform 1 0 47472 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1644511149
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1644511149
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1644511149
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1644511149
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1644511149
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1644511149
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1644511149
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1644511149
transform 1 0 39744 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1644511149
transform 1 0 44896 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1644511149
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1644511149
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1644511149
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1644511149
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1644511149
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1644511149
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1644511149
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1644511149
transform 1 0 42320 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1644511149
transform 1 0 47472 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1644511149
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1644511149
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1644511149
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1644511149
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1644511149
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1644511149
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1644511149
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1644511149
transform 1 0 39744 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1644511149
transform 1 0 44896 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1644511149
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1644511149
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1644511149
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1644511149
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1644511149
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1644511149
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1644511149
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1644511149
transform 1 0 42320 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1644511149
transform 1 0 47472 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1644511149
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1644511149
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1644511149
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1644511149
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1644511149
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1644511149
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1644511149
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1644511149
transform 1 0 39744 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1644511149
transform 1 0 44896 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1644511149
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1644511149
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1644511149
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1644511149
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1644511149
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1644511149
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1644511149
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1644511149
transform 1 0 42320 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1644511149
transform 1 0 47472 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1644511149
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1644511149
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1644511149
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1644511149
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1644511149
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1644511149
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1644511149
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1644511149
transform 1 0 39744 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1644511149
transform 1 0 44896 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1644511149
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1644511149
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1644511149
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1644511149
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1644511149
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1644511149
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1644511149
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1644511149
transform 1 0 42320 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1644511149
transform 1 0 47472 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1644511149
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1644511149
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1644511149
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1644511149
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1644511149
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1644511149
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1644511149
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1644511149
transform 1 0 39744 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1644511149
transform 1 0 44896 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1644511149
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1644511149
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1644511149
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1644511149
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1644511149
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1644511149
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1644511149
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1644511149
transform 1 0 42320 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1644511149
transform 1 0 47472 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1644511149
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1644511149
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1644511149
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1644511149
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1644511149
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1644511149
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1644511149
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1644511149
transform 1 0 39744 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1644511149
transform 1 0 44896 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1644511149
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1644511149
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1644511149
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1644511149
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1644511149
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1644511149
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1644511149
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1644511149
transform 1 0 42320 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1644511149
transform 1 0 47472 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1644511149
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1644511149
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1644511149
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1644511149
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1644511149
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1644511149
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1644511149
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1644511149
transform 1 0 39744 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1644511149
transform 1 0 44896 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1644511149
transform 1 0 3680 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1644511149
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1644511149
transform 1 0 8832 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1644511149
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1644511149
transform 1 0 13984 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1644511149
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1644511149
transform 1 0 19136 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1644511149
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1644511149
transform 1 0 24288 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1644511149
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1644511149
transform 1 0 29440 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1644511149
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1644511149
transform 1 0 34592 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1644511149
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1644511149
transform 1 0 39744 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1644511149
transform 1 0 42320 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1644511149
transform 1 0 44896 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1644511149
transform 1 0 47472 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _242_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 26956 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _243_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 28336 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _244_
timestamp 1644511149
transform 1 0 7728 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _245_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 10396 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _246_
timestamp 1644511149
transform 1 0 14260 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _247_
timestamp 1644511149
transform -1 0 2760 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _248_
timestamp 1644511149
transform 1 0 20424 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _249_
timestamp 1644511149
transform -1 0 2668 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _250_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 26956 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _251_
timestamp 1644511149
transform 1 0 47564 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _252_
timestamp 1644511149
transform -1 0 25576 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _253_
timestamp 1644511149
transform 1 0 47564 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _254_
timestamp 1644511149
transform 1 0 47564 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _255_
timestamp 1644511149
transform 1 0 42504 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _256_
timestamp 1644511149
transform 1 0 24472 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  _257_
timestamp 1644511149
transform -1 0 24748 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _258_
timestamp 1644511149
transform 1 0 15824 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _259_
timestamp 1644511149
transform 1 0 38456 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _260_
timestamp 1644511149
transform -1 0 18124 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _261_
timestamp 1644511149
transform 1 0 33764 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _262_
timestamp 1644511149
transform -1 0 15180 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _263_
timestamp 1644511149
transform 1 0 25116 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _264_
timestamp 1644511149
transform -1 0 45264 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _265_
timestamp 1644511149
transform 1 0 47564 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _266_
timestamp 1644511149
transform -1 0 18676 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _267_
timestamp 1644511149
transform 1 0 47564 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _268_
timestamp 1644511149
transform -1 0 18400 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _269_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 25116 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _270_
timestamp 1644511149
transform 1 0 46828 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _271_
timestamp 1644511149
transform -1 0 36064 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _272_
timestamp 1644511149
transform 1 0 8188 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _273_
timestamp 1644511149
transform -1 0 46828 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _274_
timestamp 1644511149
transform -1 0 4048 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_8  _275_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 25116 0 -1 15232
box -38 -48 1050 592
use sky130_fd_sc_hd__inv_2  _276_
timestamp 1644511149
transform 1 0 37260 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _277_
timestamp 1644511149
transform 1 0 12420 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _278_
timestamp 1644511149
transform 1 0 31096 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _279_
timestamp 1644511149
transform -1 0 6992 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _280_
timestamp 1644511149
transform 1 0 38456 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _281_
timestamp 1644511149
transform 1 0 25116 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _282_
timestamp 1644511149
transform 1 0 47564 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _283_
timestamp 1644511149
transform 1 0 10212 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _284_
timestamp 1644511149
transform -1 0 30176 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _285_
timestamp 1644511149
transform -1 0 5704 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _286_
timestamp 1644511149
transform 1 0 47564 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _287_
timestamp 1644511149
transform -1 0 18768 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  _288_
timestamp 1644511149
transform -1 0 18584 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _289_
timestamp 1644511149
transform 1 0 27508 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _290_
timestamp 1644511149
transform -1 0 2668 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _291_
timestamp 1644511149
transform -1 0 13616 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _292_
timestamp 1644511149
transform -1 0 2668 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _293_
timestamp 1644511149
transform 1 0 7820 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_8  _294_
timestamp 1644511149
transform 1 0 18952 0 -1 15232
box -38 -48 1050 592
use sky130_fd_sc_hd__inv_2  _295_
timestamp 1644511149
transform -1 0 43332 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _296_
timestamp 1644511149
transform 1 0 44988 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _297_
timestamp 1644511149
transform 1 0 32108 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _298_
timestamp 1644511149
transform -1 0 13616 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _299_
timestamp 1644511149
transform 1 0 42504 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _300_
timestamp 1644511149
transform -1 0 20056 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _301_
timestamp 1644511149
transform -1 0 8096 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _302_
timestamp 1644511149
transform -1 0 22632 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _303_
timestamp 1644511149
transform 1 0 39836 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _304_
timestamp 1644511149
transform 1 0 18124 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _305_
timestamp 1644511149
transform 1 0 39836 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _306_
timestamp 1644511149
transform -1 0 20056 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _307_
timestamp 1644511149
transform -1 0 2300 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _308_
timestamp 1644511149
transform 1 0 40204 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _309_
timestamp 1644511149
transform 1 0 11684 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _310_
timestamp 1644511149
transform 1 0 35880 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _311_
timestamp 1644511149
transform -1 0 4048 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _312_
timestamp 1644511149
transform 1 0 20332 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _313_
timestamp 1644511149
transform -1 0 11776 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _314_
timestamp 1644511149
transform 1 0 11776 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _315_
timestamp 1644511149
transform 1 0 40020 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _316_
timestamp 1644511149
transform 1 0 47564 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _317_
timestamp 1644511149
transform -1 0 46736 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _318_
timestamp 1644511149
transform 1 0 27692 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  _319_
timestamp 1644511149
transform -1 0 27324 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _320_
timestamp 1644511149
transform -1 0 26312 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _321_
timestamp 1644511149
transform 1 0 45172 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _322_
timestamp 1644511149
transform 1 0 26956 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _323_
timestamp 1644511149
transform -1 0 43608 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _324_
timestamp 1644511149
transform -1 0 24932 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_8  _325_
timestamp 1644511149
transform 1 0 27324 0 -1 14144
box -38 -48 1050 592
use sky130_fd_sc_hd__inv_2  _326_
timestamp 1644511149
transform 1 0 34684 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _327_
timestamp 1644511149
transform -1 0 4600 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _328_
timestamp 1644511149
transform 1 0 34684 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _329_
timestamp 1644511149
transform -1 0 22540 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _330_
timestamp 1644511149
transform -1 0 4692 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _331_
timestamp 1644511149
transform -1 0 27784 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _332_
timestamp 1644511149
transform 1 0 8188 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _333_
timestamp 1644511149
transform -1 0 4048 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _334_
timestamp 1644511149
transform 1 0 45172 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _335_
timestamp 1644511149
transform 1 0 45448 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _336_
timestamp 1644511149
transform 1 0 42320 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _337_
timestamp 1644511149
transform 1 0 26772 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _338_
timestamp 1644511149
transform -1 0 6992 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _339_
timestamp 1644511149
transform 1 0 24380 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _340_
timestamp 1644511149
transform 1 0 36524 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _341_
timestamp 1644511149
transform 1 0 9200 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _342_
timestamp 1644511149
transform 1 0 37352 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _343_
timestamp 1644511149
transform 1 0 28704 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _344_
timestamp 1644511149
transform 1 0 24472 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _345_
timestamp 1644511149
transform 1 0 31372 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _346_
timestamp 1644511149
transform 1 0 15640 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _347_
timestamp 1644511149
transform -1 0 12696 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _348_
timestamp 1644511149
transform 1 0 31556 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _349_
timestamp 1644511149
transform 1 0 32108 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _350_
timestamp 1644511149
transform -1 0 32568 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _351_
timestamp 1644511149
transform 1 0 33028 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _352_
timestamp 1644511149
transform 1 0 47564 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _353_
timestamp 1644511149
transform 1 0 35144 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _354_
timestamp 1644511149
transform 1 0 47564 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _355_
timestamp 1644511149
transform 1 0 28704 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _356_
timestamp 1644511149
transform 1 0 15916 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _357_
timestamp 1644511149
transform 1 0 28152 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _358_
timestamp 1644511149
transform 1 0 29072 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _359_
timestamp 1644511149
transform -1 0 15732 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _360_
timestamp 1644511149
transform 1 0 29532 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _361_
timestamp 1644511149
transform -1 0 31740 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _362_
timestamp 1644511149
transform -1 0 2484 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _363_
timestamp 1644511149
transform 1 0 33212 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _364_
timestamp 1644511149
transform 1 0 19964 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _365_
timestamp 1644511149
transform -1 0 2576 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _366_
timestamp 1644511149
transform -1 0 2484 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _367_
timestamp 1644511149
transform 1 0 30820 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _368_
timestamp 1644511149
transform -1 0 2668 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _369_
timestamp 1644511149
transform -1 0 2668 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _370_
timestamp 1644511149
transform 1 0 27968 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _371_
timestamp 1644511149
transform 1 0 47564 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _372_
timestamp 1644511149
transform 1 0 45632 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _373_
timestamp 1644511149
transform 1 0 19228 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _374_
timestamp 1644511149
transform 1 0 28336 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _375_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 41952 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _376_
timestamp 1644511149
transform -1 0 5888 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _377_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 42044 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _378__2 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 5980 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _379__3
timestamp 1644511149
transform -1 0 10672 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _380__4
timestamp 1644511149
transform -1 0 14536 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _381__5
timestamp 1644511149
transform -1 0 2484 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _382__6
timestamp 1644511149
transform 1 0 21068 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _383__7
timestamp 1644511149
transform 1 0 1472 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _384__8
timestamp 1644511149
transform -1 0 47840 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _385__9
timestamp 1644511149
transform 1 0 26220 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _386__10
timestamp 1644511149
transform 1 0 45632 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _387__11
timestamp 1644511149
transform 1 0 45264 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _388__12
timestamp 1644511149
transform -1 0 43976 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _389__13
timestamp 1644511149
transform -1 0 16008 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _390__14
timestamp 1644511149
transform -1 0 39376 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _391__15
timestamp 1644511149
transform -1 0 19504 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _392__16
timestamp 1644511149
transform 1 0 34408 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _393__17
timestamp 1644511149
transform 1 0 13616 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _394__18
timestamp 1644511149
transform 1 0 44528 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _395__19
timestamp 1644511149
transform 1 0 45816 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _396__20
timestamp 1644511149
transform -1 0 18768 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _397__21
timestamp 1644511149
transform 1 0 45632 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _398__22
timestamp 1644511149
transform -1 0 17940 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _399__23
timestamp 1644511149
transform 1 0 46184 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _400__24
timestamp 1644511149
transform -1 0 36064 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _401__25
timestamp 1644511149
transform 1 0 7544 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _402__26
timestamp 1644511149
transform -1 0 47012 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _403__27
timestamp 1644511149
transform -1 0 4692 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _404__28
timestamp 1644511149
transform -1 0 38456 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _405__29
timestamp 1644511149
transform -1 0 12696 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _406__30
timestamp 1644511149
transform 1 0 31096 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _407__31
timestamp 1644511149
transform 1 0 5612 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _408__32
timestamp 1644511149
transform -1 0 39376 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _409__33
timestamp 1644511149
transform 1 0 47564 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _410__34
timestamp 1644511149
transform -1 0 29072 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _411__35
timestamp 1644511149
transform -1 0 28428 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _412__36
timestamp 1644511149
transform -1 0 5244 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _413__37
timestamp 1644511149
transform 1 0 9476 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _414__38
timestamp 1644511149
transform 1 0 47472 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _415__39
timestamp 1644511149
transform -1 0 30820 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _416__40
timestamp 1644511149
transform 1 0 45632 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _417__41
timestamp 1644511149
transform 1 0 1748 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _418__42
timestamp 1644511149
transform -1 0 13248 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _419__43
timestamp 1644511149
transform -1 0 2392 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _420__44
timestamp 1644511149
transform -1 0 45908 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _421__45
timestamp 1644511149
transform -1 0 16928 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _422__46
timestamp 1644511149
transform 1 0 1748 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _423__47
timestamp 1644511149
transform -1 0 28152 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _424__48
timestamp 1644511149
transform 1 0 44988 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _425__49
timestamp 1644511149
transform 1 0 7176 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _426__50
timestamp 1644511149
transform 1 0 44528 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _427__51
timestamp 1644511149
transform -1 0 32292 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _428__52
timestamp 1644511149
transform 1 0 12788 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _429__53
timestamp 1644511149
transform 1 0 41952 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _430__54
timestamp 1644511149
transform -1 0 6808 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _431__55
timestamp 1644511149
transform 1 0 23000 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _432__56
timestamp 1644511149
transform -1 0 40204 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _433__57
timestamp 1644511149
transform 1 0 17480 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _434__58
timestamp 1644511149
transform -1 0 40756 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _435__59
timestamp 1644511149
transform -1 0 1748 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _436__60
timestamp 1644511149
transform -1 0 41492 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _437__61
timestamp 1644511149
transform -1 0 11960 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _438__62
timestamp 1644511149
transform -1 0 36156 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _439__63
timestamp 1644511149
transform 1 0 3036 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _440__64
timestamp 1644511149
transform -1 0 11776 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _441__65
timestamp 1644511149
transform -1 0 11960 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _442__66
timestamp 1644511149
transform -1 0 40296 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _443__67
timestamp 1644511149
transform -1 0 45908 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _444__68
timestamp 1644511149
transform 1 0 44528 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _445__69
timestamp 1644511149
transform 1 0 23644 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _446__70
timestamp 1644511149
transform -1 0 45816 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _447__71
timestamp 1644511149
transform 1 0 19872 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _448__72
timestamp 1644511149
transform 1 0 26220 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _449__73
timestamp 1644511149
transform -1 0 43516 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _450__74
timestamp 1644511149
transform 1 0 23644 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _451__75
timestamp 1644511149
transform -1 0 35512 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _452__76
timestamp 1644511149
transform 1 0 4968 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _453__77
timestamp 1644511149
transform 1 0 33948 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _454__78
timestamp 1644511149
transform 1 0 21068 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _455__79
timestamp 1644511149
transform 1 0 3036 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _456__80
timestamp 1644511149
transform -1 0 9200 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _457__81
timestamp 1644511149
transform -1 0 4048 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _458__82
timestamp 1644511149
transform 1 0 44988 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _459__83
timestamp 1644511149
transform 1 0 43884 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _460__84
timestamp 1644511149
transform 1 0 41676 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _461__85
timestamp 1644511149
transform 1 0 5060 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _462__86
timestamp 1644511149
transform 1 0 23828 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _463__87
timestamp 1644511149
transform 1 0 36984 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _464__88
timestamp 1644511149
transform -1 0 10120 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _465__89
timestamp 1644511149
transform -1 0 37536 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _466__90
timestamp 1644511149
transform -1 0 27232 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _467__91
timestamp 1644511149
transform 1 0 31372 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _468__92
timestamp 1644511149
transform 1 0 14904 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _469__93
timestamp 1644511149
transform 1 0 12328 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _470__94
timestamp 1644511149
transform 1 0 31372 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _471__95
timestamp 1644511149
transform -1 0 33212 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _472__96
timestamp 1644511149
transform -1 0 33304 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _473__97
timestamp 1644511149
transform 1 0 44252 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _474__98
timestamp 1644511149
transform 1 0 36432 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _475__99
timestamp 1644511149
transform -1 0 29808 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _476__100
timestamp 1644511149
transform -1 0 30084 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _477__101
timestamp 1644511149
transform -1 0 16928 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _478__102
timestamp 1644511149
transform 1 0 28520 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _479__103
timestamp 1644511149
transform 1 0 2852 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _480__104
timestamp 1644511149
transform -1 0 33948 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _481__105
timestamp 1644511149
transform 1 0 19320 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _482__106
timestamp 1644511149
transform -1 0 2300 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _483__107
timestamp 1644511149
transform -1 0 2300 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _484__108
timestamp 1644511149
transform -1 0 2392 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _485_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 5704 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _486_
timestamp 1644511149
transform 1 0 10304 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _487_
timestamp 1644511149
transform 1 0 14168 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _488_
timestamp 1644511149
transform 1 0 2116 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _489_
timestamp 1644511149
transform -1 0 21344 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _490_
timestamp 1644511149
transform 1 0 2116 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _491_
timestamp 1644511149
transform -1 0 47104 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _492_
timestamp 1644511149
transform -1 0 26496 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _493_
timestamp 1644511149
transform 1 0 46276 0 1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _494_
timestamp 1644511149
transform 1 0 45908 0 1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _495_
timestamp 1644511149
transform 1 0 43148 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _496_
timestamp 1644511149
transform 1 0 15732 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _497_
timestamp 1644511149
transform 1 0 38916 0 -1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _498_
timestamp 1644511149
transform -1 0 18768 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _499_
timestamp 1644511149
transform 1 0 34684 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _500_
timestamp 1644511149
transform -1 0 15548 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _501_
timestamp 1644511149
transform 1 0 44712 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _502_
timestamp 1644511149
transform 1 0 46276 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _503_
timestamp 1644511149
transform 1 0 18216 0 -1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _504_
timestamp 1644511149
transform 1 0 46276 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _505_
timestamp 1644511149
transform 1 0 17664 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _506_
timestamp 1644511149
transform 1 0 46276 0 1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _507_
timestamp 1644511149
transform 1 0 35604 0 1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _508_
timestamp 1644511149
transform 1 0 8832 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _509_
timestamp 1644511149
transform 1 0 46276 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _510_
timestamp 1644511149
transform -1 0 4600 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _511_
timestamp 1644511149
transform 1 0 37260 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _512_
timestamp 1644511149
transform 1 0 12328 0 -1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _513_
timestamp 1644511149
transform 1 0 32108 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _514_
timestamp 1644511149
transform 1 0 6348 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _515_
timestamp 1644511149
transform 1 0 39100 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _516_
timestamp 1644511149
transform -1 0 48208 0 1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _517_
timestamp 1644511149
transform 1 0 28796 0 -1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _518_
timestamp 1644511149
transform 1 0 27140 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _519_
timestamp 1644511149
transform 1 0 4968 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _520_
timestamp 1644511149
transform 1 0 10120 0 1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _521_
timestamp 1644511149
transform -1 0 48208 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _522_
timestamp 1644511149
transform 1 0 29716 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _523_
timestamp 1644511149
transform 1 0 46276 0 1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _524_
timestamp 1644511149
transform 1 0 2024 0 -1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _525_
timestamp 1644511149
transform 1 0 12972 0 -1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _526_
timestamp 1644511149
transform 1 0 2024 0 -1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _527_
timestamp 1644511149
transform 1 0 45172 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _528_
timestamp 1644511149
transform 1 0 16652 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _529_
timestamp 1644511149
transform 1 0 2116 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _530_
timestamp 1644511149
transform 1 0 27876 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _531_
timestamp 1644511149
transform 1 0 46276 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _532_
timestamp 1644511149
transform 1 0 8924 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _533_
timestamp 1644511149
transform 1 0 42412 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _534_
timestamp 1644511149
transform 1 0 45172 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _535_
timestamp 1644511149
transform 1 0 32016 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _536_
timestamp 1644511149
transform 1 0 14076 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _537_
timestamp 1644511149
transform 1 0 42504 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _538_
timestamp 1644511149
transform 1 0 6532 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _539_
timestamp 1644511149
transform -1 0 23920 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _540_
timestamp 1644511149
transform 1 0 39928 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _541_
timestamp 1644511149
transform 1 0 18124 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _542_
timestamp 1644511149
transform 1 0 39928 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _543_
timestamp 1644511149
transform 1 0 1380 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _544_
timestamp 1644511149
transform 1 0 40848 0 1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _545_
timestamp 1644511149
transform 1 0 11592 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _546_
timestamp 1644511149
transform 1 0 35880 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _547_
timestamp 1644511149
transform -1 0 3312 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _548_
timestamp 1644511149
transform 1 0 11040 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _549_
timestamp 1644511149
transform 1 0 11684 0 1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _550_
timestamp 1644511149
transform 1 0 40020 0 -1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _551_
timestamp 1644511149
transform 1 0 45172 0 -1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _552_
timestamp 1644511149
transform 1 0 45172 0 -1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _553_
timestamp 1644511149
transform 1 0 25208 0 1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _554_
timestamp 1644511149
transform 1 0 45172 0 -1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _555_
timestamp 1644511149
transform -1 0 20148 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _556_
timestamp 1644511149
transform 1 0 26864 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _557_
timestamp 1644511149
transform 1 0 42596 0 1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _558_
timestamp 1644511149
transform 1 0 23920 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _559_
timestamp 1644511149
transform 1 0 34868 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _560_
timestamp 1644511149
transform -1 0 5888 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _561_
timestamp 1644511149
transform 1 0 34684 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _562_
timestamp 1644511149
transform 1 0 21988 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _563_
timestamp 1644511149
transform 1 0 3772 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _564_
timestamp 1644511149
transform 1 0 8924 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _565_
timestamp 1644511149
transform 1 0 3772 0 1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _566_
timestamp 1644511149
transform 1 0 45172 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _567_
timestamp 1644511149
transform -1 0 44528 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _568_
timestamp 1644511149
transform 1 0 42412 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _569_
timestamp 1644511149
transform 1 0 6348 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _570_
timestamp 1644511149
transform 1 0 24380 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _571_
timestamp 1644511149
transform 1 0 37260 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _572_
timestamp 1644511149
transform 1 0 9108 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _573_
timestamp 1644511149
transform 1 0 37260 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _574_
timestamp 1644511149
transform -1 0 27140 0 1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _575_
timestamp 1644511149
transform 1 0 32108 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _576_
timestamp 1644511149
transform 1 0 15548 0 1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _577_
timestamp 1644511149
transform -1 0 13616 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _578_
timestamp 1644511149
transform 1 0 32108 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _579_
timestamp 1644511149
transform 1 0 32200 0 1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _580_
timestamp 1644511149
transform 1 0 32936 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _581_
timestamp 1644511149
transform 1 0 45172 0 -1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _582_
timestamp 1644511149
transform -1 0 36984 0 1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _583_
timestamp 1644511149
transform 1 0 28796 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _584_
timestamp 1644511149
transform 1 0 29716 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _585_
timestamp 1644511149
transform 1 0 16100 0 1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _586_
timestamp 1644511149
transform -1 0 29072 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _587_
timestamp 1644511149
transform -1 0 3312 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _588_
timestamp 1644511149
transform 1 0 33672 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _589_
timestamp 1644511149
transform 1 0 19964 0 1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _590_
timestamp 1644511149
transform 1 0 2024 0 -1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _591_
timestamp 1644511149
transform 1 0 2024 0 -1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _592_
timestamp 1644511149
transform 1 0 2024 0 -1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_2  input1
timestamp 1644511149
transform 1 0 11868 0 -1 17408
box -38 -48 406 592
<< labels >>
rlabel metal2 s 11582 19200 11694 20000 6 active
port 0 nsew signal input
rlabel metal2 s 10938 0 11050 800 6 io_in[0]
port 1 nsew signal input
rlabel metal2 s 34122 19200 34234 20000 6 io_in[10]
port 2 nsew signal input
rlabel metal2 s 14158 19200 14270 20000 6 io_in[11]
port 3 nsew signal input
rlabel metal3 s 49200 14228 50000 14468 6 io_in[12]
port 4 nsew signal input
rlabel metal2 s 16734 0 16846 800 6 io_in[13]
port 5 nsew signal input
rlabel metal2 s 27682 19200 27794 20000 6 io_in[14]
port 6 nsew signal input
rlabel metal3 s 49200 15588 50000 15828 6 io_in[15]
port 7 nsew signal input
rlabel metal2 s 38630 0 38742 800 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 21886 19200 21998 20000 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 23174 19200 23286 20000 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 30258 0 30370 800 6 io_in[19]
port 11 nsew signal input
rlabel metal3 s 0 11508 800 11748 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s -10 19200 102 20000 6 io_in[20]
port 13 nsew signal input
rlabel metal3 s 0 13548 800 13788 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 46358 0 46470 800 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 21242 19200 21354 20000 6 io_in[23]
port 16 nsew signal input
rlabel metal2 s 19310 19200 19422 20000 6 io_in[24]
port 17 nsew signal input
rlabel metal2 s 26394 0 26506 800 6 io_in[25]
port 18 nsew signal input
rlabel metal2 s 25750 0 25862 800 6 io_in[26]
port 19 nsew signal input
rlabel metal2 s 43138 0 43250 800 6 io_in[27]
port 20 nsew signal input
rlabel metal2 s 23174 0 23286 800 6 io_in[28]
port 21 nsew signal input
rlabel metal2 s 49578 19200 49690 20000 6 io_in[29]
port 22 nsew signal input
rlabel metal2 s 11582 0 11694 800 6 io_in[2]
port 23 nsew signal input
rlabel metal2 s 48934 0 49046 800 6 io_in[30]
port 24 nsew signal input
rlabel metal2 s 10294 19200 10406 20000 6 io_in[31]
port 25 nsew signal input
rlabel metal2 s 21886 0 21998 800 6 io_in[32]
port 26 nsew signal input
rlabel metal3 s 0 18308 800 18548 6 io_in[33]
port 27 nsew signal input
rlabel metal2 s 41206 19200 41318 20000 6 io_in[34]
port 28 nsew signal input
rlabel metal2 s 45070 19200 45182 20000 6 io_in[35]
port 29 nsew signal input
rlabel metal3 s 49200 6748 50000 6988 6 io_in[36]
port 30 nsew signal input
rlabel metal2 s 45714 19200 45826 20000 6 io_in[37]
port 31 nsew signal input
rlabel metal2 s 34766 19200 34878 20000 6 io_in[3]
port 32 nsew signal input
rlabel metal3 s 49200 6068 50000 6308 6 io_in[4]
port 33 nsew signal input
rlabel metal3 s 49200 18308 50000 18548 6 io_in[5]
port 34 nsew signal input
rlabel metal2 s 1278 19200 1390 20000 6 io_in[6]
port 35 nsew signal input
rlabel metal3 s 0 14908 800 15148 6 io_in[7]
port 36 nsew signal input
rlabel metal3 s 49200 8108 50000 8348 6 io_in[8]
port 37 nsew signal input
rlabel metal2 s 20598 19200 20710 20000 6 io_in[9]
port 38 nsew signal input
rlabel metal2 s 18666 0 18778 800 6 io_oeb[0]
port 39 nsew signal tristate
rlabel metal3 s 0 12188 800 12428 6 io_oeb[10]
port 40 nsew signal tristate
rlabel metal3 s 49200 4708 50000 4948 6 io_oeb[11]
port 41 nsew signal tristate
rlabel metal2 s 45714 0 45826 800 6 io_oeb[12]
port 42 nsew signal tristate
rlabel metal2 s 45070 0 45182 800 6 io_oeb[13]
port 43 nsew signal tristate
rlabel metal3 s 0 3348 800 3588 6 io_oeb[14]
port 44 nsew signal tristate
rlabel metal2 s 24462 19200 24574 20000 6 io_oeb[15]
port 45 nsew signal tristate
rlabel metal2 s 37342 0 37454 800 6 io_oeb[16]
port 46 nsew signal tristate
rlabel metal2 s 9650 0 9762 800 6 io_oeb[17]
port 47 nsew signal tristate
rlabel metal2 s 39918 19200 40030 20000 6 io_oeb[18]
port 48 nsew signal tristate
rlabel metal2 s 25106 19200 25218 20000 6 io_oeb[19]
port 49 nsew signal tristate
rlabel metal2 s 27682 0 27794 800 6 io_oeb[1]
port 50 nsew signal tristate
rlabel metal3 s 49200 -52 50000 188 6 io_oeb[20]
port 51 nsew signal tristate
rlabel metal2 s 16090 19200 16202 20000 6 io_oeb[21]
port 52 nsew signal tristate
rlabel metal2 s 3854 0 3966 800 6 io_oeb[22]
port 53 nsew signal tristate
rlabel metal2 s 32190 19200 32302 20000 6 io_oeb[23]
port 54 nsew signal tristate
rlabel metal2 s 32834 19200 32946 20000 6 io_oeb[24]
port 55 nsew signal tristate
rlabel metal2 s 33478 0 33590 800 6 io_oeb[25]
port 56 nsew signal tristate
rlabel metal3 s 49200 12188 50000 12428 6 io_oeb[26]
port 57 nsew signal tristate
rlabel metal2 s 35410 19200 35522 20000 6 io_oeb[27]
port 58 nsew signal tristate
rlabel metal2 s 29614 0 29726 800 6 io_oeb[28]
port 59 nsew signal tristate
rlabel metal3 s 49200 7428 50000 7668 6 io_oeb[29]
port 60 nsew signal tristate
rlabel metal2 s 43782 19200 43894 20000 6 io_oeb[2]
port 61 nsew signal tristate
rlabel metal2 s 16734 19200 16846 20000 6 io_oeb[30]
port 62 nsew signal tristate
rlabel metal2 s 28970 0 29082 800 6 io_oeb[31]
port 63 nsew signal tristate
rlabel metal3 s 0 17628 800 17868 6 io_oeb[32]
port 64 nsew signal tristate
rlabel metal2 s 34766 0 34878 800 6 io_oeb[33]
port 65 nsew signal tristate
rlabel metal2 s 22530 19200 22642 20000 6 io_oeb[34]
port 66 nsew signal tristate
rlabel metal3 s 0 15588 800 15828 6 io_oeb[35]
port 67 nsew signal tristate
rlabel metal3 s 0 8108 800 8348 6 io_oeb[36]
port 68 nsew signal tristate
rlabel metal3 s 0 12868 800 13108 6 io_oeb[37]
port 69 nsew signal tristate
rlabel metal2 s 18022 0 18134 800 6 io_oeb[3]
port 70 nsew signal tristate
rlabel metal2 s 36054 0 36166 800 6 io_oeb[4]
port 71 nsew signal tristate
rlabel metal2 s 2566 19200 2678 20000 6 io_oeb[5]
port 72 nsew signal tristate
rlabel metal2 s 47646 0 47758 800 6 io_oeb[6]
port 73 nsew signal tristate
rlabel metal2 s 23818 19200 23930 20000 6 io_oeb[7]
port 74 nsew signal tristate
rlabel metal2 s 3210 0 3322 800 6 io_oeb[8]
port 75 nsew signal tristate
rlabel metal2 s 7718 0 7830 800 6 io_oeb[9]
port 76 nsew signal tristate
rlabel metal3 s 49200 17628 50000 17868 6 io_out[0]
port 77 nsew signal tristate
rlabel metal3 s 49200 4028 50000 4268 6 io_out[10]
port 78 nsew signal tristate
rlabel metal3 s 0 1988 800 2228 6 io_out[11]
port 79 nsew signal tristate
rlabel metal3 s 0 5388 800 5628 6 io_out[12]
port 80 nsew signal tristate
rlabel metal2 s 28326 0 28438 800 6 io_out[13]
port 81 nsew signal tristate
rlabel metal3 s 49200 12868 50000 13108 6 io_out[14]
port 82 nsew signal tristate
rlabel metal2 s 8362 19200 8474 20000 6 io_out[15]
port 83 nsew signal tristate
rlabel metal3 s 49200 3348 50000 3588 6 io_out[16]
port 84 nsew signal tristate
rlabel metal2 s 47002 19200 47114 20000 6 io_out[17]
port 85 nsew signal tristate
rlabel metal2 s 32834 0 32946 800 6 io_out[18]
port 86 nsew signal tristate
rlabel metal3 s 0 16948 800 17188 6 io_out[19]
port 87 nsew signal tristate
rlabel metal2 s 37986 19200 38098 20000 6 io_out[1]
port 88 nsew signal tristate
rlabel metal2 s 43138 19200 43250 20000 6 io_out[20]
port 89 nsew signal tristate
rlabel metal2 s 7718 19200 7830 20000 6 io_out[21]
port 90 nsew signal tristate
rlabel metal2 s 22530 0 22642 800 6 io_out[22]
port 91 nsew signal tristate
rlabel metal3 s 49200 628 50000 868 6 io_out[23]
port 92 nsew signal tristate
rlabel metal2 s 19310 0 19422 800 6 io_out[24]
port 93 nsew signal tristate
rlabel metal2 s 40562 19200 40674 20000 6 io_out[25]
port 94 nsew signal tristate
rlabel metal3 s 0 4028 800 4268 6 io_out[26]
port 95 nsew signal tristate
rlabel metal2 s 41850 19200 41962 20000 6 io_out[27]
port 96 nsew signal tristate
rlabel metal2 s 12226 0 12338 800 6 io_out[28]
port 97 nsew signal tristate
rlabel metal2 s 36698 0 36810 800 6 io_out[29]
port 98 nsew signal tristate
rlabel metal2 s 5142 0 5254 800 6 io_out[2]
port 99 nsew signal tristate
rlabel metal3 s 0 4708 800 4948 6 io_out[30]
port 100 nsew signal tristate
rlabel metal3 s 0 10148 800 10388 6 io_out[31]
port 101 nsew signal tristate
rlabel metal2 s 12226 19200 12338 20000 6 io_out[32]
port 102 nsew signal tristate
rlabel metal2 s 40562 0 40674 800 6 io_out[33]
port 103 nsew signal tristate
rlabel metal3 s 49200 13548 50000 13788 6 io_out[34]
port 104 nsew signal tristate
rlabel metal3 s 49200 11508 50000 11748 6 io_out[35]
port 105 nsew signal tristate
rlabel metal2 s 25750 19200 25862 20000 6 io_out[36]
port 106 nsew signal tristate
rlabel metal3 s 49200 16268 50000 16508 6 io_out[37]
port 107 nsew signal tristate
rlabel metal2 s 9650 19200 9762 20000 6 io_out[3]
port 108 nsew signal tristate
rlabel metal3 s 49200 5388 50000 5628 6 io_out[4]
port 109 nsew signal tristate
rlabel metal2 s 30902 19200 31014 20000 6 io_out[5]
port 110 nsew signal tristate
rlabel metal2 s 48290 19200 48402 20000 6 io_out[6]
port 111 nsew signal tristate
rlabel metal3 s 0 14228 800 14468 6 io_out[7]
port 112 nsew signal tristate
rlabel metal2 s 13514 0 13626 800 6 io_out[8]
port 113 nsew signal tristate
rlabel metal3 s 0 10828 800 11068 6 io_out[9]
port 114 nsew signal tristate
rlabel metal2 s 41206 0 41318 800 6 la1_data_in[0]
port 115 nsew signal input
rlabel metal2 s 15446 0 15558 800 6 la1_data_in[10]
port 116 nsew signal input
rlabel metal2 s 39918 0 40030 800 6 la1_data_in[11]
port 117 nsew signal input
rlabel metal2 s 5786 19200 5898 20000 6 la1_data_in[12]
port 118 nsew signal input
rlabel metal2 s 23818 0 23930 800 6 la1_data_in[13]
port 119 nsew signal input
rlabel metal3 s 0 9468 800 9708 6 la1_data_in[14]
port 120 nsew signal input
rlabel metal2 s 26394 19200 26506 20000 6 la1_data_in[15]
port 121 nsew signal input
rlabel metal2 s 36698 19200 36810 20000 6 la1_data_in[16]
port 122 nsew signal input
rlabel metal2 s 31546 19200 31658 20000 6 la1_data_in[17]
port 123 nsew signal input
rlabel metal2 s 30902 0 31014 800 6 la1_data_in[18]
port 124 nsew signal input
rlabel metal2 s 27038 19200 27150 20000 6 la1_data_in[19]
port 125 nsew signal input
rlabel metal2 s 14158 0 14270 800 6 la1_data_in[1]
port 126 nsew signal input
rlabel metal2 s 5142 19200 5254 20000 6 la1_data_in[20]
port 127 nsew signal input
rlabel metal2 s 48934 19200 49046 20000 6 la1_data_in[21]
port 128 nsew signal input
rlabel metal2 s 41850 0 41962 800 6 la1_data_in[22]
port 129 nsew signal input
rlabel metal3 s 0 628 800 868 6 la1_data_in[23]
port 130 nsew signal input
rlabel metal2 s 10294 0 10406 800 6 la1_data_in[24]
port 131 nsew signal input
rlabel metal2 s 6430 19200 6542 20000 6 la1_data_in[25]
port 132 nsew signal input
rlabel metal2 s 37986 0 38098 800 6 la1_data_in[26]
port 133 nsew signal input
rlabel metal2 s 20598 0 20710 800 6 la1_data_in[27]
port 134 nsew signal input
rlabel metal2 s 3210 19200 3322 20000 6 la1_data_in[28]
port 135 nsew signal input
rlabel metal2 s 14802 19200 14914 20000 6 la1_data_in[29]
port 136 nsew signal input
rlabel metal2 s 8362 0 8474 800 6 la1_data_in[2]
port 137 nsew signal input
rlabel metal2 s 1278 0 1390 800 6 la1_data_in[30]
port 138 nsew signal input
rlabel metal2 s 27038 0 27150 800 6 la1_data_in[31]
port 139 nsew signal input
rlabel metal2 s 1922 19200 2034 20000 6 la1_data_in[3]
port 140 nsew signal input
rlabel metal2 s 44426 19200 44538 20000 6 la1_data_in[4]
port 141 nsew signal input
rlabel metal3 s 49200 1988 50000 2228 6 la1_data_in[5]
port 142 nsew signal input
rlabel metal2 s 28326 19200 28438 20000 6 la1_data_in[6]
port 143 nsew signal input
rlabel metal3 s 0 16268 800 16508 6 la1_data_in[7]
port 144 nsew signal input
rlabel metal2 s 28970 19200 29082 20000 6 la1_data_in[8]
port 145 nsew signal input
rlabel metal2 s 3854 19200 3966 20000 6 la1_data_in[9]
port 146 nsew signal input
rlabel metal2 s 5786 0 5898 800 6 la1_data_out[0]
port 147 nsew signal tristate
rlabel metal2 s 43782 0 43894 800 6 la1_data_out[10]
port 148 nsew signal tristate
rlabel metal2 s 16090 0 16202 800 6 la1_data_out[11]
port 149 nsew signal tristate
rlabel metal3 s 49200 16948 50000 17188 6 la1_data_out[12]
port 150 nsew signal tristate
rlabel metal2 s 18022 19200 18134 20000 6 la1_data_out[13]
port 151 nsew signal tristate
rlabel metal2 s 33478 19200 33590 20000 6 la1_data_out[14]
port 152 nsew signal tristate
rlabel metal3 s 0 1308 800 1548 6 la1_data_out[15]
port 153 nsew signal tristate
rlabel metal2 s 47002 0 47114 800 6 la1_data_out[16]
port 154 nsew signal tristate
rlabel metal3 s 49200 10148 50000 10388 6 la1_data_out[17]
port 155 nsew signal tristate
rlabel metal2 s 18666 19200 18778 20000 6 la1_data_out[18]
port 156 nsew signal tristate
rlabel metal3 s 49200 2668 50000 2908 6 la1_data_out[19]
port 157 nsew signal tristate
rlabel metal2 s 10938 19200 11050 20000 6 la1_data_out[1]
port 158 nsew signal tristate
rlabel metal3 s 0 7428 800 7668 6 la1_data_out[20]
port 159 nsew signal tristate
rlabel metal3 s 49200 14908 50000 15148 6 la1_data_out[21]
port 160 nsew signal tristate
rlabel metal2 s 36054 19200 36166 20000 6 la1_data_out[22]
port 161 nsew signal tristate
rlabel metal2 s 9006 0 9118 800 6 la1_data_out[23]
port 162 nsew signal tristate
rlabel metal2 s 48290 0 48402 800 6 la1_data_out[24]
port 163 nsew signal tristate
rlabel metal3 s 0 2668 800 2908 6 la1_data_out[25]
port 164 nsew signal tristate
rlabel metal2 s 39274 0 39386 800 6 la1_data_out[26]
port 165 nsew signal tristate
rlabel metal2 s 12870 19200 12982 20000 6 la1_data_out[27]
port 166 nsew signal tristate
rlabel metal2 s 31546 0 31658 800 6 la1_data_out[28]
port 167 nsew signal tristate
rlabel metal2 s 4498 0 4610 800 6 la1_data_out[29]
port 168 nsew signal tristate
rlabel metal2 s 14802 0 14914 800 6 la1_data_out[2]
port 169 nsew signal tristate
rlabel metal2 s 44426 0 44538 800 6 la1_data_out[30]
port 170 nsew signal tristate
rlabel metal3 s 49200 18988 50000 19228 6 la1_data_out[31]
port 171 nsew signal tristate
rlabel metal3 s 0 6748 800 6988 6 la1_data_out[3]
port 172 nsew signal tristate
rlabel metal2 s 32190 0 32302 800 6 la1_data_out[4]
port 173 nsew signal tristate
rlabel metal2 s 2566 0 2678 800 6 la1_data_out[5]
port 174 nsew signal tristate
rlabel metal2 s 49578 0 49690 800 6 la1_data_out[6]
port 175 nsew signal tristate
rlabel metal2 s 634 0 746 800 6 la1_data_out[7]
port 176 nsew signal tristate
rlabel metal3 s 49200 10828 50000 11068 6 la1_data_out[8]
port 177 nsew signal tristate
rlabel metal2 s 47646 19200 47758 20000 6 la1_data_out[9]
port 178 nsew signal tristate
rlabel metal2 s 35410 0 35522 800 6 la1_oenb[0]
port 179 nsew signal input
rlabel metal2 s 46358 19200 46470 20000 6 la1_oenb[10]
port 180 nsew signal input
rlabel metal3 s 0 19668 800 19908 6 la1_oenb[11]
port 181 nsew signal input
rlabel metal2 s 634 19200 746 20000 6 la1_oenb[12]
port 182 nsew signal input
rlabel metal2 s 21242 0 21354 800 6 la1_oenb[13]
port 183 nsew signal input
rlabel metal2 s -10 0 102 800 6 la1_oenb[14]
port 184 nsew signal input
rlabel metal2 s 25106 0 25218 800 6 la1_oenb[15]
port 185 nsew signal input
rlabel metal2 s 4498 19200 4610 20000 6 la1_oenb[16]
port 186 nsew signal input
rlabel metal2 s 17378 19200 17490 20000 6 la1_oenb[17]
port 187 nsew signal input
rlabel metal2 s 30258 19200 30370 20000 6 la1_oenb[18]
port 188 nsew signal input
rlabel metal3 s 0 18988 800 19228 6 la1_oenb[19]
port 189 nsew signal input
rlabel metal2 s 6430 0 6542 800 6 la1_oenb[1]
port 190 nsew signal input
rlabel metal2 s 1922 0 2034 800 6 la1_oenb[20]
port 191 nsew signal input
rlabel metal2 s 37342 19200 37454 20000 6 la1_oenb[21]
port 192 nsew signal input
rlabel metal2 s 29614 19200 29726 20000 6 la1_oenb[22]
port 193 nsew signal input
rlabel metal2 s 17378 0 17490 800 6 la1_oenb[23]
port 194 nsew signal input
rlabel metal2 s 42494 19200 42606 20000 6 la1_oenb[24]
port 195 nsew signal input
rlabel metal2 s 42494 0 42606 800 6 la1_oenb[25]
port 196 nsew signal input
rlabel metal2 s 7074 19200 7186 20000 6 la1_oenb[26]
port 197 nsew signal input
rlabel metal3 s 49200 9468 50000 9708 6 la1_oenb[27]
port 198 nsew signal input
rlabel metal2 s 7074 0 7186 800 6 la1_oenb[28]
port 199 nsew signal input
rlabel metal2 s 12870 0 12982 800 6 la1_oenb[29]
port 200 nsew signal input
rlabel metal3 s 0 6068 800 6308 6 la1_oenb[2]
port 201 nsew signal input
rlabel metal3 s 49200 8788 50000 9028 6 la1_oenb[30]
port 202 nsew signal input
rlabel metal2 s 19954 0 20066 800 6 la1_oenb[31]
port 203 nsew signal input
rlabel metal2 s 39274 19200 39386 20000 6 la1_oenb[3]
port 204 nsew signal input
rlabel metal2 s 38630 19200 38742 20000 6 la1_oenb[4]
port 205 nsew signal input
rlabel metal2 s 13514 19200 13626 20000 6 la1_oenb[5]
port 206 nsew signal input
rlabel metal2 s 19954 19200 20066 20000 6 la1_oenb[6]
port 207 nsew signal input
rlabel metal2 s 24462 0 24574 800 6 la1_oenb[7]
port 208 nsew signal input
rlabel metal3 s 0 8788 800 9028 6 la1_oenb[8]
port 209 nsew signal input
rlabel metal2 s 9006 19200 9118 20000 6 la1_oenb[9]
port 210 nsew signal input
rlabel metal4 s 8910 2128 9230 17456 6 vccd1
port 211 nsew power input
rlabel metal4 s 24840 2128 25160 17456 6 vccd1
port 211 nsew power input
rlabel metal4 s 40771 2128 41091 17456 6 vccd1
port 211 nsew power input
rlabel metal4 s 16874 2128 17194 17456 6 vssd1
port 212 nsew ground input
rlabel metal4 s 32805 2128 33125 17456 6 vssd1
port 212 nsew ground input
rlabel metal3 s 49200 1308 50000 1548 6 wb_clk_i
port 213 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 50000 20000
<< end >>
