magic
tech sky130A
magscale 1 2
timestamp 1671183550
<< obsli1 >>
rect 1104 2159 28888 47345
<< obsm1 >>
rect 14 2048 29978 47456
<< metal2 >>
rect -10 49200 102 49800
rect 634 49200 746 49800
rect 1278 49200 1390 49800
rect 1922 49200 2034 49800
rect 2566 49200 2678 49800
rect 3210 49200 3322 49800
rect 4498 49200 4610 49800
rect 5142 49200 5254 49800
rect 5786 49200 5898 49800
rect 6430 49200 6542 49800
rect 7074 49200 7186 49800
rect 7718 49200 7830 49800
rect 8362 49200 8474 49800
rect 9650 49200 9762 49800
rect 10294 49200 10406 49800
rect 10938 49200 11050 49800
rect 11582 49200 11694 49800
rect 12226 49200 12338 49800
rect 12870 49200 12982 49800
rect 13514 49200 13626 49800
rect 14802 49200 14914 49800
rect 15446 49200 15558 49800
rect 16090 49200 16202 49800
rect 16734 49200 16846 49800
rect 17378 49200 17490 49800
rect 18022 49200 18134 49800
rect 18666 49200 18778 49800
rect 19954 49200 20066 49800
rect 20598 49200 20710 49800
rect 21242 49200 21354 49800
rect 21886 49200 21998 49800
rect 22530 49200 22642 49800
rect 23174 49200 23286 49800
rect 23818 49200 23930 49800
rect 25106 49200 25218 49800
rect 25750 49200 25862 49800
rect 26394 49200 26506 49800
rect 27038 49200 27150 49800
rect 27682 49200 27794 49800
rect 28326 49200 28438 49800
rect 28970 49200 29082 49800
rect 29614 49200 29726 49800
rect -10 200 102 800
rect 634 200 746 800
rect 1278 200 1390 800
rect 1922 200 2034 800
rect 2566 200 2678 800
rect 3210 200 3322 800
rect 3854 200 3966 800
rect 4498 200 4610 800
rect 5786 200 5898 800
rect 6430 200 6542 800
rect 7074 200 7186 800
rect 7718 200 7830 800
rect 8362 200 8474 800
rect 9006 200 9118 800
rect 9650 200 9762 800
rect 10938 200 11050 800
rect 11582 200 11694 800
rect 12226 200 12338 800
rect 12870 200 12982 800
rect 13514 200 13626 800
rect 14158 200 14270 800
rect 14802 200 14914 800
rect 16090 200 16202 800
rect 16734 200 16846 800
rect 17378 200 17490 800
rect 18022 200 18134 800
rect 18666 200 18778 800
rect 19310 200 19422 800
rect 19954 200 20066 800
rect 21242 200 21354 800
rect 21886 200 21998 800
rect 22530 200 22642 800
rect 23174 200 23286 800
rect 23818 200 23930 800
rect 24462 200 24574 800
rect 25106 200 25218 800
rect 26394 200 26506 800
rect 27038 200 27150 800
rect 27682 200 27794 800
rect 28326 200 28438 800
rect 28970 200 29082 800
rect 29614 200 29726 800
<< obsm2 >>
rect 158 49144 578 49745
rect 802 49144 1222 49745
rect 1446 49144 1866 49745
rect 2090 49144 2510 49745
rect 2734 49144 3154 49745
rect 3378 49144 4442 49745
rect 4666 49144 5086 49745
rect 5310 49144 5730 49745
rect 5954 49144 6374 49745
rect 6598 49144 7018 49745
rect 7242 49144 7662 49745
rect 7886 49144 8306 49745
rect 8530 49144 9594 49745
rect 9818 49144 10238 49745
rect 10462 49144 10882 49745
rect 11106 49144 11526 49745
rect 11750 49144 12170 49745
rect 12394 49144 12814 49745
rect 13038 49144 13458 49745
rect 13682 49144 14746 49745
rect 14970 49144 15390 49745
rect 15614 49144 16034 49745
rect 16258 49144 16678 49745
rect 16902 49144 17322 49745
rect 17546 49144 17966 49745
rect 18190 49144 18610 49745
rect 18834 49144 19898 49745
rect 20122 49144 20542 49745
rect 20766 49144 21186 49745
rect 21410 49144 21830 49745
rect 22054 49144 22474 49745
rect 22698 49144 23118 49745
rect 23342 49144 23762 49745
rect 23986 49144 25050 49745
rect 25274 49144 25694 49745
rect 25918 49144 26338 49745
rect 26562 49144 26982 49745
rect 27206 49144 27626 49745
rect 27850 49144 28270 49745
rect 28494 49144 28914 49745
rect 29138 49144 29558 49745
rect 29782 49144 29974 49745
rect 20 856 29974 49144
rect 158 800 578 856
rect 802 800 1222 856
rect 1446 800 1866 856
rect 2090 800 2510 856
rect 2734 800 3154 856
rect 3378 800 3798 856
rect 4022 800 4442 856
rect 4666 800 5730 856
rect 5954 800 6374 856
rect 6598 800 7018 856
rect 7242 800 7662 856
rect 7886 800 8306 856
rect 8530 800 8950 856
rect 9174 800 9594 856
rect 9818 800 10882 856
rect 11106 800 11526 856
rect 11750 800 12170 856
rect 12394 800 12814 856
rect 13038 800 13458 856
rect 13682 800 14102 856
rect 14326 800 14746 856
rect 14970 800 16034 856
rect 16258 800 16678 856
rect 16902 800 17322 856
rect 17546 800 17966 856
rect 18190 800 18610 856
rect 18834 800 19254 856
rect 19478 800 19898 856
rect 20122 800 21186 856
rect 21410 800 21830 856
rect 22054 800 22474 856
rect 22698 800 23118 856
rect 23342 800 23762 856
rect 23986 800 24406 856
rect 24630 800 25050 856
rect 25274 800 26338 856
rect 26562 800 26982 856
rect 27206 800 27626 856
rect 27850 800 28270 856
rect 28494 800 28914 856
rect 29138 800 29558 856
rect 29782 800 29974 856
<< metal3 >>
rect 200 49588 800 49828
rect 29200 48908 29800 49148
rect 200 48228 800 48468
rect 29200 48228 29800 48468
rect 200 47548 800 47788
rect 29200 47548 29800 47788
rect 200 46868 800 47108
rect 29200 46868 29800 47108
rect 200 46188 800 46428
rect 29200 46188 29800 46428
rect 200 45508 800 45748
rect 29200 45508 29800 45748
rect 200 44828 800 45068
rect 29200 44828 29800 45068
rect 200 44148 800 44388
rect 29200 43468 29800 43708
rect 200 42788 800 43028
rect 29200 42788 29800 43028
rect 200 42108 800 42348
rect 29200 42108 29800 42348
rect 200 41428 800 41668
rect 29200 41428 29800 41668
rect 200 40748 800 40988
rect 29200 40748 29800 40988
rect 200 40068 800 40308
rect 29200 40068 29800 40308
rect 200 39388 800 39628
rect 29200 39388 29800 39628
rect 200 38708 800 38948
rect 29200 38028 29800 38268
rect 200 37348 800 37588
rect 29200 37348 29800 37588
rect 200 36668 800 36908
rect 29200 36668 29800 36908
rect 200 35988 800 36228
rect 29200 35988 29800 36228
rect 200 35308 800 35548
rect 29200 35308 29800 35548
rect 200 34628 800 34868
rect 29200 34628 29800 34868
rect 200 33948 800 34188
rect 29200 33948 29800 34188
rect 200 33268 800 33508
rect 29200 32588 29800 32828
rect 200 31908 800 32148
rect 29200 31908 29800 32148
rect 200 31228 800 31468
rect 29200 31228 29800 31468
rect 200 30548 800 30788
rect 29200 30548 29800 30788
rect 200 29868 800 30108
rect 29200 29868 29800 30108
rect 200 29188 800 29428
rect 29200 29188 29800 29428
rect 200 28508 800 28748
rect 29200 28508 29800 28748
rect 200 27828 800 28068
rect 29200 27148 29800 27388
rect 200 26468 800 26708
rect 29200 26468 29800 26708
rect 200 25788 800 26028
rect 29200 25788 29800 26028
rect 200 25108 800 25348
rect 29200 25108 29800 25348
rect 200 24428 800 24668
rect 29200 24428 29800 24668
rect 200 23748 800 23988
rect 29200 23748 29800 23988
rect 200 23068 800 23308
rect 29200 23068 29800 23308
rect 200 22388 800 22628
rect 29200 21708 29800 21948
rect 200 21028 800 21268
rect 29200 21028 29800 21268
rect 200 20348 800 20588
rect 29200 20348 29800 20588
rect 200 19668 800 19908
rect 29200 19668 29800 19908
rect 200 18988 800 19228
rect 29200 18988 29800 19228
rect 200 18308 800 18548
rect 29200 18308 29800 18548
rect 200 17628 800 17868
rect 29200 17628 29800 17868
rect 200 16948 800 17188
rect 29200 16268 29800 16508
rect 200 15588 800 15828
rect 29200 15588 29800 15828
rect 200 14908 800 15148
rect 29200 14908 29800 15148
rect 200 14228 800 14468
rect 29200 14228 29800 14468
rect 200 13548 800 13788
rect 29200 13548 29800 13788
rect 200 12868 800 13108
rect 29200 12868 29800 13108
rect 200 12188 800 12428
rect 29200 12188 29800 12428
rect 200 11508 800 11748
rect 29200 10828 29800 11068
rect 200 10148 800 10388
rect 29200 10148 29800 10388
rect 200 9468 800 9708
rect 29200 9468 29800 9708
rect 200 8788 800 9028
rect 29200 8788 29800 9028
rect 200 8108 800 8348
rect 29200 8108 29800 8348
rect 200 7428 800 7668
rect 29200 7428 29800 7668
rect 200 6748 800 6988
rect 29200 6748 29800 6988
rect 200 6068 800 6308
rect 29200 5388 29800 5628
rect 200 4708 800 4948
rect 29200 4708 29800 4948
rect 200 4028 800 4268
rect 29200 4028 29800 4268
rect 200 3348 800 3588
rect 29200 3348 29800 3588
rect 200 2668 800 2908
rect 29200 2668 29800 2908
rect 200 1988 800 2228
rect 29200 1988 29800 2228
rect 200 1308 800 1548
rect 29200 1308 29800 1548
rect 200 628 800 868
rect 29200 -52 29800 188
<< obsm3 >>
rect 880 49508 29979 49741
rect 800 49228 29979 49508
rect 800 48828 29120 49228
rect 29880 48828 29979 49228
rect 800 48548 29979 48828
rect 880 48148 29120 48548
rect 29880 48148 29979 48548
rect 800 47868 29979 48148
rect 880 47468 29120 47868
rect 29880 47468 29979 47868
rect 800 47188 29979 47468
rect 880 46788 29120 47188
rect 29880 46788 29979 47188
rect 800 46508 29979 46788
rect 880 46108 29120 46508
rect 29880 46108 29979 46508
rect 800 45828 29979 46108
rect 880 45428 29120 45828
rect 29880 45428 29979 45828
rect 800 45148 29979 45428
rect 880 44748 29120 45148
rect 29880 44748 29979 45148
rect 800 44468 29979 44748
rect 880 44068 29979 44468
rect 800 43788 29979 44068
rect 800 43388 29120 43788
rect 29880 43388 29979 43788
rect 800 43108 29979 43388
rect 880 42708 29120 43108
rect 29880 42708 29979 43108
rect 800 42428 29979 42708
rect 880 42028 29120 42428
rect 29880 42028 29979 42428
rect 800 41748 29979 42028
rect 880 41348 29120 41748
rect 29880 41348 29979 41748
rect 800 41068 29979 41348
rect 880 40668 29120 41068
rect 29880 40668 29979 41068
rect 800 40388 29979 40668
rect 880 39988 29120 40388
rect 29880 39988 29979 40388
rect 800 39708 29979 39988
rect 880 39308 29120 39708
rect 29880 39308 29979 39708
rect 800 39028 29979 39308
rect 880 38628 29979 39028
rect 800 38348 29979 38628
rect 800 37948 29120 38348
rect 29880 37948 29979 38348
rect 800 37668 29979 37948
rect 880 37268 29120 37668
rect 29880 37268 29979 37668
rect 800 36988 29979 37268
rect 880 36588 29120 36988
rect 29880 36588 29979 36988
rect 800 36308 29979 36588
rect 880 35908 29120 36308
rect 29880 35908 29979 36308
rect 800 35628 29979 35908
rect 880 35228 29120 35628
rect 29880 35228 29979 35628
rect 800 34948 29979 35228
rect 880 34548 29120 34948
rect 29880 34548 29979 34948
rect 800 34268 29979 34548
rect 880 33868 29120 34268
rect 29880 33868 29979 34268
rect 800 33588 29979 33868
rect 880 33188 29979 33588
rect 800 32908 29979 33188
rect 800 32508 29120 32908
rect 29880 32508 29979 32908
rect 800 32228 29979 32508
rect 880 31828 29120 32228
rect 29880 31828 29979 32228
rect 800 31548 29979 31828
rect 880 31148 29120 31548
rect 29880 31148 29979 31548
rect 800 30868 29979 31148
rect 880 30468 29120 30868
rect 29880 30468 29979 30868
rect 800 30188 29979 30468
rect 880 29788 29120 30188
rect 29880 29788 29979 30188
rect 800 29508 29979 29788
rect 880 29108 29120 29508
rect 29880 29108 29979 29508
rect 800 28828 29979 29108
rect 880 28428 29120 28828
rect 29880 28428 29979 28828
rect 800 28148 29979 28428
rect 880 27748 29979 28148
rect 800 27468 29979 27748
rect 800 27068 29120 27468
rect 29880 27068 29979 27468
rect 800 26788 29979 27068
rect 880 26388 29120 26788
rect 29880 26388 29979 26788
rect 800 26108 29979 26388
rect 880 25708 29120 26108
rect 29880 25708 29979 26108
rect 800 25428 29979 25708
rect 880 25028 29120 25428
rect 29880 25028 29979 25428
rect 800 24748 29979 25028
rect 880 24348 29120 24748
rect 29880 24348 29979 24748
rect 800 24068 29979 24348
rect 880 23668 29120 24068
rect 29880 23668 29979 24068
rect 800 23388 29979 23668
rect 880 22988 29120 23388
rect 29880 22988 29979 23388
rect 800 22708 29979 22988
rect 880 22308 29979 22708
rect 800 22028 29979 22308
rect 800 21628 29120 22028
rect 29880 21628 29979 22028
rect 800 21348 29979 21628
rect 880 20948 29120 21348
rect 29880 20948 29979 21348
rect 800 20668 29979 20948
rect 880 20268 29120 20668
rect 29880 20268 29979 20668
rect 800 19988 29979 20268
rect 880 19588 29120 19988
rect 29880 19588 29979 19988
rect 800 19308 29979 19588
rect 880 18908 29120 19308
rect 29880 18908 29979 19308
rect 800 18628 29979 18908
rect 880 18228 29120 18628
rect 29880 18228 29979 18628
rect 800 17948 29979 18228
rect 880 17548 29120 17948
rect 29880 17548 29979 17948
rect 800 17268 29979 17548
rect 880 16868 29979 17268
rect 800 16588 29979 16868
rect 800 16188 29120 16588
rect 29880 16188 29979 16588
rect 800 15908 29979 16188
rect 880 15508 29120 15908
rect 29880 15508 29979 15908
rect 800 15228 29979 15508
rect 880 14828 29120 15228
rect 29880 14828 29979 15228
rect 800 14548 29979 14828
rect 880 14148 29120 14548
rect 29880 14148 29979 14548
rect 800 13868 29979 14148
rect 880 13468 29120 13868
rect 29880 13468 29979 13868
rect 800 13188 29979 13468
rect 880 12788 29120 13188
rect 29880 12788 29979 13188
rect 800 12508 29979 12788
rect 880 12108 29120 12508
rect 29880 12108 29979 12508
rect 800 11828 29979 12108
rect 880 11428 29979 11828
rect 800 11148 29979 11428
rect 800 10748 29120 11148
rect 29880 10748 29979 11148
rect 800 10468 29979 10748
rect 880 10068 29120 10468
rect 29880 10068 29979 10468
rect 800 9788 29979 10068
rect 880 9388 29120 9788
rect 29880 9388 29979 9788
rect 800 9108 29979 9388
rect 880 8708 29120 9108
rect 29880 8708 29979 9108
rect 800 8428 29979 8708
rect 880 8028 29120 8428
rect 29880 8028 29979 8428
rect 800 7748 29979 8028
rect 880 7348 29120 7748
rect 29880 7348 29979 7748
rect 800 7068 29979 7348
rect 880 6668 29120 7068
rect 29880 6668 29979 7068
rect 800 6388 29979 6668
rect 880 5988 29979 6388
rect 800 5708 29979 5988
rect 800 5308 29120 5708
rect 29880 5308 29979 5708
rect 800 5028 29979 5308
rect 880 4628 29120 5028
rect 29880 4628 29979 5028
rect 800 4348 29979 4628
rect 880 3948 29120 4348
rect 29880 3948 29979 4348
rect 800 3668 29979 3948
rect 880 3268 29120 3668
rect 29880 3268 29979 3668
rect 800 2988 29979 3268
rect 880 2588 29120 2988
rect 29880 2588 29979 2988
rect 800 2308 29979 2588
rect 880 1908 29120 2308
rect 29880 1908 29979 2308
rect 800 1628 29979 1908
rect 880 1395 29120 1628
rect 29880 1395 29979 1628
<< metal4 >>
rect 4417 2128 4737 47376
rect 7890 2128 8210 47376
rect 11363 2128 11683 47376
rect 14836 2128 15156 47376
rect 18309 2128 18629 47376
rect 21782 2128 22102 47376
rect 25255 2128 25575 47376
rect 28728 2128 29048 47376
<< obsm4 >>
rect 18827 11867 18893 27981
<< labels >>
rlabel metal3 s 200 36668 800 36908 6 active
port 1 nsew signal input
rlabel metal2 s 12226 200 12338 800 6 io_in[0]
port 2 nsew signal input
rlabel metal2 s 12226 49200 12338 49800 6 io_in[10]
port 3 nsew signal input
rlabel metal3 s 200 40068 800 40308 6 io_in[11]
port 4 nsew signal input
rlabel metal3 s 29200 43468 29800 43708 6 io_in[12]
port 5 nsew signal input
rlabel metal2 s 18666 200 18778 800 6 io_in[13]
port 6 nsew signal input
rlabel metal2 s 5142 49200 5254 49800 6 io_in[14]
port 7 nsew signal input
rlabel metal3 s 29200 45508 29800 45748 6 io_in[15]
port 8 nsew signal input
rlabel metal3 s 29200 13548 29800 13788 6 io_in[16]
port 9 nsew signal input
rlabel metal3 s 200 48228 800 48468 6 io_in[17]
port 10 nsew signal input
rlabel metal2 s -10 49200 102 49800 6 io_in[18]
port 11 nsew signal input
rlabel metal3 s 29200 4028 29800 4268 6 io_in[19]
port 12 nsew signal input
rlabel metal3 s 200 12868 800 13108 6 io_in[1]
port 13 nsew signal input
rlabel metal3 s 200 23068 800 23308 6 io_in[20]
port 14 nsew signal input
rlabel metal3 s 200 14908 800 15148 6 io_in[21]
port 15 nsew signal input
rlabel metal3 s 29200 23068 29800 23308 6 io_in[22]
port 16 nsew signal input
rlabel metal3 s 200 47548 800 47788 6 io_in[23]
port 17 nsew signal input
rlabel metal3 s 200 45508 800 45748 6 io_in[24]
port 18 nsew signal input
rlabel metal2 s 29614 200 29726 800 6 io_in[25]
port 19 nsew signal input
rlabel metal2 s 28970 200 29082 800 6 io_in[26]
port 20 nsew signal input
rlabel metal3 s 29200 18988 29800 19228 6 io_in[27]
port 21 nsew signal input
rlabel metal2 s 26394 200 26506 800 6 io_in[28]
port 22 nsew signal input
rlabel metal2 s 29614 49200 29726 49800 6 io_in[29]
port 23 nsew signal input
rlabel metal2 s 12870 200 12982 800 6 io_in[2]
port 24 nsew signal input
rlabel metal3 s 29200 25788 29800 26028 6 io_in[30]
port 25 nsew signal input
rlabel metal3 s 200 35308 800 35548 6 io_in[31]
port 26 nsew signal input
rlabel metal2 s 24462 200 24574 800 6 io_in[32]
port 27 nsew signal input
rlabel metal3 s 200 20348 800 20588 6 io_in[33]
port 28 nsew signal input
rlabel metal2 s 20598 49200 20710 49800 6 io_in[34]
port 29 nsew signal input
rlabel metal2 s 25106 49200 25218 49800 6 io_in[35]
port 30 nsew signal input
rlabel metal3 s 29200 35308 29800 35548 6 io_in[36]
port 31 nsew signal input
rlabel metal2 s 25750 49200 25862 49800 6 io_in[37]
port 32 nsew signal input
rlabel metal2 s 12870 49200 12982 49800 6 io_in[3]
port 33 nsew signal input
rlabel metal3 s 29200 34628 29800 34868 6 io_in[4]
port 34 nsew signal input
rlabel metal3 s 29200 48228 29800 48468 6 io_in[5]
port 35 nsew signal input
rlabel metal3 s 200 24428 800 24668 6 io_in[6]
port 36 nsew signal input
rlabel metal3 s 200 16948 800 17188 6 io_in[7]
port 37 nsew signal input
rlabel metal3 s 29200 36668 29800 36908 6 io_in[8]
port 38 nsew signal input
rlabel metal3 s 200 46868 800 47108 6 io_in[9]
port 39 nsew signal input
rlabel metal2 s 21242 200 21354 800 6 io_oeb[0]
port 40 nsew signal output
rlabel metal3 s 200 13548 800 13788 6 io_oeb[10]
port 41 nsew signal output
rlabel metal3 s 29200 32588 29800 32828 6 io_oeb[11]
port 42 nsew signal output
rlabel metal3 s 29200 21708 29800 21948 6 io_oeb[12]
port 43 nsew signal output
rlabel metal3 s 29200 21028 29800 21268 6 io_oeb[13]
port 44 nsew signal output
rlabel metal3 s 200 3348 800 3588 6 io_oeb[14]
port 45 nsew signal output
rlabel metal2 s 1278 49200 1390 49800 6 io_oeb[15]
port 46 nsew signal output
rlabel metal3 s 29200 12188 29800 12428 6 io_oeb[16]
port 47 nsew signal output
rlabel metal2 s 10938 200 11050 800 6 io_oeb[17]
port 48 nsew signal output
rlabel metal2 s 18666 49200 18778 49800 6 io_oeb[18]
port 49 nsew signal output
rlabel metal2 s 1922 49200 2034 49800 6 io_oeb[19]
port 50 nsew signal output
rlabel metal3 s 29200 1308 29800 1548 6 io_oeb[1]
port 51 nsew signal output
rlabel metal3 s 29200 27148 29800 27388 6 io_oeb[20]
port 52 nsew signal output
rlabel metal3 s 200 41428 800 41668 6 io_oeb[21]
port 53 nsew signal output
rlabel metal2 s 3854 200 3966 800 6 io_oeb[22]
port 54 nsew signal output
rlabel metal2 s 10294 49200 10406 49800 6 io_oeb[23]
port 55 nsew signal output
rlabel metal2 s 10938 49200 11050 49800 6 io_oeb[24]
port 56 nsew signal output
rlabel metal3 s 29200 8108 29800 8348 6 io_oeb[25]
port 57 nsew signal output
rlabel metal3 s 29200 41428 29800 41668 6 io_oeb[26]
port 58 nsew signal output
rlabel metal2 s 13514 49200 13626 49800 6 io_oeb[27]
port 59 nsew signal output
rlabel metal3 s 29200 3348 29800 3588 6 io_oeb[28]
port 60 nsew signal output
rlabel metal3 s 29200 35988 29800 36228 6 io_oeb[29]
port 61 nsew signal output
rlabel metal2 s 23174 49200 23286 49800 6 io_oeb[2]
port 62 nsew signal output
rlabel metal3 s 200 42108 800 42348 6 io_oeb[30]
port 63 nsew signal output
rlabel metal3 s 29200 2668 29800 2908 6 io_oeb[31]
port 64 nsew signal output
rlabel metal3 s 200 19668 800 19908 6 io_oeb[32]
port 65 nsew signal output
rlabel metal3 s 29200 8788 29800 9028 6 io_oeb[33]
port 66 nsew signal output
rlabel metal3 s 200 49588 800 49828 6 io_oeb[34]
port 67 nsew signal output
rlabel metal3 s 200 17628 800 17868 6 io_oeb[35]
port 68 nsew signal output
rlabel metal3 s 200 8788 800 9028 6 io_oeb[36]
port 69 nsew signal output
rlabel metal3 s 200 14228 800 14468 6 io_oeb[37]
port 70 nsew signal output
rlabel metal2 s 19954 200 20066 800 6 io_oeb[3]
port 71 nsew signal output
rlabel metal3 s 29200 10148 29800 10388 6 io_oeb[4]
port 72 nsew signal output
rlabel metal3 s 200 25788 800 26028 6 io_oeb[5]
port 73 nsew signal output
rlabel metal3 s 29200 24428 29800 24668 6 io_oeb[6]
port 74 nsew signal output
rlabel metal2 s 634 49200 746 49800 6 io_oeb[7]
port 75 nsew signal output
rlabel metal2 s 3210 200 3322 800 6 io_oeb[8]
port 76 nsew signal output
rlabel metal2 s 8362 200 8474 800 6 io_oeb[9]
port 77 nsew signal output
rlabel metal3 s 29200 47548 29800 47788 6 io_out[0]
port 78 nsew signal output
rlabel metal3 s 29200 31908 29800 32148 6 io_out[10]
port 79 nsew signal output
rlabel metal3 s 200 1988 800 2228 6 io_out[11]
port 80 nsew signal output
rlabel metal3 s 200 6068 800 6308 6 io_out[12]
port 81 nsew signal output
rlabel metal3 s 29200 1988 29800 2228 6 io_out[13]
port 82 nsew signal output
rlabel metal3 s 29200 42108 29800 42348 6 io_out[14]
port 83 nsew signal output
rlabel metal3 s 200 33268 800 33508 6 io_out[15]
port 84 nsew signal output
rlabel metal3 s 29200 31228 29800 31468 6 io_out[16]
port 85 nsew signal output
rlabel metal2 s 27038 49200 27150 49800 6 io_out[17]
port 86 nsew signal output
rlabel metal3 s 29200 7428 29800 7668 6 io_out[18]
port 87 nsew signal output
rlabel metal3 s 200 18988 800 19228 6 io_out[19]
port 88 nsew signal output
rlabel metal2 s 16734 49200 16846 49800 6 io_out[1]
port 89 nsew signal output
rlabel metal2 s 22530 49200 22642 49800 6 io_out[20]
port 90 nsew signal output
rlabel metal3 s 200 31908 800 32148 6 io_out[21]
port 91 nsew signal output
rlabel metal2 s 25106 200 25218 800 6 io_out[22]
port 92 nsew signal output
rlabel metal3 s 29200 28508 29800 28748 6 io_out[23]
port 93 nsew signal output
rlabel metal2 s 21886 200 21998 800 6 io_out[24]
port 94 nsew signal output
rlabel metal2 s 19954 49200 20066 49800 6 io_out[25]
port 95 nsew signal output
rlabel metal3 s 200 4028 800 4268 6 io_out[26]
port 96 nsew signal output
rlabel metal2 s 21242 49200 21354 49800 6 io_out[27]
port 97 nsew signal output
rlabel metal2 s 13514 200 13626 800 6 io_out[28]
port 98 nsew signal output
rlabel metal3 s 29200 10828 29800 11068 6 io_out[29]
port 99 nsew signal output
rlabel metal2 s 5786 200 5898 800 6 io_out[2]
port 100 nsew signal output
rlabel metal3 s 200 4708 800 4948 6 io_out[30]
port 101 nsew signal output
rlabel metal3 s 200 11508 800 11748 6 io_out[31]
port 102 nsew signal output
rlabel metal3 s 200 37348 800 37588 6 io_out[32]
port 103 nsew signal output
rlabel metal3 s 29200 15588 29800 15828 6 io_out[33]
port 104 nsew signal output
rlabel metal3 s 29200 42788 29800 43028 6 io_out[34]
port 105 nsew signal output
rlabel metal3 s 29200 40748 29800 40988 6 io_out[35]
port 106 nsew signal output
rlabel metal2 s 2566 49200 2678 49800 6 io_out[36]
port 107 nsew signal output
rlabel metal3 s 29200 46188 29800 46428 6 io_out[37]
port 108 nsew signal output
rlabel metal3 s 200 34628 800 34868 6 io_out[3]
port 109 nsew signal output
rlabel metal3 s 29200 33948 29800 34188 6 io_out[4]
port 110 nsew signal output
rlabel metal2 s 8362 49200 8474 49800 6 io_out[5]
port 111 nsew signal output
rlabel metal2 s 28326 49200 28438 49800 6 io_out[6]
port 112 nsew signal output
rlabel metal3 s 200 15588 800 15828 6 io_out[7]
port 113 nsew signal output
rlabel metal2 s 14802 200 14914 800 6 io_out[8]
port 114 nsew signal output
rlabel metal3 s 200 12188 800 12428 6 io_out[9]
port 115 nsew signal output
rlabel metal3 s 29200 16268 29800 16508 6 la1_data_in[0]
port 116 nsew signal input
rlabel metal2 s 17378 200 17490 800 6 la1_data_in[10]
port 117 nsew signal input
rlabel metal3 s 29200 14908 29800 15148 6 la1_data_in[11]
port 118 nsew signal input
rlabel metal3 s 200 29868 800 30108 6 la1_data_in[12]
port 119 nsew signal input
rlabel metal2 s 27038 200 27150 800 6 la1_data_in[13]
port 120 nsew signal input
rlabel metal3 s 200 10148 800 10388 6 la1_data_in[14]
port 121 nsew signal input
rlabel metal2 s 3210 49200 3322 49800 6 la1_data_in[15]
port 122 nsew signal input
rlabel metal2 s 15446 49200 15558 49800 6 la1_data_in[16]
port 123 nsew signal input
rlabel metal2 s 9650 49200 9762 49800 6 la1_data_in[17]
port 124 nsew signal input
rlabel metal3 s 29200 4708 29800 4948 6 la1_data_in[18]
port 125 nsew signal input
rlabel metal2 s 4498 49200 4610 49800 6 la1_data_in[19]
port 126 nsew signal input
rlabel metal2 s 16090 200 16202 800 6 la1_data_in[1]
port 127 nsew signal input
rlabel metal3 s 200 29188 800 29428 6 la1_data_in[20]
port 128 nsew signal input
rlabel metal2 s 28970 49200 29082 49800 6 la1_data_in[21]
port 129 nsew signal input
rlabel metal3 s 29200 17628 29800 17868 6 la1_data_in[22]
port 130 nsew signal input
rlabel metal3 s 200 628 800 868 6 la1_data_in[23]
port 131 nsew signal input
rlabel metal2 s 11582 200 11694 800 6 la1_data_in[24]
port 132 nsew signal input
rlabel metal3 s 200 30548 800 30788 6 la1_data_in[25]
port 133 nsew signal input
rlabel metal3 s 29200 12868 29800 13108 6 la1_data_in[26]
port 134 nsew signal input
rlabel metal2 s 23174 200 23286 800 6 la1_data_in[27]
port 135 nsew signal input
rlabel metal3 s 200 26468 800 26708 6 la1_data_in[28]
port 136 nsew signal input
rlabel metal3 s 200 40748 800 40988 6 la1_data_in[29]
port 137 nsew signal input
rlabel metal2 s 9006 200 9118 800 6 la1_data_in[2]
port 138 nsew signal input
rlabel metal2 s 1278 200 1390 800 6 la1_data_in[30]
port 139 nsew signal input
rlabel metal3 s 29200 -52 29800 188 6 la1_data_in[31]
port 140 nsew signal input
rlabel metal3 s 200 25108 800 25348 6 la1_data_in[3]
port 141 nsew signal input
rlabel metal2 s 23818 49200 23930 49800 6 la1_data_in[4]
port 142 nsew signal input
rlabel metal3 s 29200 29868 29800 30108 6 la1_data_in[5]
port 143 nsew signal input
rlabel metal2 s 5786 49200 5898 49800 6 la1_data_in[6]
port 144 nsew signal input
rlabel metal3 s 200 18308 800 18548 6 la1_data_in[7]
port 145 nsew signal input
rlabel metal2 s 6430 49200 6542 49800 6 la1_data_in[8]
port 146 nsew signal input
rlabel metal3 s 200 27828 800 28068 6 la1_data_in[9]
port 147 nsew signal input
rlabel metal2 s 6430 200 6542 800 6 la1_data_out[0]
port 148 nsew signal output
rlabel metal3 s 29200 19668 29800 19908 6 la1_data_out[10]
port 149 nsew signal output
rlabel metal2 s 18022 200 18134 800 6 la1_data_out[11]
port 150 nsew signal output
rlabel metal3 s 29200 46868 29800 47108 6 la1_data_out[12]
port 151 nsew signal output
rlabel metal3 s 200 44148 800 44388 6 la1_data_out[13]
port 152 nsew signal output
rlabel metal2 s 11582 49200 11694 49800 6 la1_data_out[14]
port 153 nsew signal output
rlabel metal3 s 200 1308 800 1548 6 la1_data_out[15]
port 154 nsew signal output
rlabel metal3 s 29200 23748 29800 23988 6 la1_data_out[16]
port 155 nsew signal output
rlabel metal3 s 29200 39388 29800 39628 6 la1_data_out[17]
port 156 nsew signal output
rlabel metal3 s 200 44828 800 45068 6 la1_data_out[18]
port 157 nsew signal output
rlabel metal3 s 29200 30548 29800 30788 6 la1_data_out[19]
port 158 nsew signal output
rlabel metal3 s 200 35988 800 36228 6 la1_data_out[1]
port 159 nsew signal output
rlabel metal3 s 200 8108 800 8348 6 la1_data_out[20]
port 160 nsew signal output
rlabel metal3 s 29200 44828 29800 45068 6 la1_data_out[21]
port 161 nsew signal output
rlabel metal2 s 14802 49200 14914 49800 6 la1_data_out[22]
port 162 nsew signal output
rlabel metal2 s 9650 200 9762 800 6 la1_data_out[23]
port 163 nsew signal output
rlabel metal3 s 29200 25108 29800 25348 6 la1_data_out[24]
port 164 nsew signal output
rlabel metal3 s 200 2668 800 2908 6 la1_data_out[25]
port 165 nsew signal output
rlabel metal3 s 29200 14228 29800 14468 6 la1_data_out[26]
port 166 nsew signal output
rlabel metal3 s 200 38708 800 38948 6 la1_data_out[27]
port 167 nsew signal output
rlabel metal3 s 29200 5388 29800 5628 6 la1_data_out[28]
port 168 nsew signal output
rlabel metal2 s 4498 200 4610 800 6 la1_data_out[29]
port 169 nsew signal output
rlabel metal2 s 16734 200 16846 800 6 la1_data_out[2]
port 170 nsew signal output
rlabel metal3 s 29200 20348 29800 20588 6 la1_data_out[30]
port 171 nsew signal output
rlabel metal3 s 29200 48908 29800 49148 6 la1_data_out[31]
port 172 nsew signal output
rlabel metal3 s 200 7428 800 7668 6 la1_data_out[3]
port 173 nsew signal output
rlabel metal3 s 29200 6748 29800 6988 6 la1_data_out[4]
port 174 nsew signal output
rlabel metal2 s 2566 200 2678 800 6 la1_data_out[5]
port 175 nsew signal output
rlabel metal3 s 29200 26468 29800 26708 6 la1_data_out[6]
port 176 nsew signal output
rlabel metal2 s 634 200 746 800 6 la1_data_out[7]
port 177 nsew signal output
rlabel metal3 s 29200 40068 29800 40308 6 la1_data_out[8]
port 178 nsew signal output
rlabel metal2 s 27682 49200 27794 49800 6 la1_data_out[9]
port 179 nsew signal output
rlabel metal3 s 29200 9468 29800 9708 6 la1_oenb[0]
port 180 nsew signal input
rlabel metal2 s 26394 49200 26506 49800 6 la1_oenb[10]
port 181 nsew signal input
rlabel metal3 s 200 22388 800 22628 6 la1_oenb[11]
port 182 nsew signal input
rlabel metal3 s 200 23748 800 23988 6 la1_oenb[12]
port 183 nsew signal input
rlabel metal2 s 23818 200 23930 800 6 la1_oenb[13]
port 184 nsew signal input
rlabel metal2 s -10 200 102 800 6 la1_oenb[14]
port 185 nsew signal input
rlabel metal2 s 28326 200 28438 800 6 la1_oenb[15]
port 186 nsew signal input
rlabel metal3 s 200 28508 800 28748 6 la1_oenb[16]
port 187 nsew signal input
rlabel metal3 s 200 42788 800 43028 6 la1_oenb[17]
port 188 nsew signal input
rlabel metal2 s 7718 49200 7830 49800 6 la1_oenb[18]
port 189 nsew signal input
rlabel metal3 s 200 21028 800 21268 6 la1_oenb[19]
port 190 nsew signal input
rlabel metal2 s 7074 200 7186 800 6 la1_oenb[1]
port 191 nsew signal input
rlabel metal2 s 1922 200 2034 800 6 la1_oenb[20]
port 192 nsew signal input
rlabel metal2 s 16090 49200 16202 49800 6 la1_oenb[21]
port 193 nsew signal input
rlabel metal2 s 7074 49200 7186 49800 6 la1_oenb[22]
port 194 nsew signal input
rlabel metal2 s 19310 200 19422 800 6 la1_oenb[23]
port 195 nsew signal input
rlabel metal2 s 21886 49200 21998 49800 6 la1_oenb[24]
port 196 nsew signal input
rlabel metal3 s 29200 18308 29800 18548 6 la1_oenb[25]
port 197 nsew signal input
rlabel metal3 s 200 31228 800 31468 6 la1_oenb[26]
port 198 nsew signal input
rlabel metal3 s 29200 38028 29800 38268 6 la1_oenb[27]
port 199 nsew signal input
rlabel metal2 s 7718 200 7830 800 6 la1_oenb[28]
port 200 nsew signal input
rlabel metal2 s 14158 200 14270 800 6 la1_oenb[29]
port 201 nsew signal input
rlabel metal3 s 200 6748 800 6988 6 la1_oenb[2]
port 202 nsew signal input
rlabel metal3 s 29200 37348 29800 37588 6 la1_oenb[30]
port 203 nsew signal input
rlabel metal2 s 22530 200 22642 800 6 la1_oenb[31]
port 204 nsew signal input
rlabel metal2 s 18022 49200 18134 49800 6 la1_oenb[3]
port 205 nsew signal input
rlabel metal2 s 17378 49200 17490 49800 6 la1_oenb[4]
port 206 nsew signal input
rlabel metal3 s 200 39388 800 39628 6 la1_oenb[5]
port 207 nsew signal input
rlabel metal3 s 200 46188 800 46428 6 la1_oenb[6]
port 208 nsew signal input
rlabel metal2 s 27682 200 27794 800 6 la1_oenb[7]
port 209 nsew signal input
rlabel metal3 s 200 9468 800 9708 6 la1_oenb[8]
port 210 nsew signal input
rlabel metal3 s 200 33948 800 34188 6 la1_oenb[9]
port 211 nsew signal input
rlabel metal4 s 4417 2128 4737 47376 6 vccd1
port 212 nsew power bidirectional
rlabel metal4 s 11363 2128 11683 47376 6 vccd1
port 212 nsew power bidirectional
rlabel metal4 s 18309 2128 18629 47376 6 vccd1
port 212 nsew power bidirectional
rlabel metal4 s 25255 2128 25575 47376 6 vccd1
port 212 nsew power bidirectional
rlabel metal4 s 7890 2128 8210 47376 6 vssd1
port 213 nsew ground bidirectional
rlabel metal4 s 14836 2128 15156 47376 6 vssd1
port 213 nsew ground bidirectional
rlabel metal4 s 21782 2128 22102 47376 6 vssd1
port 213 nsew ground bidirectional
rlabel metal4 s 28728 2128 29048 47376 6 vssd1
port 213 nsew ground bidirectional
rlabel metal3 s 29200 29188 29800 29428 6 wb_clk_i
port 214 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 30000 50000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 2227630
string GDS_FILE /openlane/designs/wrapped_frequency_counter/runs/RUN_2022.12.16_09.38.01/results/signoff/wrapped_frequency_counter.magic.gds
string GDS_START 434220
<< end >>

