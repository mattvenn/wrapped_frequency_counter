magic
tech sky130A
magscale 1 2
timestamp 1671720230
<< viali >>
rect 21465 47141 21499 47175
rect 1961 47073 1995 47107
rect 10333 47073 10367 47107
rect 23213 47073 23247 47107
rect 26617 47073 26651 47107
rect 3433 47005 3467 47039
rect 5825 47005 5859 47039
rect 6561 47005 6595 47039
rect 7757 47005 7791 47039
rect 9321 47005 9355 47039
rect 11713 47005 11747 47039
rect 13185 47005 13219 47039
rect 14473 47005 14507 47039
rect 16865 47005 16899 47039
rect 18521 47005 18555 47039
rect 20821 47005 20855 47039
rect 22201 47005 22235 47039
rect 24777 47005 24811 47039
rect 27353 47005 27387 47039
rect 27813 47005 27847 47039
rect 3249 46937 3283 46971
rect 9505 46937 9539 46971
rect 22385 46937 22419 46971
rect 24961 46937 24995 46971
rect 27905 46937 27939 46971
rect 6009 46869 6043 46903
rect 6745 46869 6779 46903
rect 24961 46597 24995 46631
rect 7021 46529 7055 46563
rect 13921 46529 13955 46563
rect 14381 46529 14415 46563
rect 16865 46529 16899 46563
rect 19165 46529 19199 46563
rect 22017 46529 22051 46563
rect 27169 46529 27203 46563
rect 2513 46461 2547 46495
rect 2973 46461 3007 46495
rect 3157 46461 3191 46495
rect 4169 46461 4203 46495
rect 7205 46461 7239 46495
rect 8401 46461 8435 46495
rect 9321 46461 9355 46495
rect 9505 46461 9539 46495
rect 10977 46461 11011 46495
rect 13461 46461 13495 46495
rect 13737 46461 13771 46495
rect 14565 46461 14599 46495
rect 14841 46461 14875 46495
rect 17049 46461 17083 46495
rect 17325 46461 17359 46495
rect 19349 46461 19383 46495
rect 19625 46461 19659 46495
rect 22201 46461 22235 46495
rect 22477 46461 22511 46495
rect 24777 46461 24811 46495
rect 26617 46461 26651 46495
rect 27813 46393 27847 46427
rect 1685 46325 1719 46359
rect 27261 46325 27295 46359
rect 4077 46121 4111 46155
rect 7849 46121 7883 46155
rect 9873 46121 9907 46155
rect 10517 46121 10551 46155
rect 13553 46121 13587 46155
rect 14565 46121 14599 46155
rect 16405 46121 16439 46155
rect 18521 46121 18555 46155
rect 1593 45985 1627 46019
rect 2973 45985 3007 46019
rect 11161 45985 11195 46019
rect 11805 45985 11839 46019
rect 19993 45985 20027 46019
rect 22109 45985 22143 46019
rect 22569 45985 22603 46019
rect 26985 45985 27019 46019
rect 27445 45985 27479 46019
rect 4169 45917 4203 45951
rect 7941 45917 7975 45951
rect 9965 45917 9999 45951
rect 10609 45917 10643 45951
rect 13645 45917 13679 45951
rect 14473 45917 14507 45951
rect 16321 45911 16355 45945
rect 18429 45917 18463 45951
rect 19441 45917 19475 45951
rect 24777 45917 24811 45951
rect 27905 45917 27939 45951
rect 1777 45849 1811 45883
rect 11345 45849 11379 45883
rect 19625 45849 19659 45883
rect 22293 45849 22327 45883
rect 27261 45849 27295 45883
rect 24593 45781 24627 45815
rect 1961 45577 1995 45611
rect 11805 45577 11839 45611
rect 19441 45577 19475 45611
rect 22385 45577 22419 45611
rect 27261 45577 27295 45611
rect 2605 45509 2639 45543
rect 23029 45509 23063 45543
rect 26433 45509 26467 45543
rect 2053 45441 2087 45475
rect 2513 45441 2547 45475
rect 3341 45441 3375 45475
rect 9689 45441 9723 45475
rect 10333 45441 10367 45475
rect 11897 45441 11931 45475
rect 19349 45441 19383 45475
rect 19993 45441 20027 45475
rect 20637 45441 20671 45475
rect 20729 45441 20763 45475
rect 22477 45441 22511 45475
rect 23121 45441 23155 45475
rect 24317 45441 24351 45475
rect 26617 45441 26651 45475
rect 27353 45441 27387 45475
rect 27905 45441 27939 45475
rect 26157 45373 26191 45407
rect 27997 45237 28031 45271
rect 22477 45033 22511 45067
rect 24777 45033 24811 45067
rect 25329 45033 25363 45067
rect 28365 44897 28399 44931
rect 2237 44829 2271 44863
rect 3249 44829 3283 44863
rect 25421 44829 25455 44863
rect 25881 44829 25915 44863
rect 26525 44829 26559 44863
rect 26709 44761 26743 44795
rect 27261 44489 27295 44523
rect 26433 44421 26467 44455
rect 2329 44353 2363 44387
rect 3157 44353 3191 44387
rect 27353 44353 27387 44387
rect 27813 44353 27847 44387
rect 3341 44285 3375 44319
rect 3617 44285 3651 44319
rect 26065 44285 26099 44319
rect 26617 44285 26651 44319
rect 2237 44149 2271 44183
rect 4077 43945 4111 43979
rect 1593 43809 1627 43843
rect 3433 43809 3467 43843
rect 25881 43809 25915 43843
rect 26341 43809 26375 43843
rect 4169 43741 4203 43775
rect 4629 43741 4663 43775
rect 28181 43741 28215 43775
rect 3249 43673 3283 43707
rect 26065 43673 26099 43707
rect 25973 43401 26007 43435
rect 1961 43333 1995 43367
rect 3617 43333 3651 43367
rect 3801 43265 3835 43299
rect 25881 43265 25915 43299
rect 27445 43265 27479 43299
rect 27353 43061 27387 43095
rect 28089 43061 28123 43095
rect 2513 42721 2547 42755
rect 28365 42721 28399 42755
rect 1961 42653 1995 42687
rect 2421 42653 2455 42687
rect 26525 42585 26559 42619
rect 28181 42585 28215 42619
rect 27813 42313 27847 42347
rect 26433 42245 26467 42279
rect 2421 42177 2455 42211
rect 26617 42177 26651 42211
rect 27721 42177 27755 42211
rect 26065 42109 26099 42143
rect 1777 41973 1811 42007
rect 2513 41973 2547 42007
rect 1593 41633 1627 41667
rect 3249 41633 3283 41667
rect 3433 41633 3467 41667
rect 27537 41633 27571 41667
rect 26525 41565 26559 41599
rect 26709 41497 26743 41531
rect 1685 41089 1719 41123
rect 27905 41089 27939 41123
rect 1869 41021 1903 41055
rect 2789 41021 2823 41055
rect 27169 40885 27203 40919
rect 2237 40681 2271 40715
rect 26525 40545 26559 40579
rect 28365 40545 28399 40579
rect 2329 40477 2363 40511
rect 26709 40409 26743 40443
rect 27353 40001 27387 40035
rect 27445 40001 27479 40035
rect 1777 39797 1811 39831
rect 27905 39797 27939 39831
rect 26525 39457 26559 39491
rect 28365 39457 28399 39491
rect 1961 39389 1995 39423
rect 2605 39389 2639 39423
rect 3249 39389 3283 39423
rect 26709 39321 26743 39355
rect 1869 39253 1903 39287
rect 3157 39253 3191 39287
rect 19993 39049 20027 39083
rect 26525 39049 26559 39083
rect 2973 38981 3007 39015
rect 1777 38913 1811 38947
rect 2789 38913 2823 38947
rect 18981 38913 19015 38947
rect 19809 38913 19843 38947
rect 20085 38913 20119 38947
rect 20729 38913 20763 38947
rect 21189 38913 21223 38947
rect 21373 38913 21407 38947
rect 26433 38913 26467 38947
rect 27353 38913 27387 38947
rect 4261 38845 4295 38879
rect 19165 38777 19199 38811
rect 27813 38777 27847 38811
rect 1593 38709 1627 38743
rect 19625 38709 19659 38743
rect 20545 38709 20579 38743
rect 21281 38709 21315 38743
rect 27261 38709 27295 38743
rect 18705 38505 18739 38539
rect 18889 38505 18923 38539
rect 20361 38505 20395 38539
rect 20545 38505 20579 38539
rect 21189 38505 21223 38539
rect 22201 38505 22235 38539
rect 25973 38505 26007 38539
rect 19993 38437 20027 38471
rect 1593 38369 1627 38403
rect 1777 38369 1811 38403
rect 2789 38369 2823 38403
rect 26525 38369 26559 38403
rect 26709 38369 26743 38403
rect 28365 38369 28399 38403
rect 21833 38301 21867 38335
rect 25881 38301 25915 38335
rect 18521 38233 18555 38267
rect 18737 38233 18771 38267
rect 21005 38233 21039 38267
rect 21221 38233 21255 38267
rect 22017 38233 22051 38267
rect 20361 38165 20395 38199
rect 21373 38165 21407 38199
rect 20361 37961 20395 37995
rect 20269 37893 20303 37927
rect 21249 37893 21283 37927
rect 21465 37893 21499 37927
rect 18429 37825 18463 37859
rect 18613 37825 18647 37859
rect 19073 37825 19107 37859
rect 19257 37825 19291 37859
rect 20085 37825 20119 37859
rect 20453 37825 20487 37859
rect 22017 37825 22051 37859
rect 27353 37825 27387 37859
rect 1685 37757 1719 37791
rect 3341 37757 3375 37791
rect 3525 37757 3559 37791
rect 3985 37757 4019 37791
rect 19165 37757 19199 37791
rect 27721 37757 27755 37791
rect 20637 37689 20671 37723
rect 18521 37621 18555 37655
rect 21097 37621 21131 37655
rect 21281 37621 21315 37655
rect 22201 37621 22235 37655
rect 18245 37417 18279 37451
rect 19625 37417 19659 37451
rect 20453 37417 20487 37451
rect 3065 37281 3099 37315
rect 16865 37281 16899 37315
rect 19717 37281 19751 37315
rect 1777 37213 1811 37247
rect 1869 37213 1903 37247
rect 3249 37213 3283 37247
rect 4813 37213 4847 37247
rect 16957 37213 16991 37247
rect 19993 37213 20027 37247
rect 20637 37213 20671 37247
rect 20913 37213 20947 37247
rect 28365 37213 28399 37247
rect 4169 37145 4203 37179
rect 18061 37145 18095 37179
rect 18277 37145 18311 37179
rect 26525 37145 26559 37179
rect 28181 37145 28215 37179
rect 17049 37077 17083 37111
rect 17417 37077 17451 37111
rect 18429 37077 18463 37111
rect 19441 37077 19475 37111
rect 20821 37077 20855 37111
rect 21373 36873 21407 36907
rect 27905 36873 27939 36907
rect 2605 36737 2639 36771
rect 3249 36737 3283 36771
rect 4721 36737 4755 36771
rect 17049 36737 17083 36771
rect 18429 36737 18463 36771
rect 21465 36737 21499 36771
rect 22201 36737 22235 36771
rect 26361 36737 26395 36771
rect 26617 36737 26651 36771
rect 27353 36737 27387 36771
rect 27813 36737 27847 36771
rect 2421 36669 2455 36703
rect 4077 36669 4111 36703
rect 5549 36669 5583 36703
rect 16865 36669 16899 36703
rect 27169 36601 27203 36635
rect 17233 36533 17267 36567
rect 18613 36533 18647 36567
rect 22477 36533 22511 36567
rect 25237 36533 25271 36567
rect 21465 36329 21499 36363
rect 28273 36329 28307 36363
rect 1961 36193 1995 36227
rect 4813 36193 4847 36227
rect 15853 36193 15887 36227
rect 23581 36193 23615 36227
rect 23765 36193 23799 36227
rect 24777 36193 24811 36227
rect 27445 36193 27479 36227
rect 2421 36125 2455 36159
rect 3985 36125 4019 36159
rect 5549 36125 5583 36159
rect 16957 36125 16991 36159
rect 17785 36125 17819 36159
rect 20085 36125 20119 36159
rect 20352 36125 20386 36159
rect 22661 36125 22695 36159
rect 25789 36125 25823 36159
rect 3249 36057 3283 36091
rect 5917 36057 5951 36091
rect 16129 36057 16163 36091
rect 25973 36057 26007 36091
rect 16037 35989 16071 36023
rect 16497 35989 16531 36023
rect 17141 35989 17175 36023
rect 17601 35989 17635 36023
rect 22477 35989 22511 36023
rect 23121 35989 23155 36023
rect 23489 35989 23523 36023
rect 25329 35989 25363 36023
rect 26249 35785 26283 35819
rect 1685 35717 1719 35751
rect 16313 35717 16347 35751
rect 17132 35717 17166 35751
rect 3525 35649 3559 35683
rect 3985 35649 4019 35683
rect 16129 35649 16163 35683
rect 18705 35649 18739 35683
rect 18961 35649 18995 35683
rect 22385 35649 22419 35683
rect 22652 35649 22686 35683
rect 24225 35649 24259 35683
rect 24492 35649 24526 35683
rect 26341 35649 26375 35683
rect 3341 35581 3375 35615
rect 4353 35581 4387 35615
rect 15945 35581 15979 35615
rect 16865 35581 16899 35615
rect 18245 35513 18279 35547
rect 20085 35445 20119 35479
rect 23765 35445 23799 35479
rect 25605 35445 25639 35479
rect 27169 35445 27203 35479
rect 3065 35241 3099 35275
rect 20821 35241 20855 35275
rect 21281 35241 21315 35275
rect 23489 35241 23523 35275
rect 24777 35241 24811 35275
rect 25421 35241 25455 35275
rect 2421 35105 2455 35139
rect 26525 35105 26559 35139
rect 27537 35105 27571 35139
rect 1593 35037 1627 35071
rect 2973 35037 3007 35071
rect 16865 35037 16899 35071
rect 19441 35037 19475 35071
rect 22394 35037 22428 35071
rect 22661 35037 22695 35071
rect 23121 35037 23155 35071
rect 23305 35037 23339 35071
rect 24593 35037 24627 35071
rect 24777 35037 24811 35071
rect 25237 35037 25271 35071
rect 25881 35037 25915 35071
rect 17132 34969 17166 35003
rect 19708 34969 19742 35003
rect 25973 34969 26007 35003
rect 26709 34969 26743 35003
rect 18245 34901 18279 34935
rect 19441 34697 19475 34731
rect 26617 34697 26651 34731
rect 25504 34629 25538 34663
rect 19533 34561 19567 34595
rect 25237 34561 25271 34595
rect 27721 34561 27755 34595
rect 1685 34493 1719 34527
rect 1869 34493 1903 34527
rect 2789 34493 2823 34527
rect 27169 34357 27203 34391
rect 2145 34153 2179 34187
rect 21097 34153 21131 34187
rect 26709 34017 26743 34051
rect 2237 33949 2271 33983
rect 22477 33949 22511 33983
rect 23121 33949 23155 33983
rect 24685 33949 24719 33983
rect 24869 33949 24903 33983
rect 26249 33949 26283 33983
rect 22210 33881 22244 33915
rect 26433 33881 26467 33915
rect 23029 33813 23063 33847
rect 24777 33813 24811 33847
rect 22201 33609 22235 33643
rect 27261 33609 27295 33643
rect 18981 33541 19015 33575
rect 19197 33541 19231 33575
rect 20361 33541 20395 33575
rect 1777 33473 1811 33507
rect 17969 33473 18003 33507
rect 18245 33473 18279 33507
rect 18337 33473 18371 33507
rect 20177 33473 20211 33507
rect 20453 33473 20487 33507
rect 20545 33473 20579 33507
rect 22017 33473 22051 33507
rect 23397 33473 23431 33507
rect 24041 33473 24075 33507
rect 25809 33473 25843 33507
rect 26065 33473 26099 33507
rect 27353 33473 27387 33507
rect 23949 33405 23983 33439
rect 18061 33337 18095 33371
rect 18521 33269 18555 33303
rect 19165 33269 19199 33303
rect 19349 33269 19383 33303
rect 20729 33269 20763 33303
rect 23213 33269 23247 33303
rect 24685 33269 24719 33303
rect 28089 33269 28123 33303
rect 16957 33065 16991 33099
rect 19441 33065 19475 33099
rect 20729 33065 20763 33099
rect 24041 33065 24075 33099
rect 16221 32929 16255 32963
rect 17417 32929 17451 32963
rect 19901 32929 19935 32963
rect 25145 32929 25179 32963
rect 25237 32929 25271 32963
rect 27537 32929 27571 32963
rect 1685 32861 1719 32895
rect 15301 32861 15335 32895
rect 15485 32861 15519 32895
rect 16129 32861 16163 32895
rect 16349 32861 16383 32895
rect 16865 32861 16899 32895
rect 17141 32861 17175 32895
rect 17233 32861 17267 32895
rect 18061 32861 18095 32895
rect 18429 32861 18463 32895
rect 19625 32861 19659 32895
rect 19809 32861 19843 32895
rect 19993 32861 20027 32895
rect 20177 32861 20211 32895
rect 20637 32861 20671 32895
rect 20913 32861 20947 32895
rect 21005 32861 21039 32895
rect 21189 32861 21223 32895
rect 21649 32861 21683 32895
rect 21925 32861 21959 32895
rect 22661 32861 22695 32895
rect 22928 32861 22962 32895
rect 24869 32861 24903 32895
rect 24961 32861 24995 32895
rect 26525 32861 26559 32895
rect 15945 32793 15979 32827
rect 16221 32793 16255 32827
rect 18153 32793 18187 32827
rect 18245 32793 18279 32827
rect 22109 32793 22143 32827
rect 26709 32793 26743 32827
rect 15485 32725 15519 32759
rect 17877 32725 17911 32759
rect 21741 32725 21775 32759
rect 24685 32725 24719 32759
rect 15961 32521 15995 32555
rect 20545 32521 20579 32555
rect 24317 32521 24351 32555
rect 28089 32521 28123 32555
rect 15301 32453 15335 32487
rect 15761 32453 15795 32487
rect 18337 32453 18371 32487
rect 18935 32453 18969 32487
rect 19073 32453 19107 32487
rect 19165 32453 19199 32487
rect 24409 32453 24443 32487
rect 1685 32385 1719 32419
rect 15117 32385 15151 32419
rect 16865 32385 16899 32419
rect 18061 32385 18095 32419
rect 18153 32385 18187 32419
rect 19257 32385 19291 32419
rect 19993 32385 20027 32419
rect 20085 32385 20119 32419
rect 20269 32385 20303 32419
rect 20361 32385 20395 32419
rect 22017 32385 22051 32419
rect 22284 32385 22318 32419
rect 26617 32385 26651 32419
rect 27353 32385 27387 32419
rect 27997 32385 28031 32419
rect 1869 32317 1903 32351
rect 2789 32317 2823 32351
rect 18337 32317 18371 32351
rect 18797 32317 18831 32351
rect 24501 32317 24535 32351
rect 16129 32249 16163 32283
rect 14933 32181 14967 32215
rect 15945 32181 15979 32215
rect 17049 32181 17083 32215
rect 19441 32181 19475 32215
rect 23397 32181 23431 32215
rect 23949 32181 23983 32215
rect 27445 32181 27479 32215
rect 2053 31977 2087 32011
rect 16221 31977 16255 32011
rect 19533 31977 19567 32011
rect 21649 31977 21683 32011
rect 22109 31977 22143 32011
rect 23305 31977 23339 32011
rect 25605 31909 25639 31943
rect 16129 31841 16163 31875
rect 16957 31841 16991 31875
rect 21005 31841 21039 31875
rect 26709 31841 26743 31875
rect 28365 31841 28399 31875
rect 2145 31773 2179 31807
rect 16221 31773 16255 31807
rect 17213 31773 17247 31807
rect 19441 31773 19475 31807
rect 20729 31773 20763 31807
rect 21557 31773 21591 31807
rect 21833 31773 21867 31807
rect 23489 31773 23523 31807
rect 23673 31773 23707 31807
rect 25329 31773 25363 31807
rect 25421 31773 25455 31807
rect 26525 31773 26559 31807
rect 25605 31705 25639 31739
rect 15853 31637 15887 31671
rect 18337 31637 18371 31671
rect 18429 31433 18463 31467
rect 22661 31433 22695 31467
rect 24317 31433 24351 31467
rect 15853 31297 15887 31331
rect 16037 31297 16071 31331
rect 18337 31297 18371 31331
rect 22569 31297 22603 31331
rect 22753 31297 22787 31331
rect 24225 31297 24259 31331
rect 24409 31297 24443 31331
rect 26350 31297 26384 31331
rect 27445 31297 27479 31331
rect 27537 31297 27571 31331
rect 27629 31297 27663 31331
rect 28181 31297 28215 31331
rect 26617 31229 26651 31263
rect 27353 31229 27387 31263
rect 15945 31093 15979 31127
rect 25237 31093 25271 31127
rect 27169 31093 27203 31127
rect 28273 31093 28307 31127
rect 16037 30889 16071 30923
rect 17877 30889 17911 30923
rect 25421 30889 25455 30923
rect 26065 30889 26099 30923
rect 8493 30753 8527 30787
rect 10793 30753 10827 30787
rect 27445 30753 27479 30787
rect 28181 30753 28215 30787
rect 28365 30753 28399 30787
rect 8401 30685 8435 30719
rect 9137 30685 9171 30719
rect 10977 30685 11011 30719
rect 17969 30685 18003 30719
rect 24869 30685 24903 30719
rect 25053 30685 25087 30719
rect 25237 30685 25271 30719
rect 25881 30685 25915 30719
rect 26065 30685 26099 30719
rect 15853 30617 15887 30651
rect 16053 30617 16087 30651
rect 22569 30617 22603 30651
rect 25145 30617 25179 30651
rect 16221 30549 16255 30583
rect 21281 30549 21315 30583
rect 18245 30345 18279 30379
rect 19901 30277 19935 30311
rect 1593 30209 1627 30243
rect 16129 30209 16163 30243
rect 16865 30209 16899 30243
rect 17121 30209 17155 30243
rect 19993 30209 20027 30243
rect 20821 30209 20855 30243
rect 21005 30209 21039 30243
rect 26617 30209 26651 30243
rect 20177 30141 20211 30175
rect 16313 30073 16347 30107
rect 26433 30073 26467 30107
rect 1777 30005 1811 30039
rect 19533 30005 19567 30039
rect 21005 30005 21039 30039
rect 27905 30005 27939 30039
rect 17693 29801 17727 29835
rect 18337 29801 18371 29835
rect 18705 29801 18739 29835
rect 25145 29801 25179 29835
rect 23397 29733 23431 29767
rect 20545 29665 20579 29699
rect 20821 29665 20855 29699
rect 22661 29665 22695 29699
rect 27537 29665 27571 29699
rect 28365 29665 28399 29699
rect 15853 29597 15887 29631
rect 16037 29597 16071 29631
rect 16589 29597 16623 29631
rect 17785 29597 17819 29631
rect 18245 29597 18279 29631
rect 19441 29597 19475 29631
rect 19625 29597 19659 29631
rect 22845 29597 22879 29631
rect 22937 29597 22971 29631
rect 23673 29597 23707 29631
rect 23397 29529 23431 29563
rect 25329 29529 25363 29563
rect 28181 29529 28215 29563
rect 15945 29461 15979 29495
rect 16773 29461 16807 29495
rect 19533 29461 19567 29495
rect 21925 29461 21959 29495
rect 22937 29461 22971 29495
rect 23581 29461 23615 29495
rect 24961 29461 24995 29495
rect 25129 29461 25163 29495
rect 21182 29257 21216 29291
rect 23949 29257 23983 29291
rect 27721 29257 27755 29291
rect 19993 29189 20027 29223
rect 25421 29189 25455 29223
rect 26157 29189 26191 29223
rect 15853 29121 15887 29155
rect 16037 29121 16071 29155
rect 21005 29121 21039 29155
rect 21097 29121 21131 29155
rect 21281 29121 21315 29155
rect 22109 29121 22143 29155
rect 22376 29121 22410 29155
rect 24225 29121 24259 29155
rect 24317 29121 24351 29155
rect 24409 29121 24443 29155
rect 24593 29121 24627 29155
rect 25237 29121 25271 29155
rect 25881 29121 25915 29155
rect 25973 29121 26007 29155
rect 27629 29121 27663 29155
rect 18245 29053 18279 29087
rect 25053 29053 25087 29087
rect 23489 28985 23523 29019
rect 15945 28917 15979 28951
rect 26157 28917 26191 28951
rect 16129 28713 16163 28747
rect 16313 28713 16347 28747
rect 18245 28713 18279 28747
rect 20821 28713 20855 28747
rect 21649 28713 21683 28747
rect 23949 28713 23983 28747
rect 25145 28713 25179 28747
rect 16865 28577 16899 28611
rect 19441 28577 19475 28611
rect 26065 28577 26099 28611
rect 15761 28509 15795 28543
rect 17121 28509 17155 28543
rect 19697 28509 19731 28543
rect 21465 28509 21499 28543
rect 23673 28509 23707 28543
rect 23949 28509 23983 28543
rect 24869 28509 24903 28543
rect 24961 28509 24995 28543
rect 25237 28509 25271 28543
rect 16129 28441 16163 28475
rect 23765 28441 23799 28475
rect 26310 28441 26344 28475
rect 24869 28373 24903 28407
rect 27445 28373 27479 28407
rect 19993 28169 20027 28203
rect 24501 28169 24535 28203
rect 26157 28169 26191 28203
rect 18245 28101 18279 28135
rect 1593 28033 1627 28067
rect 18061 28033 18095 28067
rect 18337 28033 18371 28067
rect 18797 28033 18831 28067
rect 18889 28033 18923 28067
rect 19073 28033 19107 28067
rect 19165 28033 19199 28067
rect 19901 28033 19935 28067
rect 23397 28033 23431 28067
rect 23673 28033 23707 28067
rect 24133 28033 24167 28067
rect 25513 28033 25547 28067
rect 25697 28033 25731 28067
rect 25789 28033 25823 28067
rect 25881 28033 25915 28067
rect 27353 28033 27387 28067
rect 27537 28033 27571 28067
rect 24225 27965 24259 27999
rect 23581 27897 23615 27931
rect 1777 27829 1811 27863
rect 17877 27829 17911 27863
rect 19349 27829 19383 27863
rect 23213 27829 23247 27863
rect 24317 27829 24351 27863
rect 27169 27829 27203 27863
rect 27353 27829 27387 27863
rect 28181 27829 28215 27863
rect 25145 27625 25179 27659
rect 18061 27557 18095 27591
rect 22109 27557 22143 27591
rect 15393 27489 15427 27523
rect 19993 27489 20027 27523
rect 27537 27489 27571 27523
rect 28365 27489 28399 27523
rect 16681 27421 16715 27455
rect 21833 27421 21867 27455
rect 22109 27421 22143 27455
rect 23857 27421 23891 27455
rect 24041 27421 24075 27455
rect 25329 27421 25363 27455
rect 25605 27421 25639 27455
rect 15485 27353 15519 27387
rect 15577 27353 15611 27387
rect 16948 27353 16982 27387
rect 20260 27353 20294 27387
rect 21925 27353 21959 27387
rect 25513 27353 25547 27387
rect 28181 27353 28215 27387
rect 15945 27285 15979 27319
rect 21373 27285 21407 27319
rect 23949 27285 23983 27319
rect 17049 27081 17083 27115
rect 25881 27081 25915 27115
rect 27905 27081 27939 27115
rect 15577 27013 15611 27047
rect 15761 27013 15795 27047
rect 18521 27013 18555 27047
rect 18705 27013 18739 27047
rect 22201 27013 22235 27047
rect 22385 27013 22419 27047
rect 15945 26945 15979 26979
rect 16865 26945 16899 26979
rect 18797 26945 18831 26979
rect 21281 26945 21315 26979
rect 21465 26945 21499 26979
rect 26157 26945 26191 26979
rect 27813 26945 27847 26979
rect 25881 26877 25915 26911
rect 22017 26809 22051 26843
rect 18521 26741 18555 26775
rect 21465 26741 21499 26775
rect 26065 26741 26099 26775
rect 27169 26741 27203 26775
rect 19533 26537 19567 26571
rect 23305 26537 23339 26571
rect 17049 26469 17083 26503
rect 21005 26401 21039 26435
rect 21925 26401 21959 26435
rect 26525 26401 26559 26435
rect 28365 26401 28399 26435
rect 1777 26333 1811 26367
rect 16865 26333 16899 26367
rect 19441 26333 19475 26367
rect 21465 26333 21499 26367
rect 22181 26333 22215 26367
rect 24593 26333 24627 26367
rect 21373 26265 21407 26299
rect 26709 26265 26743 26299
rect 21281 26197 21315 26231
rect 24685 26197 24719 26231
rect 15945 25993 15979 26027
rect 18245 25993 18279 26027
rect 21097 25993 21131 26027
rect 27261 25993 27295 26027
rect 23949 25925 23983 25959
rect 26525 25925 26559 25959
rect 1685 25857 1719 25891
rect 16865 25857 16899 25891
rect 17132 25857 17166 25891
rect 18797 25857 18831 25891
rect 19053 25857 19087 25891
rect 21005 25857 21039 25891
rect 24685 25857 24719 25891
rect 24869 25857 24903 25891
rect 25697 25857 25731 25891
rect 26341 25857 26375 25891
rect 26617 25857 26651 25891
rect 27169 25857 27203 25891
rect 1869 25789 1903 25823
rect 2789 25789 2823 25823
rect 15669 25789 15703 25823
rect 15853 25789 15887 25823
rect 21189 25789 21223 25823
rect 25145 25789 25179 25823
rect 26341 25721 26375 25755
rect 16313 25653 16347 25687
rect 20177 25653 20211 25687
rect 20637 25653 20671 25687
rect 22477 25653 22511 25687
rect 25881 25653 25915 25687
rect 27997 25653 28031 25687
rect 2421 25449 2455 25483
rect 17141 25449 17175 25483
rect 18889 25449 18923 25483
rect 20821 25449 20855 25483
rect 23397 25449 23431 25483
rect 24685 25449 24719 25483
rect 25697 25449 25731 25483
rect 21281 25313 21315 25347
rect 23305 25313 23339 25347
rect 24777 25313 24811 25347
rect 27537 25313 27571 25347
rect 28365 25313 28399 25347
rect 1593 25245 1627 25279
rect 2513 25245 2547 25279
rect 16129 25245 16163 25279
rect 16497 25245 16531 25279
rect 16957 25245 16991 25279
rect 18705 25245 18739 25279
rect 19441 25245 19475 25279
rect 19625 25245 19659 25279
rect 19717 25245 19751 25279
rect 21005 25245 21039 25279
rect 21189 25245 21223 25279
rect 23581 25245 23615 25279
rect 24685 25245 24719 25279
rect 25513 25245 25547 25279
rect 25697 25245 25731 25279
rect 16313 25177 16347 25211
rect 28181 25177 28215 25211
rect 1777 25109 1811 25143
rect 23765 25109 23799 25143
rect 25053 25109 25087 25143
rect 22385 24905 22419 24939
rect 28181 24905 28215 24939
rect 22753 24837 22787 24871
rect 25605 24837 25639 24871
rect 22523 24803 22557 24837
rect 17049 24769 17083 24803
rect 23489 24769 23523 24803
rect 23765 24769 23799 24803
rect 24225 24769 24259 24803
rect 24409 24769 24443 24803
rect 25237 24769 25271 24803
rect 25421 24769 25455 24803
rect 25513 24769 25547 24803
rect 25743 24769 25777 24803
rect 25881 24769 25915 24803
rect 26617 24769 26651 24803
rect 27445 24769 27479 24803
rect 28089 24769 28123 24803
rect 26341 24701 26375 24735
rect 27169 24701 27203 24735
rect 27629 24633 27663 24667
rect 16865 24565 16899 24599
rect 22569 24565 22603 24599
rect 23213 24565 23247 24599
rect 23673 24565 23707 24599
rect 24501 24565 24535 24599
rect 26433 24565 26467 24599
rect 26525 24565 26559 24599
rect 27261 24565 27295 24599
rect 18153 24361 18187 24395
rect 15669 24225 15703 24259
rect 26525 24225 26559 24259
rect 28365 24225 28399 24259
rect 15945 24157 15979 24191
rect 16773 24157 16807 24191
rect 17029 24157 17063 24191
rect 18797 24157 18831 24191
rect 21189 24157 21223 24191
rect 21649 24157 21683 24191
rect 22569 24157 22603 24191
rect 22836 24089 22870 24123
rect 26709 24089 26743 24123
rect 15853 24021 15887 24055
rect 16313 24021 16347 24055
rect 18613 24021 18647 24055
rect 21465 24021 21499 24055
rect 21557 24021 21591 24055
rect 23949 24021 23983 24055
rect 17233 23817 17267 23851
rect 20085 23817 20119 23851
rect 22845 23817 22879 23851
rect 24961 23817 24995 23851
rect 25789 23817 25823 23851
rect 26249 23817 26283 23851
rect 16865 23749 16899 23783
rect 17049 23749 17083 23783
rect 18512 23749 18546 23783
rect 22169 23749 22203 23783
rect 22385 23749 22419 23783
rect 21198 23681 21232 23715
rect 23121 23681 23155 23715
rect 23213 23681 23247 23715
rect 23305 23681 23339 23715
rect 23489 23681 23523 23715
rect 24777 23681 24811 23715
rect 25421 23681 25455 23715
rect 25605 23681 25639 23715
rect 26433 23681 26467 23715
rect 26617 23681 26651 23715
rect 27261 23681 27295 23715
rect 18245 23613 18279 23647
rect 21465 23613 21499 23647
rect 24593 23613 24627 23647
rect 19625 23477 19659 23511
rect 22017 23477 22051 23511
rect 22201 23477 22235 23511
rect 26617 23477 26651 23511
rect 27353 23477 27387 23511
rect 27905 23477 27939 23511
rect 18797 23273 18831 23307
rect 21005 23273 21039 23307
rect 21373 23273 21407 23307
rect 19441 23205 19475 23239
rect 19993 23137 20027 23171
rect 21465 23137 21499 23171
rect 26525 23137 26559 23171
rect 26709 23137 26743 23171
rect 28365 23137 28399 23171
rect 16405 23069 16439 23103
rect 18521 23069 18555 23103
rect 18613 23069 18647 23103
rect 19809 23069 19843 23103
rect 19901 23069 19935 23103
rect 21189 23069 21223 23103
rect 25237 23069 25271 23103
rect 25421 23069 25455 23103
rect 25513 23069 25547 23103
rect 25605 23069 25639 23103
rect 16589 22933 16623 22967
rect 25881 22933 25915 22967
rect 15761 22729 15795 22763
rect 18245 22729 18279 22763
rect 22185 22729 22219 22763
rect 24593 22729 24627 22763
rect 26617 22729 26651 22763
rect 27353 22729 27387 22763
rect 17110 22661 17144 22695
rect 22385 22661 22419 22695
rect 24225 22661 24259 22695
rect 24425 22661 24459 22695
rect 25504 22661 25538 22695
rect 15669 22593 15703 22627
rect 27445 22593 27479 22627
rect 27905 22593 27939 22627
rect 15485 22525 15519 22559
rect 16865 22525 16899 22559
rect 25237 22525 25271 22559
rect 16129 22389 16163 22423
rect 22017 22389 22051 22423
rect 22201 22389 22235 22423
rect 24409 22389 24443 22423
rect 15761 22185 15795 22219
rect 22937 22185 22971 22219
rect 23949 22185 23983 22219
rect 24961 22117 24995 22151
rect 24869 22049 24903 22083
rect 27537 22049 27571 22083
rect 16129 21981 16163 22015
rect 16589 21981 16623 22015
rect 20913 21981 20947 22015
rect 21373 21981 21407 22015
rect 23673 21981 23707 22015
rect 24593 21981 24627 22015
rect 24777 21981 24811 22015
rect 25053 21981 25087 22015
rect 28365 21981 28399 22015
rect 15945 21913 15979 21947
rect 22905 21913 22939 21947
rect 23121 21913 23155 21947
rect 23949 21913 23983 21947
rect 28181 21913 28215 21947
rect 16773 21845 16807 21879
rect 21189 21845 21223 21879
rect 21281 21845 21315 21879
rect 22753 21845 22787 21879
rect 23765 21845 23799 21879
rect 25237 21845 25271 21879
rect 15945 21641 15979 21675
rect 18245 21641 18279 21675
rect 28181 21641 28215 21675
rect 15853 21505 15887 21539
rect 16865 21505 16899 21539
rect 17121 21505 17155 21539
rect 18705 21505 18739 21539
rect 18972 21505 19006 21539
rect 21005 21505 21039 21539
rect 21281 21505 21315 21539
rect 22569 21505 22603 21539
rect 22753 21505 22787 21539
rect 25145 21505 25179 21539
rect 25329 21505 25363 21539
rect 27629 21505 27663 21539
rect 28089 21505 28123 21539
rect 15761 21437 15795 21471
rect 22845 21437 22879 21471
rect 21189 21369 21223 21403
rect 16313 21301 16347 21335
rect 20085 21301 20119 21335
rect 20821 21301 20855 21335
rect 22385 21301 22419 21335
rect 25237 21301 25271 21335
rect 15025 21097 15059 21131
rect 15945 21097 15979 21131
rect 19717 21097 19751 21131
rect 18521 20961 18555 20995
rect 21097 20961 21131 20995
rect 21833 20961 21867 20995
rect 27537 20961 27571 20995
rect 16313 20893 16347 20927
rect 18705 20893 18739 20927
rect 20830 20893 20864 20927
rect 22100 20893 22134 20927
rect 25421 20893 25455 20927
rect 25605 20893 25639 20927
rect 25697 20893 25731 20927
rect 25835 20893 25869 20927
rect 28365 20893 28399 20927
rect 15209 20825 15243 20859
rect 15393 20825 15427 20859
rect 16129 20825 16163 20859
rect 28181 20825 28215 20859
rect 18889 20757 18923 20791
rect 23213 20757 23247 20791
rect 26065 20757 26099 20791
rect 12633 20553 12667 20587
rect 18889 20553 18923 20587
rect 19533 20553 19567 20587
rect 19901 20553 19935 20587
rect 22477 20553 22511 20587
rect 28181 20553 28215 20587
rect 14749 20485 14783 20519
rect 19993 20485 20027 20519
rect 2513 20417 2547 20451
rect 12817 20417 12851 20451
rect 13001 20417 13035 20451
rect 13093 20417 13127 20451
rect 14657 20417 14691 20451
rect 14933 20417 14967 20451
rect 18705 20417 18739 20451
rect 22293 20417 22327 20451
rect 22385 20417 22419 20451
rect 23765 20417 23799 20451
rect 25053 20417 25087 20451
rect 25237 20417 25271 20451
rect 25329 20417 25363 20451
rect 25421 20417 25455 20451
rect 28089 20417 28123 20451
rect 20085 20349 20119 20383
rect 22753 20349 22787 20383
rect 23673 20349 23707 20383
rect 24133 20349 24167 20383
rect 27629 20349 27663 20383
rect 15117 20281 15151 20315
rect 1685 20213 1719 20247
rect 2421 20213 2455 20247
rect 25697 20213 25731 20247
rect 13369 20009 13403 20043
rect 14657 20009 14691 20043
rect 14841 20009 14875 20043
rect 15853 20009 15887 20043
rect 25145 20009 25179 20043
rect 27169 20009 27203 20043
rect 1593 19873 1627 19907
rect 1777 19873 1811 19907
rect 2789 19873 2823 19907
rect 24685 19873 24719 19907
rect 25789 19873 25823 19907
rect 13553 19805 13587 19839
rect 15117 19805 15151 19839
rect 15577 19805 15611 19839
rect 16773 19805 16807 19839
rect 24593 19805 24627 19839
rect 24869 19805 24903 19839
rect 24961 19805 24995 19839
rect 25145 19805 25179 19839
rect 26056 19805 26090 19839
rect 27905 19805 27939 19839
rect 13277 19737 13311 19771
rect 13461 19737 13495 19771
rect 15853 19737 15887 19771
rect 15669 19669 15703 19703
rect 16957 19669 16991 19703
rect 12909 19465 12943 19499
rect 14473 19465 14507 19499
rect 15025 19465 15059 19499
rect 16313 19465 16347 19499
rect 19257 19465 19291 19499
rect 19625 19465 19659 19499
rect 15669 19397 15703 19431
rect 17224 19397 17258 19431
rect 12725 19329 12759 19363
rect 13737 19329 13771 19363
rect 13921 19329 13955 19363
rect 14381 19329 14415 19363
rect 16129 19329 16163 19363
rect 16957 19329 16991 19363
rect 19717 19329 19751 19363
rect 21189 19329 21223 19363
rect 1685 19261 1719 19295
rect 1869 19261 1903 19295
rect 2145 19261 2179 19295
rect 12541 19261 12575 19295
rect 15209 19261 15243 19295
rect 15301 19261 15335 19295
rect 19901 19261 19935 19295
rect 13921 19125 13955 19159
rect 18337 19125 18371 19159
rect 21005 19125 21039 19159
rect 27905 19125 27939 19159
rect 1777 18921 1811 18955
rect 2513 18921 2547 18955
rect 12909 18921 12943 18955
rect 16037 18921 16071 18955
rect 16221 18921 16255 18955
rect 25053 18921 25087 18955
rect 23213 18853 23247 18887
rect 20821 18785 20855 18819
rect 24685 18785 24719 18819
rect 26525 18785 26559 18819
rect 28365 18785 28399 18819
rect 2605 18717 2639 18751
rect 12725 18717 12759 18751
rect 12909 18717 12943 18751
rect 13369 18717 13403 18751
rect 13553 18717 13587 18751
rect 15669 18717 15703 18751
rect 16681 18717 16715 18751
rect 16948 18717 16982 18751
rect 18705 18717 18739 18751
rect 19809 18717 19843 18751
rect 21088 18717 21122 18751
rect 22937 18717 22971 18751
rect 24777 18717 24811 18751
rect 25881 18717 25915 18751
rect 14289 18649 14323 18683
rect 14473 18649 14507 18683
rect 19515 18649 19549 18683
rect 20085 18649 20119 18683
rect 23213 18649 23247 18683
rect 28181 18649 28215 18683
rect 13461 18581 13495 18615
rect 14657 18581 14691 18615
rect 16037 18581 16071 18615
rect 18061 18581 18095 18615
rect 18521 18581 18555 18615
rect 19993 18581 20027 18615
rect 22201 18581 22235 18615
rect 23029 18581 23063 18615
rect 25973 18581 26007 18615
rect 16313 18377 16347 18411
rect 17233 18377 17267 18411
rect 21281 18377 21315 18411
rect 22385 18377 22419 18411
rect 22477 18377 22511 18411
rect 23581 18377 23615 18411
rect 27353 18377 27387 18411
rect 27997 18377 28031 18411
rect 13737 18309 13771 18343
rect 16129 18309 16163 18343
rect 18245 18309 18279 18343
rect 19993 18309 20027 18343
rect 24409 18309 24443 18343
rect 25412 18309 25446 18343
rect 1593 18241 1627 18275
rect 12265 18241 12299 18275
rect 12817 18241 12851 18275
rect 12909 18241 12943 18275
rect 13599 18241 13633 18275
rect 13829 18241 13863 18275
rect 14012 18241 14046 18275
rect 14105 18241 14139 18275
rect 14565 18241 14599 18275
rect 14749 18241 14783 18275
rect 14841 18241 14875 18275
rect 15761 18241 15795 18275
rect 16865 18241 16899 18275
rect 17049 18241 17083 18275
rect 21097 18241 21131 18275
rect 23397 18241 23431 18275
rect 23673 18241 23707 18275
rect 24133 18241 24167 18275
rect 24225 18241 24259 18275
rect 25145 18241 25179 18275
rect 27169 18241 27203 18275
rect 27905 18241 27939 18275
rect 12449 18173 12483 18207
rect 20913 18173 20947 18207
rect 22569 18173 22603 18207
rect 1777 18105 1811 18139
rect 22017 18105 22051 18139
rect 26525 18105 26559 18139
rect 13461 18037 13495 18071
rect 14565 18037 14599 18071
rect 16129 18037 16163 18071
rect 23213 18037 23247 18071
rect 24317 18037 24351 18071
rect 16313 17833 16347 17867
rect 18521 17833 18555 17867
rect 21281 17833 21315 17867
rect 24777 17833 24811 17867
rect 19625 17765 19659 17799
rect 2789 17697 2823 17731
rect 13645 17697 13679 17731
rect 14473 17697 14507 17731
rect 14565 17697 14599 17731
rect 20085 17697 20119 17731
rect 23213 17697 23247 17731
rect 23397 17697 23431 17731
rect 26525 17697 26559 17731
rect 26709 17697 26743 17731
rect 28365 17697 28399 17731
rect 1593 17629 1627 17663
rect 13553 17629 13587 17663
rect 13737 17629 13771 17663
rect 14657 17629 14691 17663
rect 14749 17629 14783 17663
rect 15945 17629 15979 17663
rect 18705 17629 18739 17663
rect 18797 17629 18831 17663
rect 22569 17629 22603 17663
rect 23305 17629 23339 17663
rect 23489 17629 23523 17663
rect 1777 17561 1811 17595
rect 16129 17561 16163 17595
rect 20177 17561 20211 17595
rect 24761 17561 24795 17595
rect 24961 17561 24995 17595
rect 14289 17493 14323 17527
rect 20085 17493 20119 17527
rect 23029 17493 23063 17527
rect 24593 17493 24627 17527
rect 2421 17289 2455 17323
rect 15761 17289 15795 17323
rect 19441 17289 19475 17323
rect 20269 17289 20303 17323
rect 20361 17289 20395 17323
rect 25513 17289 25547 17323
rect 18328 17221 18362 17255
rect 22091 17221 22125 17255
rect 22385 17221 22419 17255
rect 22569 17221 22603 17255
rect 22661 17221 22695 17255
rect 1685 17153 1719 17187
rect 2513 17153 2547 17187
rect 14381 17153 14415 17187
rect 14565 17153 14599 17187
rect 15945 17153 15979 17187
rect 18061 17153 18095 17187
rect 24133 17153 24167 17187
rect 24400 17153 24434 17187
rect 26249 17153 26283 17187
rect 27445 17153 27479 17187
rect 16129 17085 16163 17119
rect 20453 17085 20487 17119
rect 14565 17017 14599 17051
rect 19901 17017 19935 17051
rect 26157 16949 26191 16983
rect 27353 16949 27387 16983
rect 27905 16949 27939 16983
rect 15945 16745 15979 16779
rect 16129 16745 16163 16779
rect 24961 16677 24995 16711
rect 25697 16609 25731 16643
rect 26525 16609 26559 16643
rect 26709 16609 26743 16643
rect 1777 16541 1811 16575
rect 20637 16541 20671 16575
rect 23029 16541 23063 16575
rect 23213 16541 23247 16575
rect 23489 16541 23523 16575
rect 16097 16473 16131 16507
rect 16313 16473 16347 16507
rect 20882 16473 20916 16507
rect 24777 16473 24811 16507
rect 25973 16473 26007 16507
rect 28365 16473 28399 16507
rect 22017 16405 22051 16439
rect 23673 16405 23707 16439
rect 20637 16201 20671 16235
rect 28181 16201 28215 16235
rect 1685 16065 1719 16099
rect 16865 16065 16899 16099
rect 17132 16065 17166 16099
rect 20453 16065 20487 16099
rect 21097 16065 21131 16099
rect 21281 16065 21315 16099
rect 21465 16065 21499 16099
rect 26249 16065 26283 16099
rect 26433 16065 26467 16099
rect 27353 16065 27387 16099
rect 28365 16065 28399 16099
rect 1869 15997 1903 16031
rect 2789 15997 2823 16031
rect 26065 15997 26099 16031
rect 18245 15861 18279 15895
rect 27169 15861 27203 15895
rect 2237 15657 2271 15691
rect 20821 15657 20855 15691
rect 10793 15521 10827 15555
rect 13001 15521 13035 15555
rect 13185 15521 13219 15555
rect 21649 15521 21683 15555
rect 26157 15521 26191 15555
rect 2329 15453 2363 15487
rect 10701 15453 10735 15487
rect 17233 15453 17267 15487
rect 19441 15453 19475 15487
rect 25513 15453 25547 15487
rect 26424 15453 26458 15487
rect 27997 15453 28031 15487
rect 11345 15385 11379 15419
rect 17478 15385 17512 15419
rect 19708 15385 19742 15419
rect 21894 15385 21928 15419
rect 18613 15317 18647 15351
rect 23029 15317 23063 15351
rect 25697 15317 25731 15351
rect 27537 15317 27571 15351
rect 28089 15317 28123 15351
rect 22017 15113 22051 15147
rect 22385 15113 22419 15147
rect 23213 15113 23247 15147
rect 27169 15113 27203 15147
rect 27629 15113 27663 15147
rect 24326 15045 24360 15079
rect 17978 14977 18012 15011
rect 18245 14977 18279 15011
rect 20370 14977 20404 15011
rect 20637 14977 20671 15011
rect 24593 14977 24627 15011
rect 26166 14977 26200 15011
rect 26433 14977 26467 15011
rect 27537 14977 27571 15011
rect 22477 14909 22511 14943
rect 22569 14909 22603 14943
rect 27721 14909 27755 14943
rect 19257 14841 19291 14875
rect 16865 14773 16899 14807
rect 25053 14773 25087 14807
rect 16405 14569 16439 14603
rect 17049 14569 17083 14603
rect 17877 14569 17911 14603
rect 19625 14569 19659 14603
rect 26065 14433 26099 14467
rect 27537 14433 27571 14467
rect 28181 14433 28215 14467
rect 3433 14365 3467 14399
rect 16037 14365 16071 14399
rect 17693 14365 17727 14399
rect 19441 14365 19475 14399
rect 28365 14365 28399 14399
rect 1593 14297 1627 14331
rect 3249 14297 3283 14331
rect 16221 14297 16255 14331
rect 16865 14297 16899 14331
rect 25798 14297 25832 14331
rect 17065 14229 17099 14263
rect 17233 14229 17267 14263
rect 24685 14229 24719 14263
rect 2881 14025 2915 14059
rect 16313 14025 16347 14059
rect 17141 14025 17175 14059
rect 19441 14025 19475 14059
rect 20269 14025 20303 14059
rect 23137 14025 23171 14059
rect 23857 14025 23891 14059
rect 23949 14025 23983 14059
rect 24777 14025 24811 14059
rect 25789 14025 25823 14059
rect 22937 13957 22971 13991
rect 2329 13889 2363 13923
rect 2973 13889 3007 13923
rect 16129 13889 16163 13923
rect 16313 13889 16347 13923
rect 17233 13889 17267 13923
rect 17325 13889 17359 13923
rect 17877 13889 17911 13923
rect 18521 13889 18555 13923
rect 19625 13889 19659 13923
rect 19809 13889 19843 13923
rect 20453 13889 20487 13923
rect 23765 13889 23799 13923
rect 24133 13889 24167 13923
rect 24593 13889 24627 13923
rect 25605 13889 25639 13923
rect 28089 13889 28123 13923
rect 16865 13821 16899 13855
rect 22017 13821 22051 13855
rect 22477 13821 22511 13855
rect 18613 13753 18647 13787
rect 22201 13753 22235 13787
rect 3433 13685 3467 13719
rect 17969 13685 18003 13719
rect 23121 13685 23155 13719
rect 23305 13685 23339 13719
rect 24041 13685 24075 13719
rect 18061 13481 18095 13515
rect 19901 13481 19935 13515
rect 22293 13481 22327 13515
rect 24593 13481 24627 13515
rect 24777 13481 24811 13515
rect 25605 13481 25639 13515
rect 1593 13345 1627 13379
rect 3433 13345 3467 13379
rect 20361 13345 20395 13379
rect 20545 13345 20579 13379
rect 21649 13345 21683 13379
rect 22477 13345 22511 13379
rect 23495 13345 23529 13379
rect 23765 13345 23799 13379
rect 17969 13277 18003 13311
rect 18245 13277 18279 13311
rect 18337 13277 18371 13311
rect 20269 13277 20303 13311
rect 21465 13277 21499 13311
rect 21557 13277 21591 13311
rect 22569 13277 22603 13311
rect 22937 13277 22971 13311
rect 23581 13277 23615 13311
rect 23673 13277 23707 13311
rect 25789 13277 25823 13311
rect 25973 13277 26007 13311
rect 3249 13209 3283 13243
rect 24961 13209 24995 13243
rect 18521 13141 18555 13175
rect 21097 13141 21131 13175
rect 22753 13141 22787 13175
rect 22845 13141 22879 13175
rect 23949 13141 23983 13175
rect 24751 13141 24785 13175
rect 1961 12937 1995 12971
rect 20545 12937 20579 12971
rect 22385 12937 22419 12971
rect 23765 12937 23799 12971
rect 25881 12937 25915 12971
rect 26249 12937 26283 12971
rect 23397 12869 23431 12903
rect 23581 12869 23615 12903
rect 2053 12801 2087 12835
rect 16865 12801 16899 12835
rect 18705 12801 18739 12835
rect 19165 12801 19199 12835
rect 20177 12801 20211 12835
rect 20361 12801 20395 12835
rect 22569 12801 22603 12835
rect 22661 12801 22695 12835
rect 26341 12801 26375 12835
rect 27445 12801 27479 12835
rect 17141 12733 17175 12767
rect 22753 12733 22787 12767
rect 22845 12733 22879 12767
rect 26433 12733 26467 12767
rect 27905 12665 27939 12699
rect 18245 12597 18279 12631
rect 18613 12597 18647 12631
rect 19257 12597 19291 12631
rect 27353 12597 27387 12631
rect 17325 12393 17359 12427
rect 21833 12393 21867 12427
rect 21097 12325 21131 12359
rect 16497 12257 16531 12291
rect 26525 12257 26559 12291
rect 26709 12257 26743 12291
rect 28365 12257 28399 12291
rect 1685 12189 1719 12223
rect 16681 12189 16715 12223
rect 16865 12189 16899 12223
rect 17509 12189 17543 12223
rect 21281 12189 21315 12223
rect 22017 12189 22051 12223
rect 16865 11849 16899 11883
rect 18797 11849 18831 11883
rect 18245 11781 18279 11815
rect 1685 11713 1719 11747
rect 17233 11713 17267 11747
rect 17325 11713 17359 11747
rect 18797 11713 18831 11747
rect 27169 11713 27203 11747
rect 1869 11645 1903 11679
rect 2789 11645 2823 11679
rect 17509 11645 17543 11679
rect 18889 11645 18923 11679
rect 27261 11509 27295 11543
rect 1869 11305 1903 11339
rect 18705 11305 18739 11339
rect 18889 11305 18923 11339
rect 4353 11169 4387 11203
rect 26709 11169 26743 11203
rect 1777 11101 1811 11135
rect 3985 11101 4019 11135
rect 17693 11101 17727 11135
rect 26525 11101 26559 11135
rect 18521 11033 18555 11067
rect 28365 11033 28399 11067
rect 17785 10965 17819 10999
rect 18731 10965 18765 10999
rect 18245 10761 18279 10795
rect 18705 10761 18739 10795
rect 17877 10625 17911 10659
rect 18889 10625 18923 10659
rect 18981 10625 19015 10659
rect 19165 10625 19199 10659
rect 19257 10625 19291 10659
rect 19717 10625 19751 10659
rect 19901 10625 19935 10659
rect 19993 10625 20027 10659
rect 20269 10625 20303 10659
rect 27169 10625 27203 10659
rect 17785 10557 17819 10591
rect 20177 10557 20211 10591
rect 17601 10421 17635 10455
rect 27997 10421 28031 10455
rect 18245 10217 18279 10251
rect 18061 10149 18095 10183
rect 19441 10149 19475 10183
rect 18153 10081 18187 10115
rect 19809 10081 19843 10115
rect 27537 10081 27571 10115
rect 28365 10081 28399 10115
rect 1685 10013 1719 10047
rect 3065 10013 3099 10047
rect 17969 10013 18003 10047
rect 19625 10013 19659 10047
rect 17785 9945 17819 9979
rect 28181 9945 28215 9979
rect 2973 9877 3007 9911
rect 27813 9673 27847 9707
rect 1685 9537 1719 9571
rect 20453 9537 20487 9571
rect 27721 9537 27755 9571
rect 1869 9469 1903 9503
rect 2789 9469 2823 9503
rect 4169 9333 4203 9367
rect 20545 9333 20579 9367
rect 2973 8993 3007 9027
rect 1593 8925 1627 8959
rect 26525 8925 26559 8959
rect 28365 8925 28399 8959
rect 1777 8857 1811 8891
rect 26709 8857 26743 8891
rect 1869 8585 1903 8619
rect 27261 8585 27295 8619
rect 4077 8517 4111 8551
rect 1961 8449 1995 8483
rect 4261 8449 4295 8483
rect 27353 8449 27387 8483
rect 27813 8449 27847 8483
rect 3341 8381 3375 8415
rect 26617 8245 26651 8279
rect 1685 8041 1719 8075
rect 2421 8041 2455 8075
rect 2513 7837 2547 7871
rect 3341 7837 3375 7871
rect 3985 7837 4019 7871
rect 25881 7837 25915 7871
rect 26525 7837 26559 7871
rect 26709 7769 26743 7803
rect 28365 7769 28399 7803
rect 4077 7701 4111 7735
rect 25973 7701 26007 7735
rect 3065 7429 3099 7463
rect 4721 7429 4755 7463
rect 26433 7429 26467 7463
rect 4905 7361 4939 7395
rect 26617 7361 26651 7395
rect 27813 7361 27847 7395
rect 26157 7293 26191 7327
rect 1777 7157 1811 7191
rect 27169 7157 27203 7191
rect 5457 6817 5491 6851
rect 7665 6817 7699 6851
rect 7849 6817 7883 6851
rect 26525 6817 26559 6851
rect 28365 6817 28399 6851
rect 1593 6749 1627 6783
rect 2421 6749 2455 6783
rect 2881 6749 2915 6783
rect 4353 6749 4387 6783
rect 5365 6749 5399 6783
rect 25881 6749 25915 6783
rect 6009 6681 6043 6715
rect 25973 6681 26007 6715
rect 26709 6681 26743 6715
rect 2329 6613 2363 6647
rect 4261 6613 4295 6647
rect 27261 6409 27295 6443
rect 4169 6341 4203 6375
rect 1685 6273 1719 6307
rect 27353 6273 27387 6307
rect 27997 6273 28031 6307
rect 1869 6205 1903 6239
rect 3157 6205 3191 6239
rect 3985 6205 4019 6239
rect 4445 6205 4479 6239
rect 27905 6069 27939 6103
rect 4077 5865 4111 5899
rect 1593 5729 1627 5763
rect 2789 5729 2823 5763
rect 27537 5729 27571 5763
rect 28181 5729 28215 5763
rect 28365 5661 28399 5695
rect 1777 5593 1811 5627
rect 1961 5321 1995 5355
rect 3065 5253 3099 5287
rect 2053 5185 2087 5219
rect 2881 5185 2915 5219
rect 12817 5185 12851 5219
rect 28089 5185 28123 5219
rect 4721 5117 4755 5151
rect 5181 4981 5215 5015
rect 12909 4981 12943 5015
rect 1961 4777 1995 4811
rect 20637 4641 20671 4675
rect 21281 4641 21315 4675
rect 27537 4641 27571 4675
rect 2053 4573 2087 4607
rect 3157 4573 3191 4607
rect 3985 4573 4019 4607
rect 4813 4573 4847 4607
rect 5273 4573 5307 4607
rect 6009 4573 6043 4607
rect 12909 4573 12943 4607
rect 20453 4573 20487 4607
rect 25789 4573 25823 4607
rect 26525 4573 26559 4607
rect 26709 4505 26743 4539
rect 4721 4437 4755 4471
rect 6101 4437 6135 4471
rect 25881 4437 25915 4471
rect 27261 4233 27295 4267
rect 4169 4165 4203 4199
rect 13001 4165 13035 4199
rect 3985 4097 4019 4131
rect 11989 4097 12023 4131
rect 12817 4097 12851 4131
rect 17141 4097 17175 4131
rect 20545 4097 20579 4131
rect 27353 4097 27387 4131
rect 1685 4029 1719 4063
rect 3341 4029 3375 4063
rect 3525 4029 3559 4063
rect 4997 4029 5031 4063
rect 7757 4029 7791 4063
rect 7941 4029 7975 4063
rect 8401 4029 8435 4063
rect 13553 4029 13587 4063
rect 26157 4029 26191 4063
rect 26433 4029 26467 4063
rect 26617 4029 26651 4063
rect 27905 4029 27939 4063
rect 6561 3893 6595 3927
rect 12081 3893 12115 3927
rect 17233 3893 17267 3927
rect 7849 3689 7883 3723
rect 18061 3689 18095 3723
rect 28089 3689 28123 3723
rect 3433 3553 3467 3587
rect 5825 3553 5859 3587
rect 11897 3553 11931 3587
rect 12081 3553 12115 3587
rect 12449 3553 12483 3587
rect 25697 3553 25731 3587
rect 25881 3553 25915 3587
rect 4629 3485 4663 3519
rect 5089 3485 5123 3519
rect 9137 3485 9171 3519
rect 9965 3485 9999 3519
rect 10609 3485 10643 3519
rect 11437 3485 11471 3519
rect 14381 3485 14415 3519
rect 16313 3485 16347 3519
rect 16773 3485 16807 3519
rect 17417 3485 17451 3519
rect 18245 3485 18279 3519
rect 19441 3485 19475 3519
rect 20269 3485 20303 3519
rect 21557 3485 21591 3519
rect 22017 3485 22051 3519
rect 23857 3485 23891 3519
rect 24593 3485 24627 3519
rect 27997 3485 28031 3519
rect 1593 3417 1627 3451
rect 3249 3417 3283 3451
rect 5273 3417 5307 3451
rect 27537 3417 27571 3451
rect 9873 3349 9907 3383
rect 10701 3349 10735 3383
rect 16865 3349 16899 3383
rect 20177 3349 20211 3383
rect 22109 3349 22143 3383
rect 23949 3349 23983 3383
rect 1869 3145 1903 3179
rect 2513 3145 2547 3179
rect 9137 3077 9171 3111
rect 11897 3077 11931 3111
rect 17049 3077 17083 3111
rect 19441 3077 19475 3111
rect 22201 3077 22235 3111
rect 24501 3077 24535 3111
rect 1961 3009 1995 3043
rect 2605 3009 2639 3043
rect 6561 3009 6595 3043
rect 8953 3009 8987 3043
rect 11713 3009 11747 3043
rect 14289 3009 14323 3043
rect 16865 3009 16899 3043
rect 19257 3009 19291 3043
rect 22017 3009 22051 3043
rect 24317 3009 24351 3043
rect 27169 3009 27203 3043
rect 27997 3009 28031 3043
rect 3249 2941 3283 2975
rect 3709 2941 3743 2975
rect 3893 2941 3927 2975
rect 4169 2941 4203 2975
rect 6745 2941 6779 2975
rect 7021 2941 7055 2975
rect 9689 2941 9723 2975
rect 12173 2941 12207 2975
rect 14473 2941 14507 2975
rect 14749 2941 14783 2975
rect 17325 2941 17359 2975
rect 19993 2941 20027 2975
rect 22477 2941 22511 2975
rect 25145 2941 25179 2975
rect 27905 2805 27939 2839
rect 4077 2601 4111 2635
rect 5273 2601 5307 2635
rect 8033 2601 8067 2635
rect 14381 2601 14415 2635
rect 16221 2601 16255 2635
rect 27169 2601 27203 2635
rect 2789 2465 2823 2499
rect 3433 2465 3467 2499
rect 9413 2465 9447 2499
rect 17049 2465 17083 2499
rect 17233 2465 17267 2499
rect 18061 2465 18095 2499
rect 26157 2465 26191 2499
rect 26433 2465 26467 2499
rect 26617 2465 26651 2499
rect 27813 2465 27847 2499
rect 4169 2397 4203 2431
rect 5181 2397 5215 2431
rect 6009 2397 6043 2431
rect 8125 2397 8159 2431
rect 9137 2397 9171 2431
rect 14289 2397 14323 2431
rect 27353 2397 27387 2431
rect 3249 2329 3283 2363
rect 5917 2329 5951 2363
rect 16129 2329 16163 2363
<< metal1 >>
rect 14 47404 20 47456
rect 72 47444 78 47456
rect 934 47444 940 47456
rect 72 47416 940 47444
rect 72 47404 78 47416
rect 934 47404 940 47416
rect 992 47404 998 47456
rect 1104 47354 28888 47376
rect 1104 47302 4423 47354
rect 4475 47302 4487 47354
rect 4539 47302 4551 47354
rect 4603 47302 4615 47354
rect 4667 47302 4679 47354
rect 4731 47302 11369 47354
rect 11421 47302 11433 47354
rect 11485 47302 11497 47354
rect 11549 47302 11561 47354
rect 11613 47302 11625 47354
rect 11677 47302 18315 47354
rect 18367 47302 18379 47354
rect 18431 47302 18443 47354
rect 18495 47302 18507 47354
rect 18559 47302 18571 47354
rect 18623 47302 25261 47354
rect 25313 47302 25325 47354
rect 25377 47302 25389 47354
rect 25441 47302 25453 47354
rect 25505 47302 25517 47354
rect 25569 47302 28888 47354
rect 1104 47280 28888 47302
rect 21453 47175 21511 47181
rect 21453 47141 21465 47175
rect 21499 47172 21511 47175
rect 22186 47172 22192 47184
rect 21499 47144 22192 47172
rect 21499 47141 21511 47144
rect 21453 47135 21511 47141
rect 22186 47132 22192 47144
rect 22244 47132 22250 47184
rect 1946 47104 1952 47116
rect 1907 47076 1952 47104
rect 1946 47064 1952 47076
rect 2004 47064 2010 47116
rect 10318 47104 10324 47116
rect 10279 47076 10324 47104
rect 10318 47064 10324 47076
rect 10376 47064 10382 47116
rect 22462 47104 22468 47116
rect 22204 47076 22468 47104
rect 3421 47039 3479 47045
rect 3421 47005 3433 47039
rect 3467 47036 3479 47039
rect 3510 47036 3516 47048
rect 3467 47008 3516 47036
rect 3467 47005 3479 47008
rect 3421 46999 3479 47005
rect 3510 46996 3516 47008
rect 3568 46996 3574 47048
rect 5810 47036 5816 47048
rect 5771 47008 5816 47036
rect 5810 46996 5816 47008
rect 5868 46996 5874 47048
rect 6454 46996 6460 47048
rect 6512 47036 6518 47048
rect 6549 47039 6607 47045
rect 6549 47036 6561 47039
rect 6512 47008 6561 47036
rect 6512 46996 6518 47008
rect 6549 47005 6561 47008
rect 6595 47005 6607 47039
rect 6549 46999 6607 47005
rect 7006 46996 7012 47048
rect 7064 47036 7070 47048
rect 7745 47039 7803 47045
rect 7745 47036 7757 47039
rect 7064 47008 7757 47036
rect 7064 46996 7070 47008
rect 7745 47005 7757 47008
rect 7791 47005 7803 47039
rect 9306 47036 9312 47048
rect 9267 47008 9312 47036
rect 7745 46999 7803 47005
rect 9306 46996 9312 47008
rect 9364 46996 9370 47048
rect 11698 47036 11704 47048
rect 11659 47008 11704 47036
rect 11698 46996 11704 47008
rect 11756 46996 11762 47048
rect 13173 47039 13231 47045
rect 13173 47005 13185 47039
rect 13219 47036 13231 47039
rect 13906 47036 13912 47048
rect 13219 47008 13912 47036
rect 13219 47005 13231 47008
rect 13173 46999 13231 47005
rect 13906 46996 13912 47008
rect 13964 46996 13970 47048
rect 14366 46996 14372 47048
rect 14424 47036 14430 47048
rect 14461 47039 14519 47045
rect 14461 47036 14473 47039
rect 14424 47008 14473 47036
rect 14424 46996 14430 47008
rect 14461 47005 14473 47008
rect 14507 47005 14519 47039
rect 16850 47036 16856 47048
rect 16811 47008 16856 47036
rect 14461 46999 14519 47005
rect 16850 46996 16856 47008
rect 16908 46996 16914 47048
rect 18506 47036 18512 47048
rect 18467 47008 18512 47036
rect 18506 46996 18512 47008
rect 18564 46996 18570 47048
rect 20806 47036 20812 47048
rect 20767 47008 20812 47036
rect 20806 46996 20812 47008
rect 20864 46996 20870 47048
rect 22204 47045 22232 47076
rect 22462 47064 22468 47076
rect 22520 47064 22526 47116
rect 23198 47104 23204 47116
rect 23159 47076 23204 47104
rect 23198 47064 23204 47076
rect 23256 47064 23262 47116
rect 26602 47104 26608 47116
rect 26563 47076 26608 47104
rect 26602 47064 26608 47076
rect 26660 47064 26666 47116
rect 22189 47039 22247 47045
rect 22189 47005 22201 47039
rect 22235 47005 22247 47039
rect 24762 47036 24768 47048
rect 24723 47008 24768 47036
rect 22189 46999 22247 47005
rect 24762 46996 24768 47008
rect 24820 46996 24826 47048
rect 27341 47039 27399 47045
rect 27341 47005 27353 47039
rect 27387 47036 27399 47039
rect 27430 47036 27436 47048
rect 27387 47008 27436 47036
rect 27387 47005 27399 47008
rect 27341 46999 27399 47005
rect 27430 46996 27436 47008
rect 27488 46996 27494 47048
rect 27798 47036 27804 47048
rect 27759 47008 27804 47036
rect 27798 46996 27804 47008
rect 27856 46996 27862 47048
rect 3234 46968 3240 46980
rect 3195 46940 3240 46968
rect 3234 46928 3240 46940
rect 3292 46928 3298 46980
rect 9493 46971 9551 46977
rect 9493 46937 9505 46971
rect 9539 46968 9551 46971
rect 9858 46968 9864 46980
rect 9539 46940 9864 46968
rect 9539 46937 9551 46940
rect 9493 46931 9551 46937
rect 9858 46928 9864 46940
rect 9916 46928 9922 46980
rect 22373 46971 22431 46977
rect 22373 46937 22385 46971
rect 22419 46968 22431 46971
rect 23014 46968 23020 46980
rect 22419 46940 23020 46968
rect 22419 46937 22431 46940
rect 22373 46931 22431 46937
rect 23014 46928 23020 46940
rect 23072 46928 23078 46980
rect 24946 46968 24952 46980
rect 24907 46940 24952 46968
rect 24946 46928 24952 46940
rect 25004 46928 25010 46980
rect 26694 46928 26700 46980
rect 26752 46968 26758 46980
rect 27893 46971 27951 46977
rect 27893 46968 27905 46971
rect 26752 46940 27905 46968
rect 26752 46928 26758 46940
rect 27893 46937 27905 46940
rect 27939 46937 27951 46971
rect 27893 46931 27951 46937
rect 5994 46900 6000 46912
rect 5955 46872 6000 46900
rect 5994 46860 6000 46872
rect 6052 46860 6058 46912
rect 6730 46900 6736 46912
rect 6691 46872 6736 46900
rect 6730 46860 6736 46872
rect 6788 46860 6794 46912
rect 1104 46810 29048 46832
rect 1104 46758 7896 46810
rect 7948 46758 7960 46810
rect 8012 46758 8024 46810
rect 8076 46758 8088 46810
rect 8140 46758 8152 46810
rect 8204 46758 14842 46810
rect 14894 46758 14906 46810
rect 14958 46758 14970 46810
rect 15022 46758 15034 46810
rect 15086 46758 15098 46810
rect 15150 46758 21788 46810
rect 21840 46758 21852 46810
rect 21904 46758 21916 46810
rect 21968 46758 21980 46810
rect 22032 46758 22044 46810
rect 22096 46758 28734 46810
rect 28786 46758 28798 46810
rect 28850 46758 28862 46810
rect 28914 46758 28926 46810
rect 28978 46758 28990 46810
rect 29042 46758 29048 46810
rect 1104 46736 29048 46758
rect 24949 46631 25007 46637
rect 24949 46597 24961 46631
rect 24995 46628 25007 46631
rect 26694 46628 26700 46640
rect 24995 46600 26700 46628
rect 24995 46597 25007 46600
rect 24949 46591 25007 46597
rect 26694 46588 26700 46600
rect 26752 46588 26758 46640
rect 27614 46628 27620 46640
rect 26988 46600 27620 46628
rect 7006 46560 7012 46572
rect 6967 46532 7012 46560
rect 7006 46520 7012 46532
rect 7064 46520 7070 46572
rect 13906 46520 13912 46572
rect 13964 46560 13970 46572
rect 14366 46560 14372 46572
rect 13964 46532 14009 46560
rect 14327 46532 14372 46560
rect 13964 46520 13970 46532
rect 14366 46520 14372 46532
rect 14424 46520 14430 46572
rect 16850 46560 16856 46572
rect 16811 46532 16856 46560
rect 16850 46520 16856 46532
rect 16908 46520 16914 46572
rect 18506 46520 18512 46572
rect 18564 46560 18570 46572
rect 19153 46563 19211 46569
rect 19153 46560 19165 46563
rect 18564 46532 19165 46560
rect 18564 46520 18570 46532
rect 19153 46529 19165 46532
rect 19199 46529 19211 46563
rect 19153 46523 19211 46529
rect 20806 46520 20812 46572
rect 20864 46560 20870 46572
rect 22005 46563 22063 46569
rect 22005 46560 22017 46563
rect 20864 46532 22017 46560
rect 20864 46520 20870 46532
rect 22005 46529 22017 46532
rect 22051 46529 22063 46563
rect 26988 46560 27016 46600
rect 27614 46588 27620 46600
rect 27672 46588 27678 46640
rect 27154 46560 27160 46572
rect 22005 46523 22063 46529
rect 26160 46532 27016 46560
rect 27115 46532 27160 46560
rect 2501 46495 2559 46501
rect 2501 46461 2513 46495
rect 2547 46492 2559 46495
rect 2961 46495 3019 46501
rect 2961 46492 2973 46495
rect 2547 46464 2973 46492
rect 2547 46461 2559 46464
rect 2501 46455 2559 46461
rect 2961 46461 2973 46464
rect 3007 46461 3019 46495
rect 2961 46455 3019 46461
rect 3145 46495 3203 46501
rect 3145 46461 3157 46495
rect 3191 46492 3203 46495
rect 4062 46492 4068 46504
rect 3191 46464 4068 46492
rect 3191 46461 3203 46464
rect 3145 46455 3203 46461
rect 4062 46452 4068 46464
rect 4120 46452 4126 46504
rect 4157 46495 4215 46501
rect 4157 46461 4169 46495
rect 4203 46461 4215 46495
rect 4157 46455 4215 46461
rect 7193 46495 7251 46501
rect 7193 46461 7205 46495
rect 7239 46492 7251 46495
rect 7834 46492 7840 46504
rect 7239 46464 7840 46492
rect 7239 46461 7251 46464
rect 7193 46455 7251 46461
rect 2590 46384 2596 46436
rect 2648 46424 2654 46436
rect 4172 46424 4200 46455
rect 7834 46452 7840 46464
rect 7892 46452 7898 46504
rect 8386 46492 8392 46504
rect 8347 46464 8392 46492
rect 8386 46452 8392 46464
rect 8444 46452 8450 46504
rect 9309 46495 9367 46501
rect 9309 46461 9321 46495
rect 9355 46461 9367 46495
rect 9309 46455 9367 46461
rect 9493 46495 9551 46501
rect 9493 46461 9505 46495
rect 9539 46492 9551 46495
rect 10502 46492 10508 46504
rect 9539 46464 10508 46492
rect 9539 46461 9551 46464
rect 9493 46455 9551 46461
rect 2648 46396 4200 46424
rect 9324 46424 9352 46455
rect 10502 46452 10508 46464
rect 10560 46452 10566 46504
rect 10962 46492 10968 46504
rect 10923 46464 10968 46492
rect 10962 46452 10968 46464
rect 11020 46452 11026 46504
rect 13446 46492 13452 46504
rect 13407 46464 13452 46492
rect 13446 46452 13452 46464
rect 13504 46452 13510 46504
rect 13538 46452 13544 46504
rect 13596 46492 13602 46504
rect 13725 46495 13783 46501
rect 13725 46492 13737 46495
rect 13596 46464 13737 46492
rect 13596 46452 13602 46464
rect 13725 46461 13737 46464
rect 13771 46461 13783 46495
rect 14550 46492 14556 46504
rect 14511 46464 14556 46492
rect 13725 46455 13783 46461
rect 14550 46452 14556 46464
rect 14608 46452 14614 46504
rect 14734 46452 14740 46504
rect 14792 46492 14798 46504
rect 14829 46495 14887 46501
rect 14829 46492 14841 46495
rect 14792 46464 14841 46492
rect 14792 46452 14798 46464
rect 14829 46461 14841 46464
rect 14875 46461 14887 46495
rect 14829 46455 14887 46461
rect 16390 46452 16396 46504
rect 16448 46492 16454 46504
rect 17037 46495 17095 46501
rect 17037 46492 17049 46495
rect 16448 46464 17049 46492
rect 16448 46452 16454 46464
rect 17037 46461 17049 46464
rect 17083 46461 17095 46495
rect 17037 46455 17095 46461
rect 17313 46495 17371 46501
rect 17313 46461 17325 46495
rect 17359 46461 17371 46495
rect 19334 46492 19340 46504
rect 19295 46464 19340 46492
rect 17313 46455 17371 46461
rect 10318 46424 10324 46436
rect 9324 46396 10324 46424
rect 2648 46384 2654 46396
rect 10318 46384 10324 46396
rect 10376 46384 10382 46436
rect 16758 46384 16764 46436
rect 16816 46424 16822 46436
rect 17328 46424 17356 46455
rect 19334 46452 19340 46464
rect 19392 46452 19398 46504
rect 19613 46495 19671 46501
rect 19613 46461 19625 46495
rect 19659 46461 19671 46495
rect 19613 46455 19671 46461
rect 22189 46495 22247 46501
rect 22189 46461 22201 46495
rect 22235 46492 22247 46495
rect 22370 46492 22376 46504
rect 22235 46464 22376 46492
rect 22235 46461 22247 46464
rect 22189 46455 22247 46461
rect 16816 46396 17356 46424
rect 16816 46384 16822 46396
rect 18690 46384 18696 46436
rect 18748 46424 18754 46436
rect 19628 46424 19656 46455
rect 22370 46452 22376 46464
rect 22428 46452 22434 46504
rect 22465 46495 22523 46501
rect 22465 46461 22477 46495
rect 22511 46461 22523 46495
rect 22465 46455 22523 46461
rect 18748 46396 19656 46424
rect 18748 46384 18754 46396
rect 21266 46384 21272 46436
rect 21324 46424 21330 46436
rect 22480 46424 22508 46455
rect 24302 46452 24308 46504
rect 24360 46492 24366 46504
rect 24765 46495 24823 46501
rect 24765 46492 24777 46495
rect 24360 46464 24777 46492
rect 24360 46452 24366 46464
rect 24765 46461 24777 46464
rect 24811 46461 24823 46495
rect 24765 46455 24823 46461
rect 21324 46396 22508 46424
rect 21324 46384 21330 46396
rect 1578 46316 1584 46368
rect 1636 46356 1642 46368
rect 1673 46359 1731 46365
rect 1673 46356 1685 46359
rect 1636 46328 1685 46356
rect 1636 46316 1642 46328
rect 1673 46325 1685 46328
rect 1719 46325 1731 46359
rect 1673 46319 1731 46325
rect 10594 46316 10600 46368
rect 10652 46356 10658 46368
rect 18138 46356 18144 46368
rect 10652 46328 18144 46356
rect 10652 46316 10658 46328
rect 18138 46316 18144 46328
rect 18196 46356 18202 46368
rect 26160 46356 26188 46532
rect 27154 46520 27160 46532
rect 27212 46520 27218 46572
rect 26605 46495 26663 46501
rect 26605 46461 26617 46495
rect 26651 46492 26663 46495
rect 28350 46492 28356 46504
rect 26651 46464 28356 46492
rect 26651 46461 26663 46464
rect 26605 46455 26663 46461
rect 28350 46452 28356 46464
rect 28408 46452 28414 46504
rect 26694 46384 26700 46436
rect 26752 46424 26758 46436
rect 27801 46427 27859 46433
rect 27801 46424 27813 46427
rect 26752 46396 27813 46424
rect 26752 46384 26758 46396
rect 27801 46393 27813 46396
rect 27847 46393 27859 46427
rect 27801 46387 27859 46393
rect 18196 46328 26188 46356
rect 18196 46316 18202 46328
rect 26418 46316 26424 46368
rect 26476 46356 26482 46368
rect 27249 46359 27307 46365
rect 27249 46356 27261 46359
rect 26476 46328 27261 46356
rect 26476 46316 26482 46328
rect 27249 46325 27261 46328
rect 27295 46325 27307 46359
rect 27249 46319 27307 46325
rect 1104 46266 28888 46288
rect 1104 46214 4423 46266
rect 4475 46214 4487 46266
rect 4539 46214 4551 46266
rect 4603 46214 4615 46266
rect 4667 46214 4679 46266
rect 4731 46214 11369 46266
rect 11421 46214 11433 46266
rect 11485 46214 11497 46266
rect 11549 46214 11561 46266
rect 11613 46214 11625 46266
rect 11677 46214 18315 46266
rect 18367 46214 18379 46266
rect 18431 46214 18443 46266
rect 18495 46214 18507 46266
rect 18559 46214 18571 46266
rect 18623 46214 25261 46266
rect 25313 46214 25325 46266
rect 25377 46214 25389 46266
rect 25441 46214 25453 46266
rect 25505 46214 25517 46266
rect 25569 46214 28888 46266
rect 1104 46192 28888 46214
rect 4062 46152 4068 46164
rect 4023 46124 4068 46152
rect 4062 46112 4068 46124
rect 4120 46112 4126 46164
rect 7834 46152 7840 46164
rect 7795 46124 7840 46152
rect 7834 46112 7840 46124
rect 7892 46112 7898 46164
rect 9858 46152 9864 46164
rect 9819 46124 9864 46152
rect 9858 46112 9864 46124
rect 9916 46112 9922 46164
rect 10502 46152 10508 46164
rect 10463 46124 10508 46152
rect 10502 46112 10508 46124
rect 10560 46112 10566 46164
rect 13538 46152 13544 46164
rect 13499 46124 13544 46152
rect 13538 46112 13544 46124
rect 13596 46112 13602 46164
rect 14550 46152 14556 46164
rect 14511 46124 14556 46152
rect 14550 46112 14556 46124
rect 14608 46112 14614 46164
rect 16390 46152 16396 46164
rect 16351 46124 16396 46152
rect 16390 46112 16396 46124
rect 16448 46112 16454 46164
rect 18509 46155 18567 46161
rect 18509 46121 18521 46155
rect 18555 46152 18567 46155
rect 19334 46152 19340 46164
rect 18555 46124 19340 46152
rect 18555 46121 18567 46124
rect 18509 46115 18567 46121
rect 19334 46112 19340 46124
rect 19392 46112 19398 46164
rect 27338 46152 27344 46164
rect 22066 46124 27344 46152
rect 22066 46084 22094 46124
rect 27338 46112 27344 46124
rect 27396 46112 27402 46164
rect 7944 46056 14412 46084
rect 1578 46016 1584 46028
rect 1539 45988 1584 46016
rect 1578 45976 1584 45988
rect 1636 45976 1642 46028
rect 2958 46016 2964 46028
rect 2919 45988 2964 46016
rect 2958 45976 2964 45988
rect 3016 45976 3022 46028
rect 4157 45951 4215 45957
rect 4157 45917 4169 45951
rect 4203 45948 4215 45951
rect 4798 45948 4804 45960
rect 4203 45920 4804 45948
rect 4203 45917 4215 45920
rect 4157 45911 4215 45917
rect 4798 45908 4804 45920
rect 4856 45908 4862 45960
rect 7742 45908 7748 45960
rect 7800 45948 7806 45960
rect 7944 45957 7972 46056
rect 11149 46019 11207 46025
rect 11149 45985 11161 46019
rect 11195 46016 11207 46019
rect 11698 46016 11704 46028
rect 11195 45988 11704 46016
rect 11195 45985 11207 45988
rect 11149 45979 11207 45985
rect 11698 45976 11704 45988
rect 11756 45976 11762 46028
rect 11790 45976 11796 46028
rect 11848 46016 11854 46028
rect 11848 45988 11893 46016
rect 11848 45976 11854 45988
rect 7929 45951 7987 45957
rect 7929 45948 7941 45951
rect 7800 45920 7941 45948
rect 7800 45908 7806 45920
rect 7929 45917 7941 45920
rect 7975 45917 7987 45951
rect 9950 45948 9956 45960
rect 9863 45920 9956 45948
rect 7929 45911 7987 45917
rect 9950 45908 9956 45920
rect 10008 45948 10014 45960
rect 10594 45948 10600 45960
rect 10008 45920 10600 45948
rect 10008 45908 10014 45920
rect 10594 45908 10600 45920
rect 10652 45908 10658 45960
rect 13630 45948 13636 45960
rect 13591 45920 13636 45948
rect 13630 45908 13636 45920
rect 13688 45908 13694 45960
rect 1765 45883 1823 45889
rect 1765 45849 1777 45883
rect 1811 45880 1823 45883
rect 1946 45880 1952 45892
rect 1811 45852 1952 45880
rect 1811 45849 1823 45852
rect 1765 45843 1823 45849
rect 1946 45840 1952 45852
rect 2004 45840 2010 45892
rect 11333 45883 11391 45889
rect 11333 45849 11345 45883
rect 11379 45880 11391 45883
rect 11790 45880 11796 45892
rect 11379 45852 11796 45880
rect 11379 45849 11391 45852
rect 11333 45843 11391 45849
rect 11790 45840 11796 45852
rect 11848 45840 11854 45892
rect 14384 45812 14412 46056
rect 14476 46056 22094 46084
rect 14476 45960 14504 46056
rect 22186 46044 22192 46096
rect 22244 46044 22250 46096
rect 19978 46016 19984 46028
rect 19939 45988 19984 46016
rect 19978 45976 19984 45988
rect 20036 45976 20042 46028
rect 22097 46019 22155 46025
rect 22097 45985 22109 46019
rect 22143 46016 22155 46019
rect 22204 46016 22232 46044
rect 22554 46016 22560 46028
rect 22143 45988 22232 46016
rect 22515 45988 22560 46016
rect 22143 45985 22155 45988
rect 22097 45979 22155 45985
rect 22554 45976 22560 45988
rect 22612 45976 22618 46028
rect 26973 46019 27031 46025
rect 26973 45985 26985 46019
rect 27019 46016 27031 46019
rect 27062 46016 27068 46028
rect 27019 45988 27068 46016
rect 27019 45985 27031 45988
rect 26973 45979 27031 45985
rect 27062 45976 27068 45988
rect 27120 45976 27126 46028
rect 27430 46016 27436 46028
rect 27391 45988 27436 46016
rect 27430 45976 27436 45988
rect 27488 45976 27494 46028
rect 14458 45908 14464 45960
rect 14516 45948 14522 45960
rect 14516 45920 14609 45948
rect 16309 45945 16367 45951
rect 14516 45908 14522 45920
rect 16309 45911 16321 45945
rect 16355 45942 16367 45945
rect 16355 45914 16436 45942
rect 16355 45911 16367 45914
rect 16309 45905 16367 45911
rect 16408 45812 16436 45914
rect 18138 45908 18144 45960
rect 18196 45948 18202 45960
rect 18417 45951 18475 45957
rect 18417 45948 18429 45951
rect 18196 45920 18429 45948
rect 18196 45908 18202 45920
rect 18417 45917 18429 45920
rect 18463 45917 18475 45951
rect 19426 45948 19432 45960
rect 19387 45920 19432 45948
rect 18417 45911 18475 45917
rect 19426 45908 19432 45920
rect 19484 45908 19490 45960
rect 23842 45908 23848 45960
rect 23900 45948 23906 45960
rect 24765 45951 24823 45957
rect 24765 45948 24777 45951
rect 23900 45920 24777 45948
rect 23900 45908 23906 45920
rect 24765 45917 24777 45920
rect 24811 45917 24823 45951
rect 24765 45911 24823 45917
rect 27522 45908 27528 45960
rect 27580 45948 27586 45960
rect 27893 45951 27951 45957
rect 27893 45948 27905 45951
rect 27580 45920 27905 45948
rect 27580 45908 27586 45920
rect 27893 45917 27905 45920
rect 27939 45917 27951 45951
rect 27893 45911 27951 45917
rect 19610 45880 19616 45892
rect 19571 45852 19616 45880
rect 19610 45840 19616 45852
rect 19668 45840 19674 45892
rect 22278 45880 22284 45892
rect 22239 45852 22284 45880
rect 22278 45840 22284 45852
rect 22336 45840 22342 45892
rect 25130 45880 25136 45892
rect 23492 45852 25136 45880
rect 23492 45812 23520 45852
rect 25130 45840 25136 45852
rect 25188 45840 25194 45892
rect 27246 45880 27252 45892
rect 27207 45852 27252 45880
rect 27246 45840 27252 45852
rect 27304 45840 27310 45892
rect 14384 45784 23520 45812
rect 23566 45772 23572 45824
rect 23624 45812 23630 45824
rect 24581 45815 24639 45821
rect 24581 45812 24593 45815
rect 23624 45784 24593 45812
rect 23624 45772 23630 45784
rect 24581 45781 24593 45784
rect 24627 45781 24639 45815
rect 24581 45775 24639 45781
rect 1104 45722 29048 45744
rect 1104 45670 7896 45722
rect 7948 45670 7960 45722
rect 8012 45670 8024 45722
rect 8076 45670 8088 45722
rect 8140 45670 8152 45722
rect 8204 45670 14842 45722
rect 14894 45670 14906 45722
rect 14958 45670 14970 45722
rect 15022 45670 15034 45722
rect 15086 45670 15098 45722
rect 15150 45670 21788 45722
rect 21840 45670 21852 45722
rect 21904 45670 21916 45722
rect 21968 45670 21980 45722
rect 22032 45670 22044 45722
rect 22096 45670 28734 45722
rect 28786 45670 28798 45722
rect 28850 45670 28862 45722
rect 28914 45670 28926 45722
rect 28978 45670 28990 45722
rect 29042 45670 29048 45722
rect 1104 45648 29048 45670
rect 1946 45608 1952 45620
rect 1907 45580 1952 45608
rect 1946 45568 1952 45580
rect 2004 45568 2010 45620
rect 11790 45608 11796 45620
rect 2516 45580 3372 45608
rect 11751 45580 11796 45608
rect 2406 45500 2412 45552
rect 2464 45540 2470 45552
rect 2516 45540 2544 45580
rect 2464 45512 2544 45540
rect 2593 45543 2651 45549
rect 2464 45500 2470 45512
rect 2593 45509 2605 45543
rect 2639 45540 2651 45543
rect 3234 45540 3240 45552
rect 2639 45512 3240 45540
rect 2639 45509 2651 45512
rect 2593 45503 2651 45509
rect 3234 45500 3240 45512
rect 3292 45500 3298 45552
rect 3344 45540 3372 45580
rect 11790 45568 11796 45580
rect 11848 45568 11854 45620
rect 19429 45611 19487 45617
rect 19429 45577 19441 45611
rect 19475 45608 19487 45611
rect 19610 45608 19616 45620
rect 19475 45580 19616 45608
rect 19475 45577 19487 45580
rect 19429 45571 19487 45577
rect 19610 45568 19616 45580
rect 19668 45568 19674 45620
rect 22278 45568 22284 45620
rect 22336 45608 22342 45620
rect 22373 45611 22431 45617
rect 22373 45608 22385 45611
rect 22336 45580 22385 45608
rect 22336 45568 22342 45580
rect 22373 45577 22385 45580
rect 22419 45577 22431 45611
rect 27246 45608 27252 45620
rect 27207 45580 27252 45608
rect 22373 45571 22431 45577
rect 27246 45568 27252 45580
rect 27304 45568 27310 45620
rect 27706 45608 27712 45620
rect 27448 45580 27712 45608
rect 13630 45540 13636 45552
rect 3344 45512 13636 45540
rect 13630 45500 13636 45512
rect 13688 45500 13694 45552
rect 23014 45540 23020 45552
rect 19352 45512 22508 45540
rect 22975 45512 23020 45540
rect 2041 45475 2099 45481
rect 2041 45441 2053 45475
rect 2087 45472 2099 45475
rect 2424 45472 2452 45500
rect 19352 45484 19380 45512
rect 2087 45444 2452 45472
rect 2501 45475 2559 45481
rect 2087 45441 2099 45444
rect 2041 45435 2099 45441
rect 2501 45441 2513 45475
rect 2547 45441 2559 45475
rect 2501 45435 2559 45441
rect 3329 45475 3387 45481
rect 3329 45441 3341 45475
rect 3375 45472 3387 45475
rect 3510 45472 3516 45484
rect 3375 45444 3516 45472
rect 3375 45441 3387 45444
rect 3329 45435 3387 45441
rect 2314 45364 2320 45416
rect 2372 45404 2378 45416
rect 2516 45404 2544 45435
rect 3510 45432 3516 45444
rect 3568 45432 3574 45484
rect 9306 45432 9312 45484
rect 9364 45472 9370 45484
rect 9677 45475 9735 45481
rect 9677 45472 9689 45475
rect 9364 45444 9689 45472
rect 9364 45432 9370 45444
rect 9677 45441 9689 45444
rect 9723 45441 9735 45475
rect 10318 45472 10324 45484
rect 10279 45444 10324 45472
rect 9677 45435 9735 45441
rect 10318 45432 10324 45444
rect 10376 45432 10382 45484
rect 11882 45472 11888 45484
rect 11843 45444 11888 45472
rect 11882 45432 11888 45444
rect 11940 45472 11946 45484
rect 19334 45472 19340 45484
rect 11940 45444 12434 45472
rect 19295 45444 19340 45472
rect 11940 45432 11946 45444
rect 9950 45404 9956 45416
rect 2372 45376 9956 45404
rect 2372 45364 2378 45376
rect 9950 45364 9956 45376
rect 10008 45364 10014 45416
rect 12406 45404 12434 45444
rect 19334 45432 19340 45444
rect 19392 45432 19398 45484
rect 19426 45432 19432 45484
rect 19484 45472 19490 45484
rect 19981 45475 20039 45481
rect 19981 45472 19993 45475
rect 19484 45444 19993 45472
rect 19484 45432 19490 45444
rect 19981 45441 19993 45444
rect 20027 45441 20039 45475
rect 20622 45472 20628 45484
rect 20583 45444 20628 45472
rect 19981 45435 20039 45441
rect 20622 45432 20628 45444
rect 20680 45432 20686 45484
rect 20717 45475 20775 45481
rect 20717 45441 20729 45475
rect 20763 45472 20775 45475
rect 22370 45472 22376 45484
rect 20763 45444 22376 45472
rect 20763 45441 20775 45444
rect 20717 45435 20775 45441
rect 22370 45432 22376 45444
rect 22428 45432 22434 45484
rect 22480 45481 22508 45512
rect 23014 45500 23020 45512
rect 23072 45500 23078 45552
rect 26234 45540 26240 45552
rect 23124 45512 26240 45540
rect 23124 45484 23152 45512
rect 26234 45500 26240 45512
rect 26292 45500 26298 45552
rect 26418 45540 26424 45552
rect 26379 45512 26424 45540
rect 26418 45500 26424 45512
rect 26476 45500 26482 45552
rect 22465 45475 22523 45481
rect 22465 45441 22477 45475
rect 22511 45441 22523 45475
rect 23106 45472 23112 45484
rect 23019 45444 23112 45472
rect 22465 45435 22523 45441
rect 23106 45432 23112 45444
rect 23164 45432 23170 45484
rect 24302 45472 24308 45484
rect 24263 45444 24308 45472
rect 24302 45432 24308 45444
rect 24360 45432 24366 45484
rect 26605 45475 26663 45481
rect 26605 45441 26617 45475
rect 26651 45472 26663 45475
rect 26694 45472 26700 45484
rect 26651 45444 26700 45472
rect 26651 45441 26663 45444
rect 26605 45435 26663 45441
rect 26694 45432 26700 45444
rect 26752 45432 26758 45484
rect 27338 45472 27344 45484
rect 27299 45444 27344 45472
rect 27338 45432 27344 45444
rect 27396 45432 27402 45484
rect 25774 45404 25780 45416
rect 12406 45376 25780 45404
rect 25774 45364 25780 45376
rect 25832 45364 25838 45416
rect 26145 45407 26203 45413
rect 26145 45373 26157 45407
rect 26191 45404 26203 45407
rect 27448 45404 27476 45580
rect 27706 45568 27712 45580
rect 27764 45568 27770 45620
rect 27890 45472 27896 45484
rect 27851 45444 27896 45472
rect 27890 45432 27896 45444
rect 27948 45432 27954 45484
rect 26191 45376 27476 45404
rect 26191 45373 26203 45376
rect 26145 45367 26203 45373
rect 20622 45296 20628 45348
rect 20680 45336 20686 45348
rect 27154 45336 27160 45348
rect 20680 45308 27160 45336
rect 20680 45296 20686 45308
rect 27154 45296 27160 45308
rect 27212 45296 27218 45348
rect 26418 45228 26424 45280
rect 26476 45268 26482 45280
rect 27985 45271 28043 45277
rect 27985 45268 27997 45271
rect 26476 45240 27997 45268
rect 26476 45228 26482 45240
rect 27985 45237 27997 45240
rect 28031 45237 28043 45271
rect 27985 45231 28043 45237
rect 1104 45178 28888 45200
rect 1104 45126 4423 45178
rect 4475 45126 4487 45178
rect 4539 45126 4551 45178
rect 4603 45126 4615 45178
rect 4667 45126 4679 45178
rect 4731 45126 11369 45178
rect 11421 45126 11433 45178
rect 11485 45126 11497 45178
rect 11549 45126 11561 45178
rect 11613 45126 11625 45178
rect 11677 45126 18315 45178
rect 18367 45126 18379 45178
rect 18431 45126 18443 45178
rect 18495 45126 18507 45178
rect 18559 45126 18571 45178
rect 18623 45126 25261 45178
rect 25313 45126 25325 45178
rect 25377 45126 25389 45178
rect 25441 45126 25453 45178
rect 25505 45126 25517 45178
rect 25569 45126 28888 45178
rect 1104 45104 28888 45126
rect 22462 45064 22468 45076
rect 22423 45036 22468 45064
rect 22462 45024 22468 45036
rect 22520 45024 22526 45076
rect 24762 45064 24768 45076
rect 24723 45036 24768 45064
rect 24762 45024 24768 45036
rect 24820 45024 24826 45076
rect 24946 45024 24952 45076
rect 25004 45064 25010 45076
rect 25317 45067 25375 45073
rect 25317 45064 25329 45067
rect 25004 45036 25329 45064
rect 25004 45024 25010 45036
rect 25317 45033 25329 45036
rect 25363 45033 25375 45067
rect 25317 45027 25375 45033
rect 26234 45024 26240 45076
rect 26292 45064 26298 45076
rect 27890 45064 27896 45076
rect 26292 45036 27896 45064
rect 26292 45024 26298 45036
rect 27890 45024 27896 45036
rect 27948 45024 27954 45076
rect 4798 44956 4804 45008
rect 4856 44996 4862 45008
rect 23106 44996 23112 45008
rect 4856 44968 23112 44996
rect 4856 44956 4862 44968
rect 23106 44956 23112 44968
rect 23164 44956 23170 45008
rect 27798 44956 27804 45008
rect 27856 44956 27862 45008
rect 25130 44888 25136 44940
rect 25188 44928 25194 44940
rect 25958 44928 25964 44940
rect 25188 44900 25964 44928
rect 25188 44888 25194 44900
rect 2225 44863 2283 44869
rect 2225 44829 2237 44863
rect 2271 44860 2283 44863
rect 3050 44860 3056 44872
rect 2271 44832 3056 44860
rect 2271 44829 2283 44832
rect 2225 44823 2283 44829
rect 3050 44820 3056 44832
rect 3108 44820 3114 44872
rect 3142 44820 3148 44872
rect 3200 44860 3206 44872
rect 25424 44869 25452 44900
rect 25958 44888 25964 44900
rect 26016 44928 26022 44940
rect 27816 44928 27844 44956
rect 28350 44928 28356 44940
rect 26016 44900 27844 44928
rect 28311 44900 28356 44928
rect 26016 44888 26022 44900
rect 28350 44888 28356 44900
rect 28408 44888 28414 44940
rect 3237 44863 3295 44869
rect 3237 44860 3249 44863
rect 3200 44832 3249 44860
rect 3200 44820 3206 44832
rect 3237 44829 3249 44832
rect 3283 44829 3295 44863
rect 3237 44823 3295 44829
rect 25409 44863 25467 44869
rect 25409 44829 25421 44863
rect 25455 44829 25467 44863
rect 25866 44860 25872 44872
rect 25827 44832 25872 44860
rect 25409 44823 25467 44829
rect 25866 44820 25872 44832
rect 25924 44820 25930 44872
rect 26513 44863 26571 44869
rect 26513 44829 26525 44863
rect 26559 44829 26571 44863
rect 26513 44823 26571 44829
rect 26528 44724 26556 44823
rect 26697 44795 26755 44801
rect 26697 44761 26709 44795
rect 26743 44792 26755 44795
rect 27246 44792 27252 44804
rect 26743 44764 27252 44792
rect 26743 44761 26755 44764
rect 26697 44755 26755 44761
rect 27246 44752 27252 44764
rect 27304 44752 27310 44804
rect 27798 44724 27804 44736
rect 26528 44696 27804 44724
rect 27798 44684 27804 44696
rect 27856 44684 27862 44736
rect 1104 44634 29048 44656
rect 1104 44582 7896 44634
rect 7948 44582 7960 44634
rect 8012 44582 8024 44634
rect 8076 44582 8088 44634
rect 8140 44582 8152 44634
rect 8204 44582 14842 44634
rect 14894 44582 14906 44634
rect 14958 44582 14970 44634
rect 15022 44582 15034 44634
rect 15086 44582 15098 44634
rect 15150 44582 21788 44634
rect 21840 44582 21852 44634
rect 21904 44582 21916 44634
rect 21968 44582 21980 44634
rect 22032 44582 22044 44634
rect 22096 44582 28734 44634
rect 28786 44582 28798 44634
rect 28850 44582 28862 44634
rect 28914 44582 28926 44634
rect 28978 44582 28990 44634
rect 29042 44582 29048 44634
rect 1104 44560 29048 44582
rect 27246 44520 27252 44532
rect 27207 44492 27252 44520
rect 27246 44480 27252 44492
rect 27304 44480 27310 44532
rect 26418 44452 26424 44464
rect 26379 44424 26424 44452
rect 26418 44412 26424 44424
rect 26476 44412 26482 44464
rect 2317 44387 2375 44393
rect 2317 44353 2329 44387
rect 2363 44384 2375 44387
rect 2406 44384 2412 44396
rect 2363 44356 2412 44384
rect 2363 44353 2375 44356
rect 2317 44347 2375 44353
rect 2406 44344 2412 44356
rect 2464 44344 2470 44396
rect 3142 44384 3148 44396
rect 3103 44356 3148 44384
rect 3142 44344 3148 44356
rect 3200 44344 3206 44396
rect 26878 44344 26884 44396
rect 26936 44384 26942 44396
rect 27338 44384 27344 44396
rect 26936 44356 27344 44384
rect 26936 44344 26942 44356
rect 27338 44344 27344 44356
rect 27396 44344 27402 44396
rect 27798 44384 27804 44396
rect 27759 44356 27804 44384
rect 27798 44344 27804 44356
rect 27856 44344 27862 44396
rect 3326 44316 3332 44328
rect 3287 44288 3332 44316
rect 3326 44276 3332 44288
rect 3384 44276 3390 44328
rect 3602 44316 3608 44328
rect 3563 44288 3608 44316
rect 3602 44276 3608 44288
rect 3660 44276 3666 44328
rect 26050 44316 26056 44328
rect 26011 44288 26056 44316
rect 26050 44276 26056 44288
rect 26108 44276 26114 44328
rect 26605 44319 26663 44325
rect 26605 44285 26617 44319
rect 26651 44316 26663 44319
rect 27522 44316 27528 44328
rect 26651 44288 27528 44316
rect 26651 44285 26663 44288
rect 26605 44279 26663 44285
rect 27522 44276 27528 44288
rect 27580 44276 27586 44328
rect 2225 44183 2283 44189
rect 2225 44149 2237 44183
rect 2271 44180 2283 44183
rect 3602 44180 3608 44192
rect 2271 44152 3608 44180
rect 2271 44149 2283 44152
rect 2225 44143 2283 44149
rect 3602 44140 3608 44152
rect 3660 44140 3666 44192
rect 1104 44090 28888 44112
rect 1104 44038 4423 44090
rect 4475 44038 4487 44090
rect 4539 44038 4551 44090
rect 4603 44038 4615 44090
rect 4667 44038 4679 44090
rect 4731 44038 11369 44090
rect 11421 44038 11433 44090
rect 11485 44038 11497 44090
rect 11549 44038 11561 44090
rect 11613 44038 11625 44090
rect 11677 44038 18315 44090
rect 18367 44038 18379 44090
rect 18431 44038 18443 44090
rect 18495 44038 18507 44090
rect 18559 44038 18571 44090
rect 18623 44038 25261 44090
rect 25313 44038 25325 44090
rect 25377 44038 25389 44090
rect 25441 44038 25453 44090
rect 25505 44038 25517 44090
rect 25569 44038 28888 44090
rect 1104 44016 28888 44038
rect 3326 43936 3332 43988
rect 3384 43976 3390 43988
rect 4065 43979 4123 43985
rect 4065 43976 4077 43979
rect 3384 43948 4077 43976
rect 3384 43936 3390 43948
rect 4065 43945 4077 43948
rect 4111 43945 4123 43979
rect 4065 43939 4123 43945
rect 106 43800 112 43852
rect 164 43840 170 43852
rect 1581 43843 1639 43849
rect 1581 43840 1593 43843
rect 164 43812 1593 43840
rect 164 43800 170 43812
rect 1581 43809 1593 43812
rect 1627 43809 1639 43843
rect 1581 43803 1639 43809
rect 3050 43800 3056 43852
rect 3108 43840 3114 43852
rect 3421 43843 3479 43849
rect 3421 43840 3433 43843
rect 3108 43812 3433 43840
rect 3108 43800 3114 43812
rect 3421 43809 3433 43812
rect 3467 43809 3479 43843
rect 11882 43840 11888 43852
rect 3421 43803 3479 43809
rect 4172 43812 11888 43840
rect 4172 43784 4200 43812
rect 11882 43800 11888 43812
rect 11940 43800 11946 43852
rect 25866 43840 25872 43852
rect 25827 43812 25872 43840
rect 25866 43800 25872 43812
rect 25924 43800 25930 43852
rect 26142 43800 26148 43852
rect 26200 43840 26206 43852
rect 26329 43843 26387 43849
rect 26329 43840 26341 43843
rect 26200 43812 26341 43840
rect 26200 43800 26206 43812
rect 26329 43809 26341 43812
rect 26375 43809 26387 43843
rect 26329 43803 26387 43809
rect 4154 43772 4160 43784
rect 4115 43744 4160 43772
rect 4154 43732 4160 43744
rect 4212 43732 4218 43784
rect 4614 43772 4620 43784
rect 4575 43744 4620 43772
rect 4614 43732 4620 43744
rect 4672 43732 4678 43784
rect 27246 43732 27252 43784
rect 27304 43772 27310 43784
rect 28169 43775 28227 43781
rect 28169 43772 28181 43775
rect 27304 43744 28181 43772
rect 27304 43732 27310 43744
rect 28169 43741 28181 43744
rect 28215 43741 28227 43775
rect 28169 43735 28227 43741
rect 3234 43704 3240 43716
rect 3195 43676 3240 43704
rect 3234 43664 3240 43676
rect 3292 43664 3298 43716
rect 26050 43704 26056 43716
rect 26011 43676 26056 43704
rect 26050 43664 26056 43676
rect 26108 43664 26114 43716
rect 1104 43546 29048 43568
rect 1104 43494 7896 43546
rect 7948 43494 7960 43546
rect 8012 43494 8024 43546
rect 8076 43494 8088 43546
rect 8140 43494 8152 43546
rect 8204 43494 14842 43546
rect 14894 43494 14906 43546
rect 14958 43494 14970 43546
rect 15022 43494 15034 43546
rect 15086 43494 15098 43546
rect 15150 43494 21788 43546
rect 21840 43494 21852 43546
rect 21904 43494 21916 43546
rect 21968 43494 21980 43546
rect 22032 43494 22044 43546
rect 22096 43494 28734 43546
rect 28786 43494 28798 43546
rect 28850 43494 28862 43546
rect 28914 43494 28926 43546
rect 28978 43494 28990 43546
rect 29042 43494 29048 43546
rect 1104 43472 29048 43494
rect 25961 43435 26019 43441
rect 25961 43401 25973 43435
rect 26007 43432 26019 43435
rect 26050 43432 26056 43444
rect 26007 43404 26056 43432
rect 26007 43401 26019 43404
rect 25961 43395 26019 43401
rect 26050 43392 26056 43404
rect 26108 43392 26114 43444
rect 14 43324 20 43376
rect 72 43364 78 43376
rect 1949 43367 2007 43373
rect 1949 43364 1961 43367
rect 72 43336 1961 43364
rect 72 43324 78 43336
rect 1949 43333 1961 43336
rect 1995 43333 2007 43367
rect 3602 43364 3608 43376
rect 3563 43336 3608 43364
rect 1949 43327 2007 43333
rect 3602 43324 3608 43336
rect 3660 43324 3666 43376
rect 3789 43299 3847 43305
rect 3789 43265 3801 43299
rect 3835 43296 3847 43299
rect 4614 43296 4620 43308
rect 3835 43268 4620 43296
rect 3835 43265 3847 43268
rect 3789 43259 3847 43265
rect 4614 43256 4620 43268
rect 4672 43256 4678 43308
rect 25774 43256 25780 43308
rect 25832 43296 25838 43308
rect 25869 43299 25927 43305
rect 25869 43296 25881 43299
rect 25832 43268 25881 43296
rect 25832 43256 25838 43268
rect 25869 43265 25881 43268
rect 25915 43296 25927 43299
rect 27062 43296 27068 43308
rect 25915 43268 27068 43296
rect 25915 43265 25927 43268
rect 25869 43259 25927 43265
rect 27062 43256 27068 43268
rect 27120 43256 27126 43308
rect 27433 43299 27491 43305
rect 27433 43265 27445 43299
rect 27479 43296 27491 43299
rect 27890 43296 27896 43308
rect 27479 43268 27896 43296
rect 27479 43265 27491 43268
rect 27433 43259 27491 43265
rect 26970 43188 26976 43240
rect 27028 43228 27034 43240
rect 27448 43228 27476 43259
rect 27890 43256 27896 43268
rect 27948 43256 27954 43308
rect 27028 43200 27476 43228
rect 27028 43188 27034 43200
rect 26418 43052 26424 43104
rect 26476 43092 26482 43104
rect 27341 43095 27399 43101
rect 27341 43092 27353 43095
rect 26476 43064 27353 43092
rect 26476 43052 26482 43064
rect 27341 43061 27353 43064
rect 27387 43061 27399 43095
rect 28074 43092 28080 43104
rect 28035 43064 28080 43092
rect 27341 43055 27399 43061
rect 28074 43052 28080 43064
rect 28132 43052 28138 43104
rect 1104 43002 28888 43024
rect 1104 42950 4423 43002
rect 4475 42950 4487 43002
rect 4539 42950 4551 43002
rect 4603 42950 4615 43002
rect 4667 42950 4679 43002
rect 4731 42950 11369 43002
rect 11421 42950 11433 43002
rect 11485 42950 11497 43002
rect 11549 42950 11561 43002
rect 11613 42950 11625 43002
rect 11677 42950 18315 43002
rect 18367 42950 18379 43002
rect 18431 42950 18443 43002
rect 18495 42950 18507 43002
rect 18559 42950 18571 43002
rect 18623 42950 25261 43002
rect 25313 42950 25325 43002
rect 25377 42950 25389 43002
rect 25441 42950 25453 43002
rect 25505 42950 25517 43002
rect 25569 42950 28888 43002
rect 1104 42928 28888 42950
rect 2501 42755 2559 42761
rect 2501 42721 2513 42755
rect 2547 42752 2559 42755
rect 3234 42752 3240 42764
rect 2547 42724 3240 42752
rect 2547 42721 2559 42724
rect 2501 42715 2559 42721
rect 3234 42712 3240 42724
rect 3292 42712 3298 42764
rect 28074 42712 28080 42764
rect 28132 42752 28138 42764
rect 28353 42755 28411 42761
rect 28353 42752 28365 42755
rect 28132 42724 28365 42752
rect 28132 42712 28138 42724
rect 28353 42721 28365 42724
rect 28399 42721 28411 42755
rect 28353 42715 28411 42721
rect 1949 42687 2007 42693
rect 1949 42653 1961 42687
rect 1995 42653 2007 42687
rect 2406 42684 2412 42696
rect 2367 42656 2412 42684
rect 1949 42647 2007 42653
rect 1964 42616 1992 42647
rect 2406 42644 2412 42656
rect 2464 42644 2470 42696
rect 3418 42616 3424 42628
rect 1964 42588 3424 42616
rect 3418 42576 3424 42588
rect 3476 42576 3482 42628
rect 26142 42576 26148 42628
rect 26200 42616 26206 42628
rect 26513 42619 26571 42625
rect 26513 42616 26525 42619
rect 26200 42588 26525 42616
rect 26200 42576 26206 42588
rect 26513 42585 26525 42588
rect 26559 42585 26571 42619
rect 26513 42579 26571 42585
rect 27798 42576 27804 42628
rect 27856 42616 27862 42628
rect 28169 42619 28227 42625
rect 28169 42616 28181 42619
rect 27856 42588 28181 42616
rect 27856 42576 27862 42588
rect 28169 42585 28181 42588
rect 28215 42585 28227 42619
rect 28169 42579 28227 42585
rect 1104 42458 29048 42480
rect 1104 42406 7896 42458
rect 7948 42406 7960 42458
rect 8012 42406 8024 42458
rect 8076 42406 8088 42458
rect 8140 42406 8152 42458
rect 8204 42406 14842 42458
rect 14894 42406 14906 42458
rect 14958 42406 14970 42458
rect 15022 42406 15034 42458
rect 15086 42406 15098 42458
rect 15150 42406 21788 42458
rect 21840 42406 21852 42458
rect 21904 42406 21916 42458
rect 21968 42406 21980 42458
rect 22032 42406 22044 42458
rect 22096 42406 28734 42458
rect 28786 42406 28798 42458
rect 28850 42406 28862 42458
rect 28914 42406 28926 42458
rect 28978 42406 28990 42458
rect 29042 42406 29048 42458
rect 1104 42384 29048 42406
rect 27798 42344 27804 42356
rect 27759 42316 27804 42344
rect 27798 42304 27804 42316
rect 27856 42304 27862 42356
rect 26418 42276 26424 42288
rect 26379 42248 26424 42276
rect 26418 42236 26424 42248
rect 26476 42236 26482 42288
rect 2409 42211 2467 42217
rect 2409 42177 2421 42211
rect 2455 42208 2467 42211
rect 2498 42208 2504 42220
rect 2455 42180 2504 42208
rect 2455 42177 2467 42180
rect 2409 42171 2467 42177
rect 2498 42168 2504 42180
rect 2556 42168 2562 42220
rect 26605 42211 26663 42217
rect 26605 42177 26617 42211
rect 26651 42208 26663 42211
rect 27246 42208 27252 42220
rect 26651 42180 27252 42208
rect 26651 42177 26663 42180
rect 26605 42171 26663 42177
rect 27246 42168 27252 42180
rect 27304 42168 27310 42220
rect 27614 42168 27620 42220
rect 27672 42208 27678 42220
rect 27709 42211 27767 42217
rect 27709 42208 27721 42211
rect 27672 42180 27721 42208
rect 27672 42168 27678 42180
rect 27709 42177 27721 42180
rect 27755 42177 27767 42211
rect 27709 42171 27767 42177
rect 26050 42140 26056 42152
rect 26011 42112 26056 42140
rect 26050 42100 26056 42112
rect 26108 42100 26114 42152
rect 1670 41964 1676 42016
rect 1728 42004 1734 42016
rect 1765 42007 1823 42013
rect 1765 42004 1777 42007
rect 1728 41976 1777 42004
rect 1728 41964 1734 41976
rect 1765 41973 1777 41976
rect 1811 41973 1823 42007
rect 1765 41967 1823 41973
rect 2501 42007 2559 42013
rect 2501 41973 2513 42007
rect 2547 42004 2559 42007
rect 3234 42004 3240 42016
rect 2547 41976 3240 42004
rect 2547 41973 2559 41976
rect 2501 41967 2559 41973
rect 3234 41964 3240 41976
rect 3292 41964 3298 42016
rect 1104 41914 28888 41936
rect 1104 41862 4423 41914
rect 4475 41862 4487 41914
rect 4539 41862 4551 41914
rect 4603 41862 4615 41914
rect 4667 41862 4679 41914
rect 4731 41862 11369 41914
rect 11421 41862 11433 41914
rect 11485 41862 11497 41914
rect 11549 41862 11561 41914
rect 11613 41862 11625 41914
rect 11677 41862 18315 41914
rect 18367 41862 18379 41914
rect 18431 41862 18443 41914
rect 18495 41862 18507 41914
rect 18559 41862 18571 41914
rect 18623 41862 25261 41914
rect 25313 41862 25325 41914
rect 25377 41862 25389 41914
rect 25441 41862 25453 41914
rect 25505 41862 25517 41914
rect 25569 41862 28888 41914
rect 1104 41840 28888 41862
rect 1578 41664 1584 41676
rect 1539 41636 1584 41664
rect 1578 41624 1584 41636
rect 1636 41624 1642 41676
rect 3234 41664 3240 41676
rect 3195 41636 3240 41664
rect 3234 41624 3240 41636
rect 3292 41624 3298 41676
rect 3418 41664 3424 41676
rect 3379 41636 3424 41664
rect 3418 41624 3424 41636
rect 3476 41624 3482 41676
rect 27522 41664 27528 41676
rect 27483 41636 27528 41664
rect 27522 41624 27528 41636
rect 27580 41624 27586 41676
rect 26513 41599 26571 41605
rect 26513 41565 26525 41599
rect 26559 41565 26571 41599
rect 26513 41559 26571 41565
rect 26528 41460 26556 41559
rect 26697 41531 26755 41537
rect 26697 41497 26709 41531
rect 26743 41528 26755 41531
rect 27338 41528 27344 41540
rect 26743 41500 27344 41528
rect 26743 41497 26755 41500
rect 26697 41491 26755 41497
rect 27338 41488 27344 41500
rect 27396 41488 27402 41540
rect 27890 41460 27896 41472
rect 26528 41432 27896 41460
rect 27890 41420 27896 41432
rect 27948 41420 27954 41472
rect 1104 41370 29048 41392
rect 1104 41318 7896 41370
rect 7948 41318 7960 41370
rect 8012 41318 8024 41370
rect 8076 41318 8088 41370
rect 8140 41318 8152 41370
rect 8204 41318 14842 41370
rect 14894 41318 14906 41370
rect 14958 41318 14970 41370
rect 15022 41318 15034 41370
rect 15086 41318 15098 41370
rect 15150 41318 21788 41370
rect 21840 41318 21852 41370
rect 21904 41318 21916 41370
rect 21968 41318 21980 41370
rect 22032 41318 22044 41370
rect 22096 41318 28734 41370
rect 28786 41318 28798 41370
rect 28850 41318 28862 41370
rect 28914 41318 28926 41370
rect 28978 41318 28990 41370
rect 29042 41318 29048 41370
rect 1104 41296 29048 41318
rect 1670 41120 1676 41132
rect 1631 41092 1676 41120
rect 1670 41080 1676 41092
rect 1728 41080 1734 41132
rect 27890 41120 27896 41132
rect 27851 41092 27896 41120
rect 27890 41080 27896 41092
rect 27948 41080 27954 41132
rect 1857 41055 1915 41061
rect 1857 41021 1869 41055
rect 1903 41052 1915 41055
rect 2222 41052 2228 41064
rect 1903 41024 2228 41052
rect 1903 41021 1915 41024
rect 1857 41015 1915 41021
rect 2222 41012 2228 41024
rect 2280 41012 2286 41064
rect 2774 41052 2780 41064
rect 2735 41024 2780 41052
rect 2774 41012 2780 41024
rect 2832 41012 2838 41064
rect 26510 40876 26516 40928
rect 26568 40916 26574 40928
rect 27157 40919 27215 40925
rect 27157 40916 27169 40919
rect 26568 40888 27169 40916
rect 26568 40876 26574 40888
rect 27157 40885 27169 40888
rect 27203 40885 27215 40919
rect 27157 40879 27215 40885
rect 1104 40826 28888 40848
rect 1104 40774 4423 40826
rect 4475 40774 4487 40826
rect 4539 40774 4551 40826
rect 4603 40774 4615 40826
rect 4667 40774 4679 40826
rect 4731 40774 11369 40826
rect 11421 40774 11433 40826
rect 11485 40774 11497 40826
rect 11549 40774 11561 40826
rect 11613 40774 11625 40826
rect 11677 40774 18315 40826
rect 18367 40774 18379 40826
rect 18431 40774 18443 40826
rect 18495 40774 18507 40826
rect 18559 40774 18571 40826
rect 18623 40774 25261 40826
rect 25313 40774 25325 40826
rect 25377 40774 25389 40826
rect 25441 40774 25453 40826
rect 25505 40774 25517 40826
rect 25569 40774 28888 40826
rect 1104 40752 28888 40774
rect 2222 40712 2228 40724
rect 2183 40684 2228 40712
rect 2222 40672 2228 40684
rect 2280 40672 2286 40724
rect 26510 40576 26516 40588
rect 26471 40548 26516 40576
rect 26510 40536 26516 40548
rect 26568 40536 26574 40588
rect 28353 40579 28411 40585
rect 28353 40545 28365 40579
rect 28399 40576 28411 40579
rect 28626 40576 28632 40588
rect 28399 40548 28632 40576
rect 28399 40545 28411 40548
rect 28353 40539 28411 40545
rect 28626 40536 28632 40548
rect 28684 40536 28690 40588
rect 2314 40508 2320 40520
rect 2275 40480 2320 40508
rect 2314 40468 2320 40480
rect 2372 40468 2378 40520
rect 26694 40440 26700 40452
rect 26655 40412 26700 40440
rect 26694 40400 26700 40412
rect 26752 40400 26758 40452
rect 1104 40282 29048 40304
rect 1104 40230 7896 40282
rect 7948 40230 7960 40282
rect 8012 40230 8024 40282
rect 8076 40230 8088 40282
rect 8140 40230 8152 40282
rect 8204 40230 14842 40282
rect 14894 40230 14906 40282
rect 14958 40230 14970 40282
rect 15022 40230 15034 40282
rect 15086 40230 15098 40282
rect 15150 40230 21788 40282
rect 21840 40230 21852 40282
rect 21904 40230 21916 40282
rect 21968 40230 21980 40282
rect 22032 40230 22044 40282
rect 22096 40230 28734 40282
rect 28786 40230 28798 40282
rect 28850 40230 28862 40282
rect 28914 40230 28926 40282
rect 28978 40230 28990 40282
rect 29042 40230 29048 40282
rect 1104 40208 29048 40230
rect 27338 40032 27344 40044
rect 27299 40004 27344 40032
rect 27338 39992 27344 40004
rect 27396 39992 27402 40044
rect 27433 40035 27491 40041
rect 27433 40001 27445 40035
rect 27479 40001 27491 40035
rect 27433 39995 27491 40001
rect 26970 39924 26976 39976
rect 27028 39964 27034 39976
rect 27448 39964 27476 39995
rect 27028 39936 27476 39964
rect 27028 39924 27034 39936
rect 1670 39788 1676 39840
rect 1728 39828 1734 39840
rect 1765 39831 1823 39837
rect 1765 39828 1777 39831
rect 1728 39800 1777 39828
rect 1728 39788 1734 39800
rect 1765 39797 1777 39800
rect 1811 39797 1823 39831
rect 27890 39828 27896 39840
rect 27851 39800 27896 39828
rect 1765 39791 1823 39797
rect 27890 39788 27896 39800
rect 27948 39788 27954 39840
rect 1104 39738 28888 39760
rect 1104 39686 4423 39738
rect 4475 39686 4487 39738
rect 4539 39686 4551 39738
rect 4603 39686 4615 39738
rect 4667 39686 4679 39738
rect 4731 39686 11369 39738
rect 11421 39686 11433 39738
rect 11485 39686 11497 39738
rect 11549 39686 11561 39738
rect 11613 39686 11625 39738
rect 11677 39686 18315 39738
rect 18367 39686 18379 39738
rect 18431 39686 18443 39738
rect 18495 39686 18507 39738
rect 18559 39686 18571 39738
rect 18623 39686 25261 39738
rect 25313 39686 25325 39738
rect 25377 39686 25389 39738
rect 25441 39686 25453 39738
rect 25505 39686 25517 39738
rect 25569 39686 28888 39738
rect 1104 39664 28888 39686
rect 26513 39491 26571 39497
rect 26513 39457 26525 39491
rect 26559 39488 26571 39491
rect 27890 39488 27896 39500
rect 26559 39460 27896 39488
rect 26559 39457 26571 39460
rect 26513 39451 26571 39457
rect 27890 39448 27896 39460
rect 27948 39448 27954 39500
rect 28353 39491 28411 39497
rect 28353 39457 28365 39491
rect 28399 39488 28411 39491
rect 29914 39488 29920 39500
rect 28399 39460 29920 39488
rect 28399 39457 28411 39460
rect 28353 39451 28411 39457
rect 29914 39448 29920 39460
rect 29972 39448 29978 39500
rect 1949 39423 2007 39429
rect 1949 39389 1961 39423
rect 1995 39389 2007 39423
rect 1949 39383 2007 39389
rect 2593 39423 2651 39429
rect 2593 39389 2605 39423
rect 2639 39420 2651 39423
rect 2774 39420 2780 39432
rect 2639 39392 2780 39420
rect 2639 39389 2651 39392
rect 2593 39383 2651 39389
rect 1964 39352 1992 39383
rect 2774 39380 2780 39392
rect 2832 39380 2838 39432
rect 3234 39420 3240 39432
rect 3147 39392 3240 39420
rect 3234 39380 3240 39392
rect 3292 39420 3298 39432
rect 3292 39392 6914 39420
rect 3292 39380 3298 39392
rect 4338 39352 4344 39364
rect 1964 39324 4344 39352
rect 4338 39312 4344 39324
rect 4396 39312 4402 39364
rect 1762 39244 1768 39296
rect 1820 39284 1826 39296
rect 1857 39287 1915 39293
rect 1857 39284 1869 39287
rect 1820 39256 1869 39284
rect 1820 39244 1826 39256
rect 1857 39253 1869 39256
rect 1903 39253 1915 39287
rect 1857 39247 1915 39253
rect 2958 39244 2964 39296
rect 3016 39284 3022 39296
rect 3145 39287 3203 39293
rect 3145 39284 3157 39287
rect 3016 39256 3157 39284
rect 3016 39244 3022 39256
rect 3145 39253 3157 39256
rect 3191 39253 3203 39287
rect 6886 39284 6914 39392
rect 26418 39312 26424 39364
rect 26476 39352 26482 39364
rect 26697 39355 26755 39361
rect 26697 39352 26709 39355
rect 26476 39324 26709 39352
rect 26476 39312 26482 39324
rect 26697 39321 26709 39324
rect 26743 39321 26755 39355
rect 26697 39315 26755 39321
rect 26326 39284 26332 39296
rect 6886 39256 26332 39284
rect 3145 39247 3203 39253
rect 26326 39244 26332 39256
rect 26384 39244 26390 39296
rect 1104 39194 29048 39216
rect 1104 39142 7896 39194
rect 7948 39142 7960 39194
rect 8012 39142 8024 39194
rect 8076 39142 8088 39194
rect 8140 39142 8152 39194
rect 8204 39142 14842 39194
rect 14894 39142 14906 39194
rect 14958 39142 14970 39194
rect 15022 39142 15034 39194
rect 15086 39142 15098 39194
rect 15150 39142 21788 39194
rect 21840 39142 21852 39194
rect 21904 39142 21916 39194
rect 21968 39142 21980 39194
rect 22032 39142 22044 39194
rect 22096 39142 28734 39194
rect 28786 39142 28798 39194
rect 28850 39142 28862 39194
rect 28914 39142 28926 39194
rect 28978 39142 28990 39194
rect 29042 39142 29048 39194
rect 1104 39120 29048 39142
rect 19981 39083 20039 39089
rect 19981 39049 19993 39083
rect 20027 39080 20039 39083
rect 26513 39083 26571 39089
rect 20027 39052 21036 39080
rect 20027 39049 20039 39052
rect 19981 39043 20039 39049
rect 2958 39012 2964 39024
rect 2919 38984 2964 39012
rect 2958 38972 2964 38984
rect 3016 38972 3022 39024
rect 1765 38947 1823 38953
rect 1765 38913 1777 38947
rect 1811 38944 1823 38947
rect 2774 38944 2780 38956
rect 1811 38916 2636 38944
rect 2735 38916 2780 38944
rect 1811 38913 1823 38916
rect 1765 38907 1823 38913
rect 2608 38876 2636 38916
rect 2774 38904 2780 38916
rect 2832 38904 2838 38956
rect 18966 38944 18972 38956
rect 18927 38916 18972 38944
rect 18966 38904 18972 38916
rect 19024 38904 19030 38956
rect 19797 38947 19855 38953
rect 19797 38913 19809 38947
rect 19843 38913 19855 38947
rect 20070 38944 20076 38956
rect 20031 38916 20076 38944
rect 19797 38907 19855 38913
rect 4246 38876 4252 38888
rect 2608 38848 2912 38876
rect 4207 38848 4252 38876
rect 2884 38820 2912 38848
rect 4246 38836 4252 38848
rect 4304 38836 4310 38888
rect 19812 38876 19840 38907
rect 20070 38904 20076 38916
rect 20128 38904 20134 38956
rect 20714 38944 20720 38956
rect 20675 38916 20720 38944
rect 20714 38904 20720 38916
rect 20772 38904 20778 38956
rect 21008 38944 21036 39052
rect 26513 39049 26525 39083
rect 26559 39080 26571 39083
rect 26694 39080 26700 39092
rect 26559 39052 26700 39080
rect 26559 39049 26571 39052
rect 26513 39043 26571 39049
rect 26694 39040 26700 39052
rect 26752 39040 26758 39092
rect 21177 38947 21235 38953
rect 21177 38944 21189 38947
rect 21008 38916 21189 38944
rect 21177 38913 21189 38916
rect 21223 38913 21235 38947
rect 21177 38907 21235 38913
rect 21361 38947 21419 38953
rect 21361 38913 21373 38947
rect 21407 38944 21419 38947
rect 21407 38916 21772 38944
rect 21407 38913 21419 38916
rect 21361 38907 21419 38913
rect 20530 38876 20536 38888
rect 19812 38848 20536 38876
rect 20530 38836 20536 38848
rect 20588 38836 20594 38888
rect 21192 38876 21220 38907
rect 21634 38876 21640 38888
rect 21192 38848 21640 38876
rect 21634 38836 21640 38848
rect 21692 38836 21698 38888
rect 2866 38768 2872 38820
rect 2924 38768 2930 38820
rect 19153 38811 19211 38817
rect 19153 38777 19165 38811
rect 19199 38808 19211 38811
rect 19702 38808 19708 38820
rect 19199 38780 19708 38808
rect 19199 38777 19211 38780
rect 19153 38771 19211 38777
rect 19702 38768 19708 38780
rect 19760 38768 19766 38820
rect 20070 38768 20076 38820
rect 20128 38808 20134 38820
rect 21744 38808 21772 38916
rect 26326 38904 26332 38956
rect 26384 38944 26390 38956
rect 26421 38947 26479 38953
rect 26421 38944 26433 38947
rect 26384 38916 26433 38944
rect 26384 38904 26390 38916
rect 26421 38913 26433 38916
rect 26467 38944 26479 38947
rect 27338 38944 27344 38956
rect 26467 38916 27344 38944
rect 26467 38913 26479 38916
rect 26421 38907 26479 38913
rect 27338 38904 27344 38916
rect 27396 38904 27402 38956
rect 21818 38808 21824 38820
rect 20128 38780 21824 38808
rect 20128 38768 20134 38780
rect 21818 38768 21824 38780
rect 21876 38768 21882 38820
rect 26510 38768 26516 38820
rect 26568 38808 26574 38820
rect 27801 38811 27859 38817
rect 27801 38808 27813 38811
rect 26568 38780 27813 38808
rect 26568 38768 26574 38780
rect 27801 38777 27813 38780
rect 27847 38777 27859 38811
rect 27801 38771 27859 38777
rect 1578 38740 1584 38752
rect 1539 38712 1584 38740
rect 1578 38700 1584 38712
rect 1636 38700 1642 38752
rect 19610 38740 19616 38752
rect 19571 38712 19616 38740
rect 19610 38700 19616 38712
rect 19668 38700 19674 38752
rect 20346 38700 20352 38752
rect 20404 38740 20410 38752
rect 20533 38743 20591 38749
rect 20533 38740 20545 38743
rect 20404 38712 20545 38740
rect 20404 38700 20410 38712
rect 20533 38709 20545 38712
rect 20579 38709 20591 38743
rect 21266 38740 21272 38752
rect 21227 38712 21272 38740
rect 20533 38703 20591 38709
rect 21266 38700 21272 38712
rect 21324 38700 21330 38752
rect 26694 38700 26700 38752
rect 26752 38740 26758 38752
rect 27249 38743 27307 38749
rect 27249 38740 27261 38743
rect 26752 38712 27261 38740
rect 26752 38700 26758 38712
rect 27249 38709 27261 38712
rect 27295 38709 27307 38743
rect 27249 38703 27307 38709
rect 1104 38650 28888 38672
rect 1104 38598 4423 38650
rect 4475 38598 4487 38650
rect 4539 38598 4551 38650
rect 4603 38598 4615 38650
rect 4667 38598 4679 38650
rect 4731 38598 11369 38650
rect 11421 38598 11433 38650
rect 11485 38598 11497 38650
rect 11549 38598 11561 38650
rect 11613 38598 11625 38650
rect 11677 38598 18315 38650
rect 18367 38598 18379 38650
rect 18431 38598 18443 38650
rect 18495 38598 18507 38650
rect 18559 38598 18571 38650
rect 18623 38598 25261 38650
rect 25313 38598 25325 38650
rect 25377 38598 25389 38650
rect 25441 38598 25453 38650
rect 25505 38598 25517 38650
rect 25569 38598 28888 38650
rect 1104 38576 28888 38598
rect 18690 38536 18696 38548
rect 18651 38508 18696 38536
rect 18690 38496 18696 38508
rect 18748 38496 18754 38548
rect 18877 38539 18935 38545
rect 18877 38505 18889 38539
rect 18923 38536 18935 38539
rect 18966 38536 18972 38548
rect 18923 38508 18972 38536
rect 18923 38505 18935 38508
rect 18877 38499 18935 38505
rect 18966 38496 18972 38508
rect 19024 38496 19030 38548
rect 20349 38539 20407 38545
rect 20349 38536 20361 38539
rect 19076 38508 20361 38536
rect 1670 38468 1676 38480
rect 1596 38440 1676 38468
rect 1596 38409 1624 38440
rect 1670 38428 1676 38440
rect 1728 38428 1734 38480
rect 19076 38468 19104 38508
rect 18524 38440 19104 38468
rect 1581 38403 1639 38409
rect 1581 38369 1593 38403
rect 1627 38369 1639 38403
rect 1762 38400 1768 38412
rect 1723 38372 1768 38400
rect 1581 38363 1639 38369
rect 1762 38360 1768 38372
rect 1820 38360 1826 38412
rect 2774 38400 2780 38412
rect 2735 38372 2780 38400
rect 2774 38360 2780 38372
rect 2832 38360 2838 38412
rect 18046 38224 18052 38276
rect 18104 38264 18110 38276
rect 18524 38273 18552 38440
rect 18509 38267 18567 38273
rect 18509 38264 18521 38267
rect 18104 38236 18521 38264
rect 18104 38224 18110 38236
rect 18509 38233 18521 38236
rect 18555 38233 18567 38267
rect 18509 38227 18567 38233
rect 18725 38267 18783 38273
rect 18725 38233 18737 38267
rect 18771 38264 18783 38267
rect 19610 38264 19616 38276
rect 18771 38236 19616 38264
rect 18771 38233 18783 38236
rect 18725 38227 18783 38233
rect 19610 38224 19616 38236
rect 19668 38224 19674 38276
rect 19904 38264 19932 38508
rect 20349 38505 20361 38508
rect 20395 38505 20407 38539
rect 20349 38499 20407 38505
rect 20533 38539 20591 38545
rect 20533 38505 20545 38539
rect 20579 38536 20591 38539
rect 20714 38536 20720 38548
rect 20579 38508 20720 38536
rect 20579 38505 20591 38508
rect 20533 38499 20591 38505
rect 20714 38496 20720 38508
rect 20772 38496 20778 38548
rect 21177 38539 21235 38545
rect 21177 38505 21189 38539
rect 21223 38536 21235 38539
rect 22189 38539 22247 38545
rect 22189 38536 22201 38539
rect 21223 38508 22201 38536
rect 21223 38505 21235 38508
rect 21177 38499 21235 38505
rect 22189 38505 22201 38508
rect 22235 38505 22247 38539
rect 22189 38499 22247 38505
rect 25961 38539 26019 38545
rect 25961 38505 25973 38539
rect 26007 38536 26019 38539
rect 26418 38536 26424 38548
rect 26007 38508 26424 38536
rect 26007 38505 26019 38508
rect 25961 38499 26019 38505
rect 26418 38496 26424 38508
rect 26476 38496 26482 38548
rect 19981 38471 20039 38477
rect 19981 38437 19993 38471
rect 20027 38468 20039 38471
rect 20070 38468 20076 38480
rect 20027 38440 20076 38468
rect 20027 38437 20039 38440
rect 19981 38431 20039 38437
rect 20070 38428 20076 38440
rect 20128 38428 20134 38480
rect 26510 38400 26516 38412
rect 26471 38372 26516 38400
rect 26510 38360 26516 38372
rect 26568 38360 26574 38412
rect 26694 38400 26700 38412
rect 26655 38372 26700 38400
rect 26694 38360 26700 38372
rect 26752 38360 26758 38412
rect 28353 38403 28411 38409
rect 28353 38369 28365 38403
rect 28399 38400 28411 38403
rect 28626 38400 28632 38412
rect 28399 38372 28632 38400
rect 28399 38369 28411 38372
rect 28353 38363 28411 38369
rect 28626 38360 28632 38372
rect 28684 38360 28690 38412
rect 21818 38332 21824 38344
rect 21779 38304 21824 38332
rect 21818 38292 21824 38304
rect 21876 38292 21882 38344
rect 25869 38335 25927 38341
rect 25869 38301 25881 38335
rect 25915 38332 25927 38335
rect 25915 38304 26234 38332
rect 25915 38301 25927 38304
rect 25869 38295 25927 38301
rect 21266 38273 21272 38276
rect 20993 38267 21051 38273
rect 20993 38264 21005 38267
rect 19904 38236 21005 38264
rect 20993 38233 21005 38236
rect 21039 38233 21051 38267
rect 20993 38227 21051 38233
rect 21209 38267 21272 38273
rect 21209 38233 21221 38267
rect 21255 38233 21272 38267
rect 21209 38227 21272 38233
rect 21266 38224 21272 38227
rect 21324 38224 21330 38276
rect 21634 38224 21640 38276
rect 21692 38264 21698 38276
rect 22005 38267 22063 38273
rect 22005 38264 22017 38267
rect 21692 38236 22017 38264
rect 21692 38224 21698 38236
rect 22005 38233 22017 38236
rect 22051 38233 22063 38267
rect 26206 38264 26234 38304
rect 26878 38264 26884 38276
rect 26206 38236 26884 38264
rect 22005 38227 22063 38233
rect 26878 38224 26884 38236
rect 26936 38224 26942 38276
rect 20349 38199 20407 38205
rect 20349 38165 20361 38199
rect 20395 38196 20407 38199
rect 20438 38196 20444 38208
rect 20395 38168 20444 38196
rect 20395 38165 20407 38168
rect 20349 38159 20407 38165
rect 20438 38156 20444 38168
rect 20496 38156 20502 38208
rect 21358 38196 21364 38208
rect 21319 38168 21364 38196
rect 21358 38156 21364 38168
rect 21416 38156 21422 38208
rect 1104 38106 29048 38128
rect 1104 38054 7896 38106
rect 7948 38054 7960 38106
rect 8012 38054 8024 38106
rect 8076 38054 8088 38106
rect 8140 38054 8152 38106
rect 8204 38054 14842 38106
rect 14894 38054 14906 38106
rect 14958 38054 14970 38106
rect 15022 38054 15034 38106
rect 15086 38054 15098 38106
rect 15150 38054 21788 38106
rect 21840 38054 21852 38106
rect 21904 38054 21916 38106
rect 21968 38054 21980 38106
rect 22032 38054 22044 38106
rect 22096 38054 28734 38106
rect 28786 38054 28798 38106
rect 28850 38054 28862 38106
rect 28914 38054 28926 38106
rect 28978 38054 28990 38106
rect 29042 38054 29048 38106
rect 1104 38032 29048 38054
rect 20349 37995 20407 38001
rect 20349 37961 20361 37995
rect 20395 37992 20407 37995
rect 20714 37992 20720 38004
rect 20395 37964 20720 37992
rect 20395 37961 20407 37964
rect 20349 37955 20407 37961
rect 20714 37952 20720 37964
rect 20772 37952 20778 38004
rect 20806 37952 20812 38004
rect 20864 37992 20870 38004
rect 20864 37964 21496 37992
rect 20864 37952 20870 37964
rect 19610 37924 19616 37936
rect 18432 37896 19616 37924
rect 18432 37865 18460 37896
rect 19610 37884 19616 37896
rect 19668 37884 19674 37936
rect 20257 37927 20315 37933
rect 20257 37893 20269 37927
rect 20303 37924 20315 37927
rect 20990 37924 20996 37936
rect 20303 37896 20996 37924
rect 20303 37893 20315 37896
rect 20257 37887 20315 37893
rect 20990 37884 20996 37896
rect 21048 37924 21054 37936
rect 21468 37933 21496 37964
rect 21237 37927 21295 37933
rect 21237 37924 21249 37927
rect 21048 37896 21249 37924
rect 21048 37884 21054 37896
rect 21237 37893 21249 37896
rect 21283 37893 21295 37927
rect 21237 37887 21295 37893
rect 21453 37927 21511 37933
rect 21453 37893 21465 37927
rect 21499 37893 21511 37927
rect 21453 37887 21511 37893
rect 18417 37859 18475 37865
rect 18417 37825 18429 37859
rect 18463 37825 18475 37859
rect 18417 37819 18475 37825
rect 18601 37859 18659 37865
rect 18601 37825 18613 37859
rect 18647 37856 18659 37859
rect 18690 37856 18696 37868
rect 18647 37828 18696 37856
rect 18647 37825 18659 37828
rect 18601 37819 18659 37825
rect 1670 37788 1676 37800
rect 1631 37760 1676 37788
rect 1670 37748 1676 37760
rect 1728 37748 1734 37800
rect 2774 37748 2780 37800
rect 2832 37788 2838 37800
rect 3329 37791 3387 37797
rect 3329 37788 3341 37791
rect 2832 37760 3341 37788
rect 2832 37748 2838 37760
rect 3329 37757 3341 37760
rect 3375 37757 3387 37791
rect 3329 37751 3387 37757
rect 3513 37791 3571 37797
rect 3513 37757 3525 37791
rect 3559 37788 3571 37791
rect 3973 37791 4031 37797
rect 3973 37788 3985 37791
rect 3559 37760 3985 37788
rect 3559 37757 3571 37760
rect 3513 37751 3571 37757
rect 3973 37757 3985 37760
rect 4019 37757 4031 37791
rect 18616 37788 18644 37819
rect 18690 37816 18696 37828
rect 18748 37816 18754 37868
rect 19058 37856 19064 37868
rect 19019 37828 19064 37856
rect 19058 37816 19064 37828
rect 19116 37816 19122 37868
rect 19245 37859 19303 37865
rect 19245 37825 19257 37859
rect 19291 37856 19303 37859
rect 19978 37856 19984 37868
rect 19291 37828 19984 37856
rect 19291 37825 19303 37828
rect 19245 37819 19303 37825
rect 19978 37816 19984 37828
rect 20036 37856 20042 37868
rect 20073 37859 20131 37865
rect 20073 37856 20085 37859
rect 20036 37828 20085 37856
rect 20036 37816 20042 37828
rect 20073 37825 20085 37828
rect 20119 37825 20131 37859
rect 20073 37819 20131 37825
rect 20441 37859 20499 37865
rect 20441 37825 20453 37859
rect 20487 37825 20499 37859
rect 20441 37819 20499 37825
rect 19153 37791 19211 37797
rect 19153 37788 19165 37791
rect 18616 37760 19165 37788
rect 3973 37751 4031 37757
rect 19153 37757 19165 37760
rect 19199 37757 19211 37791
rect 20456 37788 20484 37819
rect 21358 37816 21364 37868
rect 21416 37856 21422 37868
rect 22005 37859 22063 37865
rect 22005 37856 22017 37859
rect 21416 37828 22017 37856
rect 21416 37816 21422 37828
rect 22005 37825 22017 37828
rect 22051 37825 22063 37859
rect 27338 37856 27344 37868
rect 27251 37828 27344 37856
rect 22005 37819 22063 37825
rect 27338 37816 27344 37828
rect 27396 37856 27402 37868
rect 27982 37856 27988 37868
rect 27396 37828 27988 37856
rect 27396 37816 27402 37828
rect 27982 37816 27988 37828
rect 28040 37816 28046 37868
rect 21634 37788 21640 37800
rect 20456 37760 21640 37788
rect 19153 37751 19211 37757
rect 21634 37748 21640 37760
rect 21692 37748 21698 37800
rect 27706 37788 27712 37800
rect 27667 37760 27712 37788
rect 27706 37748 27712 37760
rect 27764 37748 27770 37800
rect 20530 37680 20536 37732
rect 20588 37720 20594 37732
rect 20625 37723 20683 37729
rect 20625 37720 20637 37723
rect 20588 37692 20637 37720
rect 20588 37680 20594 37692
rect 20625 37689 20637 37692
rect 20671 37689 20683 37723
rect 20625 37683 20683 37689
rect 20714 37680 20720 37732
rect 20772 37720 20778 37732
rect 20772 37692 21312 37720
rect 20772 37680 20778 37692
rect 18230 37612 18236 37664
rect 18288 37652 18294 37664
rect 18509 37655 18567 37661
rect 18509 37652 18521 37655
rect 18288 37624 18521 37652
rect 18288 37612 18294 37624
rect 18509 37621 18521 37624
rect 18555 37621 18567 37655
rect 18509 37615 18567 37621
rect 20070 37612 20076 37664
rect 20128 37652 20134 37664
rect 21284 37661 21312 37692
rect 21085 37655 21143 37661
rect 21085 37652 21097 37655
rect 20128 37624 21097 37652
rect 20128 37612 20134 37624
rect 21085 37621 21097 37624
rect 21131 37621 21143 37655
rect 21085 37615 21143 37621
rect 21269 37655 21327 37661
rect 21269 37621 21281 37655
rect 21315 37621 21327 37655
rect 21269 37615 21327 37621
rect 22189 37655 22247 37661
rect 22189 37621 22201 37655
rect 22235 37652 22247 37655
rect 22370 37652 22376 37664
rect 22235 37624 22376 37652
rect 22235 37621 22247 37624
rect 22189 37615 22247 37621
rect 22370 37612 22376 37624
rect 22428 37612 22434 37664
rect 1104 37562 28888 37584
rect 1104 37510 4423 37562
rect 4475 37510 4487 37562
rect 4539 37510 4551 37562
rect 4603 37510 4615 37562
rect 4667 37510 4679 37562
rect 4731 37510 11369 37562
rect 11421 37510 11433 37562
rect 11485 37510 11497 37562
rect 11549 37510 11561 37562
rect 11613 37510 11625 37562
rect 11677 37510 18315 37562
rect 18367 37510 18379 37562
rect 18431 37510 18443 37562
rect 18495 37510 18507 37562
rect 18559 37510 18571 37562
rect 18623 37510 25261 37562
rect 25313 37510 25325 37562
rect 25377 37510 25389 37562
rect 25441 37510 25453 37562
rect 25505 37510 25517 37562
rect 25569 37510 28888 37562
rect 1104 37488 28888 37510
rect 18230 37448 18236 37460
rect 18191 37420 18236 37448
rect 18230 37408 18236 37420
rect 18288 37408 18294 37460
rect 19334 37408 19340 37460
rect 19392 37448 19398 37460
rect 19610 37448 19616 37460
rect 19392 37420 19616 37448
rect 19392 37408 19398 37420
rect 19610 37408 19616 37420
rect 19668 37408 19674 37460
rect 20438 37448 20444 37460
rect 20399 37420 20444 37448
rect 20438 37408 20444 37420
rect 20496 37408 20502 37460
rect 3068 37352 19012 37380
rect 3068 37321 3096 37352
rect 3053 37315 3111 37321
rect 3053 37312 3065 37315
rect 1780 37284 3065 37312
rect 1486 37204 1492 37256
rect 1544 37244 1550 37256
rect 1780 37253 1808 37284
rect 3053 37281 3065 37284
rect 3099 37281 3111 37315
rect 16850 37312 16856 37324
rect 16811 37284 16856 37312
rect 3053 37275 3111 37281
rect 16850 37272 16856 37284
rect 16908 37272 16914 37324
rect 18984 37312 19012 37352
rect 19058 37340 19064 37392
rect 19116 37380 19122 37392
rect 20806 37380 20812 37392
rect 19116 37352 20812 37380
rect 19116 37340 19122 37352
rect 20806 37340 20812 37352
rect 20864 37340 20870 37392
rect 19518 37312 19524 37324
rect 18984 37284 19524 37312
rect 19518 37272 19524 37284
rect 19576 37272 19582 37324
rect 19705 37315 19763 37321
rect 19705 37281 19717 37315
rect 19751 37312 19763 37315
rect 21358 37312 21364 37324
rect 19751 37284 21364 37312
rect 19751 37281 19763 37284
rect 19705 37275 19763 37281
rect 21358 37272 21364 37284
rect 21416 37272 21422 37324
rect 1765 37247 1823 37253
rect 1765 37244 1777 37247
rect 1544 37216 1777 37244
rect 1544 37204 1550 37216
rect 1765 37213 1777 37216
rect 1811 37213 1823 37247
rect 1765 37207 1823 37213
rect 1857 37247 1915 37253
rect 1857 37213 1869 37247
rect 1903 37244 1915 37247
rect 2774 37244 2780 37256
rect 1903 37216 2780 37244
rect 1903 37213 1915 37216
rect 1857 37207 1915 37213
rect 2774 37204 2780 37216
rect 2832 37204 2838 37256
rect 3237 37247 3295 37253
rect 3237 37213 3249 37247
rect 3283 37244 3295 37247
rect 4801 37247 4859 37253
rect 4801 37244 4813 37247
rect 3283 37216 4813 37244
rect 3283 37213 3295 37216
rect 3237 37207 3295 37213
rect 4801 37213 4813 37216
rect 4847 37213 4859 37247
rect 4801 37207 4859 37213
rect 2682 37136 2688 37188
rect 2740 37176 2746 37188
rect 3252 37176 3280 37207
rect 5994 37204 6000 37256
rect 6052 37244 6058 37256
rect 16945 37247 17003 37253
rect 16945 37244 16957 37247
rect 6052 37216 16957 37244
rect 6052 37204 6058 37216
rect 16945 37213 16957 37216
rect 16991 37213 17003 37247
rect 19978 37244 19984 37256
rect 16945 37207 17003 37213
rect 17052 37216 18276 37244
rect 19939 37216 19984 37244
rect 2740 37148 3280 37176
rect 4157 37179 4215 37185
rect 2740 37136 2746 37148
rect 4157 37145 4169 37179
rect 4203 37176 4215 37179
rect 4338 37176 4344 37188
rect 4203 37148 4344 37176
rect 4203 37145 4215 37148
rect 4157 37139 4215 37145
rect 4338 37136 4344 37148
rect 4396 37136 4402 37188
rect 15286 37136 15292 37188
rect 15344 37176 15350 37188
rect 17052 37176 17080 37216
rect 17954 37176 17960 37188
rect 15344 37148 17080 37176
rect 17236 37148 17960 37176
rect 15344 37136 15350 37148
rect 17037 37111 17095 37117
rect 17037 37077 17049 37111
rect 17083 37108 17095 37111
rect 17236 37108 17264 37148
rect 17954 37136 17960 37148
rect 18012 37136 18018 37188
rect 18046 37136 18052 37188
rect 18104 37176 18110 37188
rect 18248 37185 18276 37216
rect 19978 37204 19984 37216
rect 20036 37204 20042 37256
rect 20625 37247 20683 37253
rect 20625 37213 20637 37247
rect 20671 37244 20683 37247
rect 20714 37244 20720 37256
rect 20671 37216 20720 37244
rect 20671 37213 20683 37216
rect 20625 37207 20683 37213
rect 20714 37204 20720 37216
rect 20772 37204 20778 37256
rect 20901 37247 20959 37253
rect 20901 37213 20913 37247
rect 20947 37244 20959 37247
rect 20990 37244 20996 37256
rect 20947 37216 20996 37244
rect 20947 37213 20959 37216
rect 20901 37207 20959 37213
rect 20990 37204 20996 37216
rect 21048 37204 21054 37256
rect 28350 37204 28356 37256
rect 28408 37244 28414 37256
rect 28408 37216 28453 37244
rect 28408 37204 28414 37216
rect 18248 37179 18323 37185
rect 18104 37148 18149 37176
rect 18248 37148 18277 37179
rect 18104 37136 18110 37148
rect 18265 37145 18277 37148
rect 18311 37176 18323 37179
rect 18311 37148 19472 37176
rect 18311 37145 18323 37148
rect 18265 37139 18323 37145
rect 17402 37108 17408 37120
rect 17083 37080 17264 37108
rect 17363 37080 17408 37108
rect 17083 37077 17095 37080
rect 17037 37071 17095 37077
rect 17402 37068 17408 37080
rect 17460 37068 17466 37120
rect 18414 37108 18420 37120
rect 18375 37080 18420 37108
rect 18414 37068 18420 37080
rect 18472 37068 18478 37120
rect 19444 37117 19472 37148
rect 26142 37136 26148 37188
rect 26200 37176 26206 37188
rect 26513 37179 26571 37185
rect 26513 37176 26525 37179
rect 26200 37148 26525 37176
rect 26200 37136 26206 37148
rect 26513 37145 26525 37148
rect 26559 37145 26571 37179
rect 26513 37139 26571 37145
rect 27890 37136 27896 37188
rect 27948 37176 27954 37188
rect 28169 37179 28227 37185
rect 28169 37176 28181 37179
rect 27948 37148 28181 37176
rect 27948 37136 27954 37148
rect 28169 37145 28181 37148
rect 28215 37145 28227 37179
rect 28169 37139 28227 37145
rect 19429 37111 19487 37117
rect 19429 37077 19441 37111
rect 19475 37077 19487 37111
rect 20806 37108 20812 37120
rect 20767 37080 20812 37108
rect 19429 37071 19487 37077
rect 20806 37068 20812 37080
rect 20864 37068 20870 37120
rect 1104 37018 29048 37040
rect 1104 36966 7896 37018
rect 7948 36966 7960 37018
rect 8012 36966 8024 37018
rect 8076 36966 8088 37018
rect 8140 36966 8152 37018
rect 8204 36966 14842 37018
rect 14894 36966 14906 37018
rect 14958 36966 14970 37018
rect 15022 36966 15034 37018
rect 15086 36966 15098 37018
rect 15150 36966 21788 37018
rect 21840 36966 21852 37018
rect 21904 36966 21916 37018
rect 21968 36966 21980 37018
rect 22032 36966 22044 37018
rect 22096 36966 28734 37018
rect 28786 36966 28798 37018
rect 28850 36966 28862 37018
rect 28914 36966 28926 37018
rect 28978 36966 28990 37018
rect 29042 36966 29048 37018
rect 1104 36944 29048 36966
rect 15746 36864 15752 36916
rect 15804 36904 15810 36916
rect 18046 36904 18052 36916
rect 15804 36876 18052 36904
rect 15804 36864 15810 36876
rect 18046 36864 18052 36876
rect 18104 36864 18110 36916
rect 21358 36904 21364 36916
rect 21319 36876 21364 36904
rect 21358 36864 21364 36876
rect 21416 36864 21422 36916
rect 27890 36904 27896 36916
rect 27851 36876 27896 36904
rect 27890 36864 27896 36876
rect 27948 36864 27954 36916
rect 4338 36796 4344 36848
rect 4396 36836 4402 36848
rect 19426 36836 19432 36848
rect 4396 36808 19432 36836
rect 4396 36796 4402 36808
rect 19426 36796 19432 36808
rect 19484 36796 19490 36848
rect 26206 36808 26648 36836
rect 2590 36768 2596 36780
rect 2551 36740 2596 36768
rect 2590 36728 2596 36740
rect 2648 36768 2654 36780
rect 3237 36771 3295 36777
rect 3237 36768 3249 36771
rect 2648 36740 3249 36768
rect 2648 36728 2654 36740
rect 3237 36737 3249 36740
rect 3283 36768 3295 36771
rect 4709 36771 4767 36777
rect 4709 36768 4721 36771
rect 3283 36740 4721 36768
rect 3283 36737 3295 36740
rect 3237 36731 3295 36737
rect 4709 36737 4721 36740
rect 4755 36737 4767 36771
rect 4709 36731 4767 36737
rect 17037 36771 17095 36777
rect 17037 36737 17049 36771
rect 17083 36768 17095 36771
rect 17402 36768 17408 36780
rect 17083 36740 17408 36768
rect 17083 36737 17095 36740
rect 17037 36731 17095 36737
rect 17402 36728 17408 36740
rect 17460 36728 17466 36780
rect 18414 36768 18420 36780
rect 18375 36740 18420 36768
rect 18414 36728 18420 36740
rect 18472 36728 18478 36780
rect 21450 36768 21456 36780
rect 21411 36740 21456 36768
rect 21450 36728 21456 36740
rect 21508 36768 21514 36780
rect 22189 36771 22247 36777
rect 22189 36768 22201 36771
rect 21508 36740 22201 36768
rect 21508 36728 21514 36740
rect 22189 36737 22201 36740
rect 22235 36737 22247 36771
rect 22189 36731 22247 36737
rect 24854 36728 24860 36780
rect 24912 36768 24918 36780
rect 26206 36768 26234 36808
rect 26620 36777 26648 36808
rect 24912 36740 26234 36768
rect 26349 36771 26407 36777
rect 24912 36728 24918 36740
rect 26349 36737 26361 36771
rect 26395 36768 26407 36771
rect 26605 36771 26663 36777
rect 26395 36740 26556 36768
rect 26395 36737 26407 36740
rect 26349 36731 26407 36737
rect 2130 36660 2136 36712
rect 2188 36700 2194 36712
rect 2406 36700 2412 36712
rect 2188 36672 2412 36700
rect 2188 36660 2194 36672
rect 2406 36660 2412 36672
rect 2464 36660 2470 36712
rect 4065 36703 4123 36709
rect 4065 36669 4077 36703
rect 4111 36700 4123 36703
rect 4154 36700 4160 36712
rect 4111 36672 4160 36700
rect 4111 36669 4123 36672
rect 4065 36663 4123 36669
rect 4080 36564 4108 36663
rect 4154 36660 4160 36672
rect 4212 36660 4218 36712
rect 5537 36703 5595 36709
rect 5537 36669 5549 36703
rect 5583 36700 5595 36703
rect 9582 36700 9588 36712
rect 5583 36672 9588 36700
rect 5583 36669 5595 36672
rect 5537 36663 5595 36669
rect 9582 36660 9588 36672
rect 9640 36660 9646 36712
rect 16666 36660 16672 36712
rect 16724 36700 16730 36712
rect 16853 36703 16911 36709
rect 16853 36700 16865 36703
rect 16724 36672 16865 36700
rect 16724 36660 16730 36672
rect 16853 36669 16865 36672
rect 16899 36669 16911 36703
rect 26528 36700 26556 36740
rect 26605 36737 26617 36771
rect 26651 36737 26663 36771
rect 27338 36768 27344 36780
rect 27299 36740 27344 36768
rect 26605 36731 26663 36737
rect 27338 36728 27344 36740
rect 27396 36728 27402 36780
rect 27798 36768 27804 36780
rect 27759 36740 27804 36768
rect 27798 36728 27804 36740
rect 27856 36728 27862 36780
rect 26528 36672 27200 36700
rect 16853 36663 16911 36669
rect 27172 36641 27200 36672
rect 27157 36635 27215 36641
rect 27157 36601 27169 36635
rect 27203 36601 27215 36635
rect 27157 36595 27215 36601
rect 10686 36564 10692 36576
rect 4080 36536 10692 36564
rect 10686 36524 10692 36536
rect 10744 36524 10750 36576
rect 17221 36567 17279 36573
rect 17221 36533 17233 36567
rect 17267 36564 17279 36567
rect 17770 36564 17776 36576
rect 17267 36536 17776 36564
rect 17267 36533 17279 36536
rect 17221 36527 17279 36533
rect 17770 36524 17776 36536
rect 17828 36524 17834 36576
rect 18601 36567 18659 36573
rect 18601 36533 18613 36567
rect 18647 36564 18659 36567
rect 18782 36564 18788 36576
rect 18647 36536 18788 36564
rect 18647 36533 18659 36536
rect 18601 36527 18659 36533
rect 18782 36524 18788 36536
rect 18840 36524 18846 36576
rect 20806 36524 20812 36576
rect 20864 36564 20870 36576
rect 22465 36567 22523 36573
rect 22465 36564 22477 36567
rect 20864 36536 22477 36564
rect 20864 36524 20870 36536
rect 22465 36533 22477 36536
rect 22511 36564 22523 36567
rect 24670 36564 24676 36576
rect 22511 36536 24676 36564
rect 22511 36533 22523 36536
rect 22465 36527 22523 36533
rect 24670 36524 24676 36536
rect 24728 36524 24734 36576
rect 24762 36524 24768 36576
rect 24820 36564 24826 36576
rect 25225 36567 25283 36573
rect 25225 36564 25237 36567
rect 24820 36536 25237 36564
rect 24820 36524 24826 36536
rect 25225 36533 25237 36536
rect 25271 36533 25283 36567
rect 25225 36527 25283 36533
rect 1104 36474 28888 36496
rect 1104 36422 4423 36474
rect 4475 36422 4487 36474
rect 4539 36422 4551 36474
rect 4603 36422 4615 36474
rect 4667 36422 4679 36474
rect 4731 36422 11369 36474
rect 11421 36422 11433 36474
rect 11485 36422 11497 36474
rect 11549 36422 11561 36474
rect 11613 36422 11625 36474
rect 11677 36422 18315 36474
rect 18367 36422 18379 36474
rect 18431 36422 18443 36474
rect 18495 36422 18507 36474
rect 18559 36422 18571 36474
rect 18623 36422 25261 36474
rect 25313 36422 25325 36474
rect 25377 36422 25389 36474
rect 25441 36422 25453 36474
rect 25505 36422 25517 36474
rect 25569 36422 28888 36474
rect 1104 36400 28888 36422
rect 20714 36320 20720 36372
rect 20772 36360 20778 36372
rect 21453 36363 21511 36369
rect 21453 36360 21465 36363
rect 20772 36332 21465 36360
rect 20772 36320 20778 36332
rect 21453 36329 21465 36332
rect 21499 36329 21511 36363
rect 21453 36323 21511 36329
rect 28261 36363 28319 36369
rect 28261 36329 28273 36363
rect 28307 36360 28319 36363
rect 28350 36360 28356 36372
rect 28307 36332 28356 36360
rect 28307 36329 28319 36332
rect 28261 36323 28319 36329
rect 28350 36320 28356 36332
rect 28408 36320 28414 36372
rect 1949 36227 2007 36233
rect 1949 36193 1961 36227
rect 1995 36224 2007 36227
rect 3510 36224 3516 36236
rect 1995 36196 3516 36224
rect 1995 36193 2007 36196
rect 1949 36187 2007 36193
rect 3510 36184 3516 36196
rect 3568 36184 3574 36236
rect 4246 36184 4252 36236
rect 4304 36224 4310 36236
rect 4798 36224 4804 36236
rect 4304 36196 4804 36224
rect 4304 36184 4310 36196
rect 4798 36184 4804 36196
rect 4856 36184 4862 36236
rect 15654 36184 15660 36236
rect 15712 36224 15718 36236
rect 15841 36227 15899 36233
rect 15841 36224 15853 36227
rect 15712 36196 15853 36224
rect 15712 36184 15718 36196
rect 15841 36193 15853 36196
rect 15887 36224 15899 36227
rect 16850 36224 16856 36236
rect 15887 36196 16856 36224
rect 15887 36193 15899 36196
rect 15841 36187 15899 36193
rect 16850 36184 16856 36196
rect 16908 36224 16914 36236
rect 23566 36224 23572 36236
rect 16908 36196 20208 36224
rect 23527 36196 23572 36224
rect 16908 36184 16914 36196
rect 2406 36156 2412 36168
rect 2367 36128 2412 36156
rect 2406 36116 2412 36128
rect 2464 36156 2470 36168
rect 2590 36156 2596 36168
rect 2464 36128 2596 36156
rect 2464 36116 2470 36128
rect 2590 36116 2596 36128
rect 2648 36156 2654 36168
rect 3970 36156 3976 36168
rect 2648 36128 3976 36156
rect 2648 36116 2654 36128
rect 3970 36116 3976 36128
rect 4028 36156 4034 36168
rect 5537 36159 5595 36165
rect 5537 36156 5549 36159
rect 4028 36128 5549 36156
rect 4028 36116 4034 36128
rect 5537 36125 5549 36128
rect 5583 36125 5595 36159
rect 5537 36119 5595 36125
rect 16574 36116 16580 36168
rect 16632 36156 16638 36168
rect 16945 36159 17003 36165
rect 16945 36156 16957 36159
rect 16632 36128 16957 36156
rect 16632 36116 16638 36128
rect 16945 36125 16957 36128
rect 16991 36125 17003 36159
rect 17770 36156 17776 36168
rect 17731 36128 17776 36156
rect 16945 36119 17003 36125
rect 17770 36116 17776 36128
rect 17828 36116 17834 36168
rect 20070 36156 20076 36168
rect 20031 36128 20076 36156
rect 20070 36116 20076 36128
rect 20128 36116 20134 36168
rect 2958 36048 2964 36100
rect 3016 36088 3022 36100
rect 3234 36088 3240 36100
rect 3016 36060 3240 36088
rect 3016 36048 3022 36060
rect 3234 36048 3240 36060
rect 3292 36048 3298 36100
rect 5902 36088 5908 36100
rect 5863 36060 5908 36088
rect 5902 36048 5908 36060
rect 5960 36048 5966 36100
rect 9582 36048 9588 36100
rect 9640 36088 9646 36100
rect 9766 36088 9772 36100
rect 9640 36060 9772 36088
rect 9640 36048 9646 36060
rect 9766 36048 9772 36060
rect 9824 36088 9830 36100
rect 14458 36088 14464 36100
rect 9824 36060 14464 36088
rect 9824 36048 9830 36060
rect 14458 36048 14464 36060
rect 14516 36048 14522 36100
rect 16117 36091 16175 36097
rect 16117 36057 16129 36091
rect 16163 36088 16175 36091
rect 18230 36088 18236 36100
rect 16163 36060 18236 36088
rect 16163 36057 16175 36060
rect 16117 36051 16175 36057
rect 18230 36048 18236 36060
rect 18288 36048 18294 36100
rect 20180 36088 20208 36196
rect 23566 36184 23572 36196
rect 23624 36184 23630 36236
rect 23753 36227 23811 36233
rect 23753 36193 23765 36227
rect 23799 36224 23811 36227
rect 24486 36224 24492 36236
rect 23799 36196 24492 36224
rect 23799 36193 23811 36196
rect 23753 36187 23811 36193
rect 20346 36165 20352 36168
rect 20340 36156 20352 36165
rect 20307 36128 20352 36156
rect 20340 36119 20352 36128
rect 20346 36116 20352 36119
rect 20404 36116 20410 36168
rect 22649 36159 22707 36165
rect 22649 36125 22661 36159
rect 22695 36156 22707 36159
rect 23474 36156 23480 36168
rect 22695 36128 23480 36156
rect 22695 36125 22707 36128
rect 22649 36119 22707 36125
rect 23474 36116 23480 36128
rect 23532 36116 23538 36168
rect 23768 36088 23796 36187
rect 24486 36184 24492 36196
rect 24544 36184 24550 36236
rect 24762 36224 24768 36236
rect 24723 36196 24768 36224
rect 24762 36184 24768 36196
rect 24820 36184 24826 36236
rect 27430 36224 27436 36236
rect 27391 36196 27436 36224
rect 27430 36184 27436 36196
rect 27488 36184 27494 36236
rect 25774 36156 25780 36168
rect 25735 36128 25780 36156
rect 25774 36116 25780 36128
rect 25832 36116 25838 36168
rect 20180 36060 23796 36088
rect 25961 36091 26019 36097
rect 25961 36057 25973 36091
rect 26007 36088 26019 36091
rect 26234 36088 26240 36100
rect 26007 36060 26240 36088
rect 26007 36057 26019 36060
rect 25961 36051 26019 36057
rect 26234 36048 26240 36060
rect 26292 36048 26298 36100
rect 6730 35980 6736 36032
rect 6788 36020 6794 36032
rect 16025 36023 16083 36029
rect 16025 36020 16037 36023
rect 6788 35992 16037 36020
rect 6788 35980 6794 35992
rect 16025 35989 16037 35992
rect 16071 35989 16083 36023
rect 16482 36020 16488 36032
rect 16443 35992 16488 36020
rect 16025 35983 16083 35989
rect 16482 35980 16488 35992
rect 16540 35980 16546 36032
rect 17126 36020 17132 36032
rect 17087 35992 17132 36020
rect 17126 35980 17132 35992
rect 17184 35980 17190 36032
rect 17586 36020 17592 36032
rect 17547 35992 17592 36020
rect 17586 35980 17592 35992
rect 17644 35980 17650 36032
rect 18138 35980 18144 36032
rect 18196 36020 18202 36032
rect 19334 36020 19340 36032
rect 18196 35992 19340 36020
rect 18196 35980 18202 35992
rect 19334 35980 19340 35992
rect 19392 35980 19398 36032
rect 22465 36023 22523 36029
rect 22465 35989 22477 36023
rect 22511 36020 22523 36023
rect 22646 36020 22652 36032
rect 22511 35992 22652 36020
rect 22511 35989 22523 35992
rect 22465 35983 22523 35989
rect 22646 35980 22652 35992
rect 22704 35980 22710 36032
rect 23106 36020 23112 36032
rect 23067 35992 23112 36020
rect 23106 35980 23112 35992
rect 23164 35980 23170 36032
rect 23477 36023 23535 36029
rect 23477 35989 23489 36023
rect 23523 36020 23535 36023
rect 23750 36020 23756 36032
rect 23523 35992 23756 36020
rect 23523 35989 23535 35992
rect 23477 35983 23535 35989
rect 23750 35980 23756 35992
rect 23808 35980 23814 36032
rect 25317 36023 25375 36029
rect 25317 35989 25329 36023
rect 25363 36020 25375 36023
rect 25682 36020 25688 36032
rect 25363 35992 25688 36020
rect 25363 35989 25375 35992
rect 25317 35983 25375 35989
rect 25682 35980 25688 35992
rect 25740 35980 25746 36032
rect 1104 35930 29048 35952
rect 1104 35878 7896 35930
rect 7948 35878 7960 35930
rect 8012 35878 8024 35930
rect 8076 35878 8088 35930
rect 8140 35878 8152 35930
rect 8204 35878 14842 35930
rect 14894 35878 14906 35930
rect 14958 35878 14970 35930
rect 15022 35878 15034 35930
rect 15086 35878 15098 35930
rect 15150 35878 21788 35930
rect 21840 35878 21852 35930
rect 21904 35878 21916 35930
rect 21968 35878 21980 35930
rect 22032 35878 22044 35930
rect 22096 35878 28734 35930
rect 28786 35878 28798 35930
rect 28850 35878 28862 35930
rect 28914 35878 28926 35930
rect 28978 35878 28990 35930
rect 29042 35878 29048 35930
rect 1104 35856 29048 35878
rect 6886 35788 24992 35816
rect 1670 35748 1676 35760
rect 1631 35720 1676 35748
rect 1670 35708 1676 35720
rect 1728 35708 1734 35760
rect 5902 35708 5908 35760
rect 5960 35748 5966 35760
rect 6886 35748 6914 35788
rect 5960 35720 6914 35748
rect 16301 35751 16359 35757
rect 5960 35708 5966 35720
rect 16301 35717 16313 35751
rect 16347 35748 16359 35751
rect 16574 35748 16580 35760
rect 16347 35720 16580 35748
rect 16347 35717 16359 35720
rect 16301 35711 16359 35717
rect 16574 35708 16580 35720
rect 16632 35708 16638 35760
rect 17126 35757 17132 35760
rect 17120 35748 17132 35757
rect 17087 35720 17132 35748
rect 17120 35711 17132 35720
rect 17126 35708 17132 35711
rect 17184 35708 17190 35760
rect 20070 35748 20076 35760
rect 18708 35720 20076 35748
rect 3510 35640 3516 35692
rect 3568 35680 3574 35692
rect 3970 35680 3976 35692
rect 3568 35652 3613 35680
rect 3931 35652 3976 35680
rect 3568 35640 3574 35652
rect 3970 35640 3976 35652
rect 4028 35640 4034 35692
rect 7742 35680 7748 35692
rect 4356 35652 7748 35680
rect 4356 35624 4384 35652
rect 7742 35640 7748 35652
rect 7800 35640 7806 35692
rect 16117 35683 16175 35689
rect 16117 35649 16129 35683
rect 16163 35680 16175 35683
rect 16482 35680 16488 35692
rect 16163 35652 16488 35680
rect 16163 35649 16175 35652
rect 16117 35643 16175 35649
rect 16482 35640 16488 35652
rect 16540 35640 16546 35692
rect 18708 35689 18736 35720
rect 20070 35708 20076 35720
rect 20128 35708 20134 35760
rect 24854 35748 24860 35760
rect 22480 35720 24860 35748
rect 22480 35692 22508 35720
rect 18693 35683 18751 35689
rect 18693 35649 18705 35683
rect 18739 35649 18751 35683
rect 18693 35643 18751 35649
rect 18782 35640 18788 35692
rect 18840 35680 18846 35692
rect 18949 35683 19007 35689
rect 18949 35680 18961 35683
rect 18840 35652 18961 35680
rect 18840 35640 18846 35652
rect 18949 35649 18961 35652
rect 18995 35649 19007 35683
rect 18949 35643 19007 35649
rect 22373 35683 22431 35689
rect 22373 35649 22385 35683
rect 22419 35680 22431 35683
rect 22462 35680 22468 35692
rect 22419 35652 22468 35680
rect 22419 35649 22431 35652
rect 22373 35643 22431 35649
rect 22462 35640 22468 35652
rect 22520 35640 22526 35692
rect 22646 35689 22652 35692
rect 22640 35680 22652 35689
rect 22607 35652 22652 35680
rect 22640 35643 22652 35652
rect 22646 35640 22652 35643
rect 22704 35640 22710 35692
rect 24228 35689 24256 35720
rect 24854 35708 24860 35720
rect 24912 35708 24918 35760
rect 24213 35683 24271 35689
rect 24213 35649 24225 35683
rect 24259 35649 24271 35683
rect 24213 35643 24271 35649
rect 24480 35683 24538 35689
rect 24480 35649 24492 35683
rect 24526 35680 24538 35683
rect 24762 35680 24768 35692
rect 24526 35652 24768 35680
rect 24526 35649 24538 35652
rect 24480 35643 24538 35649
rect 24762 35640 24768 35652
rect 24820 35640 24826 35692
rect 24964 35680 24992 35788
rect 26234 35776 26240 35828
rect 26292 35816 26298 35828
rect 26292 35788 26337 35816
rect 26292 35776 26298 35788
rect 26329 35683 26387 35689
rect 26329 35680 26341 35683
rect 24964 35652 26341 35680
rect 26329 35649 26341 35652
rect 26375 35680 26387 35683
rect 26694 35680 26700 35692
rect 26375 35652 26700 35680
rect 26375 35649 26387 35652
rect 26329 35643 26387 35649
rect 26694 35640 26700 35652
rect 26752 35640 26758 35692
rect 3050 35572 3056 35624
rect 3108 35612 3114 35624
rect 3329 35615 3387 35621
rect 3329 35612 3341 35615
rect 3108 35584 3341 35612
rect 3108 35572 3114 35584
rect 3329 35581 3341 35584
rect 3375 35581 3387 35615
rect 4338 35612 4344 35624
rect 4299 35584 4344 35612
rect 3329 35575 3387 35581
rect 4338 35572 4344 35584
rect 4396 35572 4402 35624
rect 15933 35615 15991 35621
rect 15933 35581 15945 35615
rect 15979 35612 15991 35615
rect 16666 35612 16672 35624
rect 15979 35584 16672 35612
rect 15979 35581 15991 35584
rect 15933 35575 15991 35581
rect 16666 35572 16672 35584
rect 16724 35572 16730 35624
rect 16850 35612 16856 35624
rect 16811 35584 16856 35612
rect 16850 35572 16856 35584
rect 16908 35572 16914 35624
rect 18230 35544 18236 35556
rect 18191 35516 18236 35544
rect 18230 35504 18236 35516
rect 18288 35504 18294 35556
rect 19610 35436 19616 35488
rect 19668 35476 19674 35488
rect 20073 35479 20131 35485
rect 20073 35476 20085 35479
rect 19668 35448 20085 35476
rect 19668 35436 19674 35448
rect 20073 35445 20085 35448
rect 20119 35445 20131 35479
rect 23750 35476 23756 35488
rect 23711 35448 23756 35476
rect 20073 35439 20131 35445
rect 23750 35436 23756 35448
rect 23808 35436 23814 35488
rect 24118 35436 24124 35488
rect 24176 35476 24182 35488
rect 25593 35479 25651 35485
rect 25593 35476 25605 35479
rect 24176 35448 25605 35476
rect 24176 35436 24182 35448
rect 25593 35445 25605 35448
rect 25639 35476 25651 35479
rect 26234 35476 26240 35488
rect 25639 35448 26240 35476
rect 25639 35445 25651 35448
rect 25593 35439 25651 35445
rect 26234 35436 26240 35448
rect 26292 35436 26298 35488
rect 26510 35436 26516 35488
rect 26568 35476 26574 35488
rect 27157 35479 27215 35485
rect 27157 35476 27169 35479
rect 26568 35448 27169 35476
rect 26568 35436 26574 35448
rect 27157 35445 27169 35448
rect 27203 35445 27215 35479
rect 27157 35439 27215 35445
rect 1104 35386 28888 35408
rect 1104 35334 4423 35386
rect 4475 35334 4487 35386
rect 4539 35334 4551 35386
rect 4603 35334 4615 35386
rect 4667 35334 4679 35386
rect 4731 35334 11369 35386
rect 11421 35334 11433 35386
rect 11485 35334 11497 35386
rect 11549 35334 11561 35386
rect 11613 35334 11625 35386
rect 11677 35334 18315 35386
rect 18367 35334 18379 35386
rect 18431 35334 18443 35386
rect 18495 35334 18507 35386
rect 18559 35334 18571 35386
rect 18623 35334 25261 35386
rect 25313 35334 25325 35386
rect 25377 35334 25389 35386
rect 25441 35334 25453 35386
rect 25505 35334 25517 35386
rect 25569 35334 28888 35386
rect 1104 35312 28888 35334
rect 3050 35272 3056 35284
rect 3011 35244 3056 35272
rect 3050 35232 3056 35244
rect 3108 35232 3114 35284
rect 20530 35232 20536 35284
rect 20588 35272 20594 35284
rect 20809 35275 20867 35281
rect 20809 35272 20821 35275
rect 20588 35244 20821 35272
rect 20588 35232 20594 35244
rect 20809 35241 20821 35244
rect 20855 35241 20867 35275
rect 20809 35235 20867 35241
rect 21269 35275 21327 35281
rect 21269 35241 21281 35275
rect 21315 35272 21327 35275
rect 21634 35272 21640 35284
rect 21315 35244 21640 35272
rect 21315 35241 21327 35244
rect 21269 35235 21327 35241
rect 21634 35232 21640 35244
rect 21692 35232 21698 35284
rect 23474 35272 23480 35284
rect 23435 35244 23480 35272
rect 23474 35232 23480 35244
rect 23532 35232 23538 35284
rect 24762 35272 24768 35284
rect 24723 35244 24768 35272
rect 24762 35232 24768 35244
rect 24820 35232 24826 35284
rect 25409 35275 25467 35281
rect 25409 35241 25421 35275
rect 25455 35272 25467 35275
rect 25774 35272 25780 35284
rect 25455 35244 25780 35272
rect 25455 35241 25467 35244
rect 25409 35235 25467 35241
rect 25774 35232 25780 35244
rect 25832 35232 25838 35284
rect 2406 35136 2412 35148
rect 2367 35108 2412 35136
rect 2406 35096 2412 35108
rect 2464 35096 2470 35148
rect 25958 35136 25964 35148
rect 25884 35108 25964 35136
rect 1578 35068 1584 35080
rect 1539 35040 1584 35068
rect 1578 35028 1584 35040
rect 1636 35028 1642 35080
rect 2961 35071 3019 35077
rect 2961 35037 2973 35071
rect 3007 35068 3019 35071
rect 3878 35068 3884 35080
rect 3007 35040 3884 35068
rect 3007 35037 3019 35040
rect 2961 35031 3019 35037
rect 3878 35028 3884 35040
rect 3936 35068 3942 35080
rect 5902 35068 5908 35080
rect 3936 35040 5908 35068
rect 3936 35028 3942 35040
rect 5902 35028 5908 35040
rect 5960 35028 5966 35080
rect 16850 35068 16856 35080
rect 16763 35040 16856 35068
rect 16850 35028 16856 35040
rect 16908 35068 16914 35080
rect 19429 35071 19487 35077
rect 19429 35068 19441 35071
rect 16908 35040 19441 35068
rect 16908 35028 16914 35040
rect 19429 35037 19441 35040
rect 19475 35068 19487 35071
rect 20070 35068 20076 35080
rect 19475 35040 20076 35068
rect 19475 35037 19487 35040
rect 19429 35031 19487 35037
rect 20070 35028 20076 35040
rect 20128 35028 20134 35080
rect 22370 35068 22376 35080
rect 22428 35077 22434 35080
rect 22340 35040 22376 35068
rect 22370 35028 22376 35040
rect 22428 35031 22440 35077
rect 22428 35028 22434 35031
rect 22554 35028 22560 35080
rect 22612 35068 22618 35080
rect 22649 35071 22707 35077
rect 22649 35068 22661 35071
rect 22612 35040 22661 35068
rect 22612 35028 22618 35040
rect 22649 35037 22661 35040
rect 22695 35037 22707 35071
rect 23106 35068 23112 35080
rect 23067 35040 23112 35068
rect 22649 35031 22707 35037
rect 23106 35028 23112 35040
rect 23164 35028 23170 35080
rect 23293 35071 23351 35077
rect 23293 35037 23305 35071
rect 23339 35068 23351 35071
rect 24581 35071 24639 35077
rect 24581 35068 24593 35071
rect 23339 35040 24593 35068
rect 23339 35037 23351 35040
rect 23293 35031 23351 35037
rect 24581 35037 24593 35040
rect 24627 35037 24639 35071
rect 24581 35031 24639 35037
rect 24765 35071 24823 35077
rect 24765 35037 24777 35071
rect 24811 35037 24823 35071
rect 24765 35031 24823 35037
rect 17120 35003 17178 35009
rect 17120 34969 17132 35003
rect 17166 35000 17178 35003
rect 17586 35000 17592 35012
rect 17166 34972 17592 35000
rect 17166 34969 17178 34972
rect 17120 34963 17178 34969
rect 17586 34960 17592 34972
rect 17644 34960 17650 35012
rect 19702 35009 19708 35012
rect 19696 34963 19708 35009
rect 19760 35000 19766 35012
rect 19760 34972 19796 35000
rect 19702 34960 19708 34963
rect 19760 34960 19766 34972
rect 22738 34960 22744 35012
rect 22796 35000 22802 35012
rect 23308 35000 23336 35031
rect 22796 34972 23336 35000
rect 22796 34960 22802 34972
rect 24118 34960 24124 35012
rect 24176 35000 24182 35012
rect 24780 35000 24808 35031
rect 24946 35028 24952 35080
rect 25004 35068 25010 35080
rect 25884 35077 25912 35108
rect 25958 35096 25964 35108
rect 26016 35096 26022 35148
rect 26510 35136 26516 35148
rect 26471 35108 26516 35136
rect 26510 35096 26516 35108
rect 26568 35096 26574 35148
rect 27522 35136 27528 35148
rect 27483 35108 27528 35136
rect 27522 35096 27528 35108
rect 27580 35096 27586 35148
rect 25225 35071 25283 35077
rect 25225 35068 25237 35071
rect 25004 35040 25237 35068
rect 25004 35028 25010 35040
rect 25225 35037 25237 35040
rect 25271 35037 25283 35071
rect 25225 35031 25283 35037
rect 25869 35071 25927 35077
rect 25869 35037 25881 35071
rect 25915 35037 25927 35071
rect 25869 35031 25927 35037
rect 24176 34972 24808 35000
rect 24176 34960 24182 34972
rect 17954 34892 17960 34944
rect 18012 34932 18018 34944
rect 18233 34935 18291 34941
rect 18233 34932 18245 34935
rect 18012 34904 18245 34932
rect 18012 34892 18018 34904
rect 18233 34901 18245 34904
rect 18279 34932 18291 34935
rect 18874 34932 18880 34944
rect 18279 34904 18880 34932
rect 18279 34901 18291 34904
rect 18233 34895 18291 34901
rect 18874 34892 18880 34904
rect 18932 34892 18938 34944
rect 25884 34932 25912 35031
rect 25961 35003 26019 35009
rect 25961 34969 25973 35003
rect 26007 35000 26019 35003
rect 26697 35003 26755 35009
rect 26697 35000 26709 35003
rect 26007 34972 26709 35000
rect 26007 34969 26019 34972
rect 25961 34963 26019 34969
rect 26697 34969 26709 34972
rect 26743 34969 26755 35003
rect 26697 34963 26755 34969
rect 27890 34932 27896 34944
rect 25884 34904 27896 34932
rect 27890 34892 27896 34904
rect 27948 34892 27954 34944
rect 1104 34842 29048 34864
rect 1104 34790 7896 34842
rect 7948 34790 7960 34842
rect 8012 34790 8024 34842
rect 8076 34790 8088 34842
rect 8140 34790 8152 34842
rect 8204 34790 14842 34842
rect 14894 34790 14906 34842
rect 14958 34790 14970 34842
rect 15022 34790 15034 34842
rect 15086 34790 15098 34842
rect 15150 34790 21788 34842
rect 21840 34790 21852 34842
rect 21904 34790 21916 34842
rect 21968 34790 21980 34842
rect 22032 34790 22044 34842
rect 22096 34790 28734 34842
rect 28786 34790 28798 34842
rect 28850 34790 28862 34842
rect 28914 34790 28926 34842
rect 28978 34790 28990 34842
rect 29042 34790 29048 34842
rect 1104 34768 29048 34790
rect 19334 34688 19340 34740
rect 19392 34728 19398 34740
rect 19429 34731 19487 34737
rect 19429 34728 19441 34731
rect 19392 34700 19441 34728
rect 19392 34688 19398 34700
rect 19429 34697 19441 34700
rect 19475 34697 19487 34731
rect 26602 34728 26608 34740
rect 26515 34700 26608 34728
rect 19429 34691 19487 34697
rect 26602 34688 26608 34700
rect 26660 34728 26666 34740
rect 26660 34700 27752 34728
rect 26660 34688 26666 34700
rect 14734 34620 14740 34672
rect 14792 34660 14798 34672
rect 24946 34660 24952 34672
rect 14792 34632 24952 34660
rect 14792 34620 14798 34632
rect 24946 34620 24952 34632
rect 25004 34620 25010 34672
rect 25492 34663 25550 34669
rect 25492 34629 25504 34663
rect 25538 34660 25550 34663
rect 25682 34660 25688 34672
rect 25538 34632 25688 34660
rect 25538 34629 25550 34632
rect 25492 34623 25550 34629
rect 25682 34620 25688 34632
rect 25740 34620 25746 34672
rect 19521 34595 19579 34601
rect 19521 34561 19533 34595
rect 19567 34592 19579 34595
rect 19610 34592 19616 34604
rect 19567 34564 19616 34592
rect 19567 34561 19579 34564
rect 19521 34555 19579 34561
rect 19610 34552 19616 34564
rect 19668 34552 19674 34604
rect 24854 34552 24860 34604
rect 24912 34592 24918 34604
rect 27724 34601 27752 34700
rect 25225 34595 25283 34601
rect 25225 34592 25237 34595
rect 24912 34564 25237 34592
rect 24912 34552 24918 34564
rect 25225 34561 25237 34564
rect 25271 34561 25283 34595
rect 25225 34555 25283 34561
rect 27709 34595 27767 34601
rect 27709 34561 27721 34595
rect 27755 34561 27767 34595
rect 27709 34555 27767 34561
rect 1670 34524 1676 34536
rect 1631 34496 1676 34524
rect 1670 34484 1676 34496
rect 1728 34484 1734 34536
rect 1854 34524 1860 34536
rect 1815 34496 1860 34524
rect 1854 34484 1860 34496
rect 1912 34484 1918 34536
rect 2774 34524 2780 34536
rect 2735 34496 2780 34524
rect 2774 34484 2780 34496
rect 2832 34484 2838 34536
rect 16666 34484 16672 34536
rect 16724 34524 16730 34536
rect 19702 34524 19708 34536
rect 16724 34496 19708 34524
rect 16724 34484 16730 34496
rect 19702 34484 19708 34496
rect 19760 34484 19766 34536
rect 27154 34388 27160 34400
rect 27115 34360 27160 34388
rect 27154 34348 27160 34360
rect 27212 34348 27218 34400
rect 1104 34298 28888 34320
rect 1104 34246 4423 34298
rect 4475 34246 4487 34298
rect 4539 34246 4551 34298
rect 4603 34246 4615 34298
rect 4667 34246 4679 34298
rect 4731 34246 11369 34298
rect 11421 34246 11433 34298
rect 11485 34246 11497 34298
rect 11549 34246 11561 34298
rect 11613 34246 11625 34298
rect 11677 34246 18315 34298
rect 18367 34246 18379 34298
rect 18431 34246 18443 34298
rect 18495 34246 18507 34298
rect 18559 34246 18571 34298
rect 18623 34246 25261 34298
rect 25313 34246 25325 34298
rect 25377 34246 25389 34298
rect 25441 34246 25453 34298
rect 25505 34246 25517 34298
rect 25569 34246 28888 34298
rect 1104 34224 28888 34246
rect 1854 34144 1860 34196
rect 1912 34184 1918 34196
rect 2133 34187 2191 34193
rect 2133 34184 2145 34187
rect 1912 34156 2145 34184
rect 1912 34144 1918 34156
rect 2133 34153 2145 34156
rect 2179 34153 2191 34187
rect 2133 34147 2191 34153
rect 21085 34187 21143 34193
rect 21085 34153 21097 34187
rect 21131 34184 21143 34187
rect 21450 34184 21456 34196
rect 21131 34156 21456 34184
rect 21131 34153 21143 34156
rect 21085 34147 21143 34153
rect 21450 34144 21456 34156
rect 21508 34144 21514 34196
rect 26142 34076 26148 34128
rect 26200 34116 26206 34128
rect 26200 34088 26740 34116
rect 26200 34076 26206 34088
rect 26602 34048 26608 34060
rect 24872 34020 26608 34048
rect 2225 33983 2283 33989
rect 2225 33949 2237 33983
rect 2271 33980 2283 33983
rect 2314 33980 2320 33992
rect 2271 33952 2320 33980
rect 2271 33949 2283 33952
rect 2225 33943 2283 33949
rect 2314 33940 2320 33952
rect 2372 33980 2378 33992
rect 4338 33980 4344 33992
rect 2372 33952 4344 33980
rect 2372 33940 2378 33952
rect 4338 33940 4344 33952
rect 4396 33940 4402 33992
rect 22462 33980 22468 33992
rect 22423 33952 22468 33980
rect 22462 33940 22468 33952
rect 22520 33940 22526 33992
rect 23109 33983 23167 33989
rect 23109 33949 23121 33983
rect 23155 33980 23167 33983
rect 23750 33980 23756 33992
rect 23155 33952 23756 33980
rect 23155 33949 23167 33952
rect 23109 33943 23167 33949
rect 23750 33940 23756 33952
rect 23808 33940 23814 33992
rect 24670 33980 24676 33992
rect 24631 33952 24676 33980
rect 24670 33940 24676 33952
rect 24728 33940 24734 33992
rect 24872 33989 24900 34020
rect 26602 34008 26608 34020
rect 26660 34008 26666 34060
rect 26712 34057 26740 34088
rect 26697 34051 26755 34057
rect 26697 34017 26709 34051
rect 26743 34017 26755 34051
rect 26697 34011 26755 34017
rect 24857 33983 24915 33989
rect 24857 33949 24869 33983
rect 24903 33949 24915 33983
rect 24857 33943 24915 33949
rect 26237 33983 26295 33989
rect 26237 33949 26249 33983
rect 26283 33949 26295 33983
rect 26237 33943 26295 33949
rect 22186 33912 22192 33924
rect 22244 33921 22250 33924
rect 22156 33884 22192 33912
rect 22186 33872 22192 33884
rect 22244 33875 22256 33921
rect 22244 33872 22250 33875
rect 26252 33856 26280 33943
rect 26421 33915 26479 33921
rect 26421 33881 26433 33915
rect 26467 33912 26479 33915
rect 27246 33912 27252 33924
rect 26467 33884 27252 33912
rect 26467 33881 26479 33884
rect 26421 33875 26479 33881
rect 27246 33872 27252 33884
rect 27304 33872 27310 33924
rect 20714 33804 20720 33856
rect 20772 33844 20778 33856
rect 23017 33847 23075 33853
rect 23017 33844 23029 33847
rect 20772 33816 23029 33844
rect 20772 33804 20778 33816
rect 23017 33813 23029 33816
rect 23063 33813 23075 33847
rect 23017 33807 23075 33813
rect 24765 33847 24823 33853
rect 24765 33813 24777 33847
rect 24811 33844 24823 33847
rect 24946 33844 24952 33856
rect 24811 33816 24952 33844
rect 24811 33813 24823 33816
rect 24765 33807 24823 33813
rect 24946 33804 24952 33816
rect 25004 33804 25010 33856
rect 26234 33804 26240 33856
rect 26292 33804 26298 33856
rect 1104 33754 29048 33776
rect 1104 33702 7896 33754
rect 7948 33702 7960 33754
rect 8012 33702 8024 33754
rect 8076 33702 8088 33754
rect 8140 33702 8152 33754
rect 8204 33702 14842 33754
rect 14894 33702 14906 33754
rect 14958 33702 14970 33754
rect 15022 33702 15034 33754
rect 15086 33702 15098 33754
rect 15150 33702 21788 33754
rect 21840 33702 21852 33754
rect 21904 33702 21916 33754
rect 21968 33702 21980 33754
rect 22032 33702 22044 33754
rect 22096 33702 28734 33754
rect 28786 33702 28798 33754
rect 28850 33702 28862 33754
rect 28914 33702 28926 33754
rect 28978 33702 28990 33754
rect 29042 33702 29048 33754
rect 1104 33680 29048 33702
rect 20898 33640 20904 33652
rect 20272 33612 20904 33640
rect 18690 33532 18696 33584
rect 18748 33572 18754 33584
rect 18969 33575 19027 33581
rect 18969 33572 18981 33575
rect 18748 33544 18981 33572
rect 18748 33532 18754 33544
rect 18969 33541 18981 33544
rect 19015 33541 19027 33575
rect 18969 33535 19027 33541
rect 19185 33575 19243 33581
rect 19185 33541 19197 33575
rect 19231 33572 19243 33575
rect 19426 33572 19432 33584
rect 19231 33544 19432 33572
rect 19231 33541 19243 33544
rect 19185 33535 19243 33541
rect 19426 33532 19432 33544
rect 19484 33532 19490 33584
rect 1670 33464 1676 33516
rect 1728 33504 1734 33516
rect 1765 33507 1823 33513
rect 1765 33504 1777 33507
rect 1728 33476 1777 33504
rect 1728 33464 1734 33476
rect 1765 33473 1777 33476
rect 1811 33473 1823 33507
rect 17954 33504 17960 33516
rect 17915 33476 17960 33504
rect 1765 33467 1823 33473
rect 17954 33464 17960 33476
rect 18012 33464 18018 33516
rect 18138 33464 18144 33516
rect 18196 33504 18202 33516
rect 18233 33507 18291 33513
rect 18233 33504 18245 33507
rect 18196 33476 18245 33504
rect 18196 33464 18202 33476
rect 18233 33473 18245 33476
rect 18279 33473 18291 33507
rect 18233 33467 18291 33473
rect 18325 33507 18383 33513
rect 18325 33473 18337 33507
rect 18371 33504 18383 33507
rect 18874 33504 18880 33516
rect 18371 33476 18880 33504
rect 18371 33473 18383 33476
rect 18325 33467 18383 33473
rect 18874 33464 18880 33476
rect 18932 33464 18938 33516
rect 20165 33507 20223 33513
rect 20165 33473 20177 33507
rect 20211 33504 20223 33507
rect 20272 33504 20300 33612
rect 20898 33600 20904 33612
rect 20956 33640 20962 33652
rect 21634 33640 21640 33652
rect 20956 33612 21640 33640
rect 20956 33600 20962 33612
rect 21634 33600 21640 33612
rect 21692 33600 21698 33652
rect 22186 33640 22192 33652
rect 22147 33612 22192 33640
rect 22186 33600 22192 33612
rect 22244 33600 22250 33652
rect 27246 33640 27252 33652
rect 27207 33612 27252 33640
rect 27246 33600 27252 33612
rect 27304 33600 27310 33652
rect 20349 33575 20407 33581
rect 20349 33541 20361 33575
rect 20395 33572 20407 33575
rect 20714 33572 20720 33584
rect 20395 33544 20720 33572
rect 20395 33541 20407 33544
rect 20349 33535 20407 33541
rect 20714 33532 20720 33544
rect 20772 33532 20778 33584
rect 24854 33532 24860 33584
rect 24912 33572 24918 33584
rect 24912 33544 26096 33572
rect 24912 33532 24918 33544
rect 20438 33504 20444 33516
rect 20211 33476 20300 33504
rect 20399 33476 20444 33504
rect 20211 33473 20223 33476
rect 20165 33467 20223 33473
rect 20438 33464 20444 33476
rect 20496 33464 20502 33516
rect 20533 33507 20591 33513
rect 20533 33473 20545 33507
rect 20579 33473 20591 33507
rect 20533 33467 20591 33473
rect 22005 33507 22063 33513
rect 22005 33473 22017 33507
rect 22051 33504 22063 33507
rect 22278 33504 22284 33516
rect 22051 33476 22284 33504
rect 22051 33473 22063 33476
rect 22005 33467 22063 33473
rect 19978 33396 19984 33448
rect 20036 33436 20042 33448
rect 20548 33436 20576 33467
rect 22278 33464 22284 33476
rect 22336 33464 22342 33516
rect 23382 33504 23388 33516
rect 23343 33476 23388 33504
rect 23382 33464 23388 33476
rect 23440 33464 23446 33516
rect 24026 33504 24032 33516
rect 23987 33476 24032 33504
rect 24026 33464 24032 33476
rect 24084 33464 24090 33516
rect 26068 33513 26096 33544
rect 25797 33507 25855 33513
rect 25797 33473 25809 33507
rect 25843 33504 25855 33507
rect 26053 33507 26111 33513
rect 25843 33476 26004 33504
rect 25843 33473 25855 33476
rect 25797 33467 25855 33473
rect 23937 33439 23995 33445
rect 23937 33436 23949 33439
rect 20036 33408 23949 33436
rect 20036 33396 20042 33408
rect 23937 33405 23949 33408
rect 23983 33405 23995 33439
rect 25976 33436 26004 33476
rect 26053 33473 26065 33507
rect 26099 33473 26111 33507
rect 26053 33467 26111 33473
rect 26878 33464 26884 33516
rect 26936 33504 26942 33516
rect 27341 33507 27399 33513
rect 27341 33504 27353 33507
rect 26936 33476 27353 33504
rect 26936 33464 26942 33476
rect 27341 33473 27353 33476
rect 27387 33504 27399 33507
rect 28166 33504 28172 33516
rect 27387 33476 28172 33504
rect 27387 33473 27399 33476
rect 27341 33467 27399 33473
rect 28166 33464 28172 33476
rect 28224 33464 28230 33516
rect 27154 33436 27160 33448
rect 25976 33408 27160 33436
rect 23937 33399 23995 33405
rect 27154 33396 27160 33408
rect 27212 33396 27218 33448
rect 3510 33328 3516 33380
rect 3568 33368 3574 33380
rect 9122 33368 9128 33380
rect 3568 33340 9128 33368
rect 3568 33328 3574 33340
rect 9122 33328 9128 33340
rect 9180 33328 9186 33380
rect 16758 33328 16764 33380
rect 16816 33368 16822 33380
rect 18049 33371 18107 33377
rect 18049 33368 18061 33371
rect 16816 33340 18061 33368
rect 16816 33328 16822 33340
rect 18049 33337 18061 33340
rect 18095 33368 18107 33371
rect 18966 33368 18972 33380
rect 18095 33340 18972 33368
rect 18095 33337 18107 33340
rect 18049 33331 18107 33337
rect 18966 33328 18972 33340
rect 19024 33328 19030 33380
rect 26694 33328 26700 33380
rect 26752 33368 26758 33380
rect 26878 33368 26884 33380
rect 26752 33340 26884 33368
rect 26752 33328 26758 33340
rect 26878 33328 26884 33340
rect 26936 33328 26942 33380
rect 18138 33260 18144 33312
rect 18196 33300 18202 33312
rect 18509 33303 18567 33309
rect 18509 33300 18521 33303
rect 18196 33272 18521 33300
rect 18196 33260 18202 33272
rect 18509 33269 18521 33272
rect 18555 33300 18567 33303
rect 19153 33303 19211 33309
rect 19153 33300 19165 33303
rect 18555 33272 19165 33300
rect 18555 33269 18567 33272
rect 18509 33263 18567 33269
rect 19153 33269 19165 33272
rect 19199 33269 19211 33303
rect 19334 33300 19340 33312
rect 19295 33272 19340 33300
rect 19153 33263 19211 33269
rect 19334 33260 19340 33272
rect 19392 33260 19398 33312
rect 20717 33303 20775 33309
rect 20717 33269 20729 33303
rect 20763 33300 20775 33303
rect 21910 33300 21916 33312
rect 20763 33272 21916 33300
rect 20763 33269 20775 33272
rect 20717 33263 20775 33269
rect 21910 33260 21916 33272
rect 21968 33260 21974 33312
rect 23198 33300 23204 33312
rect 23159 33272 23204 33300
rect 23198 33260 23204 33272
rect 23256 33260 23262 33312
rect 24673 33303 24731 33309
rect 24673 33269 24685 33303
rect 24719 33300 24731 33303
rect 25038 33300 25044 33312
rect 24719 33272 25044 33300
rect 24719 33269 24731 33272
rect 24673 33263 24731 33269
rect 25038 33260 25044 33272
rect 25096 33260 25102 33312
rect 28077 33303 28135 33309
rect 28077 33269 28089 33303
rect 28123 33300 28135 33303
rect 28258 33300 28264 33312
rect 28123 33272 28264 33300
rect 28123 33269 28135 33272
rect 28077 33263 28135 33269
rect 28258 33260 28264 33272
rect 28316 33260 28322 33312
rect 1104 33210 28888 33232
rect 1104 33158 4423 33210
rect 4475 33158 4487 33210
rect 4539 33158 4551 33210
rect 4603 33158 4615 33210
rect 4667 33158 4679 33210
rect 4731 33158 11369 33210
rect 11421 33158 11433 33210
rect 11485 33158 11497 33210
rect 11549 33158 11561 33210
rect 11613 33158 11625 33210
rect 11677 33158 18315 33210
rect 18367 33158 18379 33210
rect 18431 33158 18443 33210
rect 18495 33158 18507 33210
rect 18559 33158 18571 33210
rect 18623 33158 25261 33210
rect 25313 33158 25325 33210
rect 25377 33158 25389 33210
rect 25441 33158 25453 33210
rect 25505 33158 25517 33210
rect 25569 33158 28888 33210
rect 1104 33136 28888 33158
rect 16945 33099 17003 33105
rect 16945 33065 16957 33099
rect 16991 33096 17003 33099
rect 17862 33096 17868 33108
rect 16991 33068 17868 33096
rect 16991 33065 17003 33068
rect 16945 33059 17003 33065
rect 17862 33056 17868 33068
rect 17920 33056 17926 33108
rect 17954 33056 17960 33108
rect 18012 33096 18018 33108
rect 18230 33096 18236 33108
rect 18012 33068 18236 33096
rect 18012 33056 18018 33068
rect 18230 33056 18236 33068
rect 18288 33056 18294 33108
rect 19426 33096 19432 33108
rect 19387 33068 19432 33096
rect 19426 33056 19432 33068
rect 19484 33056 19490 33108
rect 19886 33056 19892 33108
rect 19944 33096 19950 33108
rect 20438 33096 20444 33108
rect 19944 33068 20444 33096
rect 19944 33056 19950 33068
rect 20438 33056 20444 33068
rect 20496 33056 20502 33108
rect 20714 33096 20720 33108
rect 20675 33068 20720 33096
rect 20714 33056 20720 33068
rect 20772 33056 20778 33108
rect 24026 33096 24032 33108
rect 20824 33068 21036 33096
rect 23987 33068 24032 33096
rect 16758 33028 16764 33040
rect 16132 33000 16764 33028
rect 1670 32892 1676 32904
rect 1631 32864 1676 32892
rect 1670 32852 1676 32864
rect 1728 32852 1734 32904
rect 15286 32892 15292 32904
rect 15247 32864 15292 32892
rect 15286 32852 15292 32864
rect 15344 32852 15350 32904
rect 16132 32901 16160 33000
rect 16758 32988 16764 33000
rect 16816 32988 16822 33040
rect 16868 33000 17264 33028
rect 16206 32920 16212 32972
rect 16264 32960 16270 32972
rect 16868 32960 16896 33000
rect 16264 32932 16309 32960
rect 16546 32932 16896 32960
rect 16264 32920 16270 32932
rect 15473 32895 15531 32901
rect 15473 32861 15485 32895
rect 15519 32892 15531 32895
rect 16117 32895 16175 32901
rect 15519 32864 15976 32892
rect 15519 32861 15531 32864
rect 15473 32855 15531 32861
rect 15948 32836 15976 32864
rect 16117 32861 16129 32895
rect 16163 32861 16175 32895
rect 16117 32855 16175 32861
rect 16337 32895 16395 32901
rect 16337 32861 16349 32895
rect 16383 32892 16395 32895
rect 16546 32892 16574 32932
rect 16383 32864 16574 32892
rect 16383 32861 16395 32864
rect 16337 32855 16395 32861
rect 16758 32852 16764 32904
rect 16816 32892 16822 32904
rect 17236 32901 17264 33000
rect 18782 32988 18788 33040
rect 18840 33028 18846 33040
rect 18840 33000 20208 33028
rect 18840 32988 18846 33000
rect 17405 32963 17463 32969
rect 17405 32929 17417 32963
rect 17451 32960 17463 32963
rect 18690 32960 18696 32972
rect 17451 32932 18696 32960
rect 17451 32929 17463 32932
rect 17405 32923 17463 32929
rect 18690 32920 18696 32932
rect 18748 32920 18754 32972
rect 19886 32960 19892 32972
rect 19847 32932 19892 32960
rect 19886 32920 19892 32932
rect 19944 32920 19950 32972
rect 16853 32895 16911 32901
rect 16853 32892 16865 32895
rect 16816 32864 16865 32892
rect 16816 32852 16822 32864
rect 16853 32861 16865 32864
rect 16899 32861 16911 32895
rect 16853 32855 16911 32861
rect 17129 32895 17187 32901
rect 17129 32861 17141 32895
rect 17175 32861 17187 32895
rect 17129 32855 17187 32861
rect 17221 32895 17279 32901
rect 17221 32861 17233 32895
rect 17267 32892 17279 32895
rect 18046 32892 18052 32904
rect 17267 32864 18052 32892
rect 17267 32861 17279 32864
rect 17221 32855 17279 32861
rect 15930 32824 15936 32836
rect 15891 32796 15936 32824
rect 15930 32784 15936 32796
rect 15988 32784 15994 32836
rect 16209 32827 16267 32833
rect 16209 32793 16221 32827
rect 16255 32824 16267 32827
rect 17144 32824 17172 32855
rect 18046 32852 18052 32864
rect 18104 32852 18110 32904
rect 18322 32852 18328 32904
rect 18380 32892 18386 32904
rect 18417 32895 18475 32901
rect 18417 32892 18429 32895
rect 18380 32864 18429 32892
rect 18380 32852 18386 32864
rect 18417 32861 18429 32864
rect 18463 32861 18475 32895
rect 19610 32892 19616 32904
rect 19571 32864 19616 32892
rect 18417 32855 18475 32861
rect 19610 32852 19616 32864
rect 19668 32852 19674 32904
rect 19794 32892 19800 32904
rect 19755 32864 19800 32892
rect 19794 32852 19800 32864
rect 19852 32852 19858 32904
rect 19978 32892 19984 32904
rect 19939 32864 19984 32892
rect 19978 32852 19984 32864
rect 20036 32852 20042 32904
rect 20180 32901 20208 33000
rect 20346 32988 20352 33040
rect 20404 33028 20410 33040
rect 20824 33028 20852 33068
rect 20404 33000 20852 33028
rect 20404 32988 20410 33000
rect 20898 32988 20904 33040
rect 20956 32988 20962 33040
rect 20916 32960 20944 32988
rect 20640 32932 20944 32960
rect 20640 32901 20668 32932
rect 20165 32895 20223 32901
rect 20165 32861 20177 32895
rect 20211 32861 20223 32895
rect 20165 32855 20223 32861
rect 20625 32895 20683 32901
rect 20625 32861 20637 32895
rect 20671 32861 20683 32895
rect 20625 32855 20683 32861
rect 20806 32852 20812 32904
rect 20864 32892 20870 32904
rect 21008 32901 21036 33068
rect 24026 33056 24032 33068
rect 24084 33056 24090 33108
rect 24670 32988 24676 33040
rect 24728 33028 24734 33040
rect 24728 33000 25268 33028
rect 24728 32988 24734 33000
rect 25130 32960 25136 32972
rect 25091 32932 25136 32960
rect 25130 32920 25136 32932
rect 25188 32920 25194 32972
rect 25240 32969 25268 33000
rect 25225 32963 25283 32969
rect 25225 32929 25237 32963
rect 25271 32929 25283 32963
rect 27522 32960 27528 32972
rect 27483 32932 27528 32960
rect 25225 32923 25283 32929
rect 27522 32920 27528 32932
rect 27580 32920 27586 32972
rect 20901 32895 20959 32901
rect 20901 32892 20913 32895
rect 20864 32864 20913 32892
rect 20864 32852 20870 32864
rect 20901 32861 20913 32864
rect 20947 32861 20959 32895
rect 20901 32855 20959 32861
rect 20993 32895 21051 32901
rect 20993 32861 21005 32895
rect 21039 32861 21051 32895
rect 20993 32855 21051 32861
rect 21177 32895 21235 32901
rect 21177 32861 21189 32895
rect 21223 32892 21235 32895
rect 21637 32895 21695 32901
rect 21637 32892 21649 32895
rect 21223 32864 21649 32892
rect 21223 32861 21235 32864
rect 21177 32855 21235 32861
rect 21637 32861 21649 32864
rect 21683 32861 21695 32895
rect 21910 32892 21916 32904
rect 21871 32864 21916 32892
rect 21637 32855 21695 32861
rect 21910 32852 21916 32864
rect 21968 32852 21974 32904
rect 22186 32852 22192 32904
rect 22244 32892 22250 32904
rect 22462 32892 22468 32904
rect 22244 32864 22468 32892
rect 22244 32852 22250 32864
rect 22462 32852 22468 32864
rect 22520 32892 22526 32904
rect 22649 32895 22707 32901
rect 22649 32892 22661 32895
rect 22520 32864 22661 32892
rect 22520 32852 22526 32864
rect 22649 32861 22661 32864
rect 22695 32861 22707 32895
rect 22649 32855 22707 32861
rect 22916 32895 22974 32901
rect 22916 32861 22928 32895
rect 22962 32892 22974 32895
rect 23198 32892 23204 32904
rect 22962 32864 23204 32892
rect 22962 32861 22974 32864
rect 22916 32855 22974 32861
rect 23198 32852 23204 32864
rect 23256 32852 23262 32904
rect 24854 32892 24860 32904
rect 24815 32864 24860 32892
rect 24854 32852 24860 32864
rect 24912 32852 24918 32904
rect 24949 32895 25007 32901
rect 24949 32861 24961 32895
rect 24995 32892 25007 32895
rect 25038 32892 25044 32904
rect 24995 32864 25044 32892
rect 24995 32861 25007 32864
rect 24949 32855 25007 32861
rect 25038 32852 25044 32864
rect 25096 32852 25102 32904
rect 26510 32892 26516 32904
rect 26471 32864 26516 32892
rect 26510 32852 26516 32864
rect 26568 32852 26574 32904
rect 18141 32827 18199 32833
rect 18141 32824 18153 32827
rect 16255 32796 16574 32824
rect 16255 32793 16267 32796
rect 16209 32787 16267 32793
rect 16546 32768 16574 32796
rect 17144 32796 18153 32824
rect 15470 32756 15476 32768
rect 15431 32728 15476 32756
rect 15470 32716 15476 32728
rect 15528 32716 15534 32768
rect 16546 32728 16580 32768
rect 16574 32716 16580 32728
rect 16632 32756 16638 32768
rect 17144 32756 17172 32796
rect 18141 32793 18153 32796
rect 18187 32793 18199 32827
rect 18141 32787 18199 32793
rect 18233 32827 18291 32833
rect 18233 32793 18245 32827
rect 18279 32824 18291 32827
rect 18966 32824 18972 32836
rect 18279 32796 18972 32824
rect 18279 32793 18291 32796
rect 18233 32787 18291 32793
rect 18966 32784 18972 32796
rect 19024 32784 19030 32836
rect 19150 32784 19156 32836
rect 19208 32824 19214 32836
rect 22097 32827 22155 32833
rect 22097 32824 22109 32827
rect 19208 32796 22109 32824
rect 19208 32784 19214 32796
rect 22097 32793 22109 32796
rect 22143 32793 22155 32827
rect 22097 32787 22155 32793
rect 26697 32827 26755 32833
rect 26697 32793 26709 32827
rect 26743 32824 26755 32827
rect 28074 32824 28080 32836
rect 26743 32796 28080 32824
rect 26743 32793 26755 32796
rect 26697 32787 26755 32793
rect 28074 32784 28080 32796
rect 28132 32784 28138 32836
rect 16632 32728 17172 32756
rect 17865 32759 17923 32765
rect 16632 32716 16638 32728
rect 17865 32725 17877 32759
rect 17911 32756 17923 32759
rect 18046 32756 18052 32768
rect 17911 32728 18052 32756
rect 17911 32725 17923 32728
rect 17865 32719 17923 32725
rect 18046 32716 18052 32728
rect 18104 32716 18110 32768
rect 20530 32716 20536 32768
rect 20588 32756 20594 32768
rect 21729 32759 21787 32765
rect 21729 32756 21741 32759
rect 20588 32728 21741 32756
rect 20588 32716 20594 32728
rect 21729 32725 21741 32728
rect 21775 32725 21787 32759
rect 24670 32756 24676 32768
rect 24631 32728 24676 32756
rect 21729 32719 21787 32725
rect 24670 32716 24676 32728
rect 24728 32716 24734 32768
rect 1104 32666 29048 32688
rect 1104 32614 7896 32666
rect 7948 32614 7960 32666
rect 8012 32614 8024 32666
rect 8076 32614 8088 32666
rect 8140 32614 8152 32666
rect 8204 32614 14842 32666
rect 14894 32614 14906 32666
rect 14958 32614 14970 32666
rect 15022 32614 15034 32666
rect 15086 32614 15098 32666
rect 15150 32614 21788 32666
rect 21840 32614 21852 32666
rect 21904 32614 21916 32666
rect 21968 32614 21980 32666
rect 22032 32614 22044 32666
rect 22096 32614 28734 32666
rect 28786 32614 28798 32666
rect 28850 32614 28862 32666
rect 28914 32614 28926 32666
rect 28978 32614 28990 32666
rect 29042 32614 29048 32666
rect 1104 32592 29048 32614
rect 15470 32512 15476 32564
rect 15528 32552 15534 32564
rect 15949 32555 16007 32561
rect 15949 32552 15961 32555
rect 15528 32524 15961 32552
rect 15528 32512 15534 32524
rect 15949 32521 15961 32524
rect 15995 32521 16007 32555
rect 15949 32515 16007 32521
rect 16206 32512 16212 32564
rect 16264 32552 16270 32564
rect 20530 32552 20536 32564
rect 16264 32524 19104 32552
rect 20491 32524 20536 32552
rect 16264 32512 16270 32524
rect 15286 32484 15292 32496
rect 15247 32456 15292 32484
rect 15286 32444 15292 32456
rect 15344 32444 15350 32496
rect 15746 32484 15752 32496
rect 15707 32456 15752 32484
rect 15746 32444 15752 32456
rect 15804 32444 15810 32496
rect 19076 32493 19104 32524
rect 20530 32512 20536 32524
rect 20588 32512 20594 32564
rect 24026 32512 24032 32564
rect 24084 32552 24090 32564
rect 24305 32555 24363 32561
rect 24305 32552 24317 32555
rect 24084 32524 24317 32552
rect 24084 32512 24090 32524
rect 24305 32521 24317 32524
rect 24351 32521 24363 32555
rect 28074 32552 28080 32564
rect 28035 32524 28080 32552
rect 24305 32515 24363 32521
rect 28074 32512 28080 32524
rect 28132 32512 28138 32564
rect 18325 32487 18383 32493
rect 18325 32453 18337 32487
rect 18371 32484 18383 32487
rect 18923 32487 18981 32493
rect 18923 32484 18935 32487
rect 18371 32456 18935 32484
rect 18371 32453 18383 32456
rect 18325 32447 18383 32453
rect 18923 32453 18935 32456
rect 18969 32453 18981 32487
rect 18923 32447 18981 32453
rect 19061 32487 19119 32493
rect 19061 32453 19073 32487
rect 19107 32453 19119 32487
rect 19061 32447 19119 32453
rect 19150 32444 19156 32496
rect 19208 32484 19214 32496
rect 20806 32484 20812 32496
rect 19208 32456 19253 32484
rect 20272 32456 20812 32484
rect 19208 32444 19214 32456
rect 1670 32416 1676 32428
rect 1631 32388 1676 32416
rect 1670 32376 1676 32388
rect 1728 32376 1734 32428
rect 15105 32419 15163 32425
rect 15105 32385 15117 32419
rect 15151 32385 15163 32419
rect 16853 32419 16911 32425
rect 16853 32416 16865 32419
rect 15105 32379 15163 32385
rect 16546 32388 16865 32416
rect 1857 32351 1915 32357
rect 1857 32317 1869 32351
rect 1903 32348 1915 32351
rect 2038 32348 2044 32360
rect 1903 32320 2044 32348
rect 1903 32317 1915 32320
rect 1857 32311 1915 32317
rect 2038 32308 2044 32320
rect 2096 32308 2102 32360
rect 2774 32348 2780 32360
rect 2735 32320 2780 32348
rect 2774 32308 2780 32320
rect 2832 32308 2838 32360
rect 15120 32348 15148 32379
rect 15930 32348 15936 32360
rect 15120 32320 15936 32348
rect 15930 32308 15936 32320
rect 15988 32308 15994 32360
rect 16117 32283 16175 32289
rect 16117 32249 16129 32283
rect 16163 32280 16175 32283
rect 16546 32280 16574 32388
rect 16853 32385 16865 32388
rect 16899 32385 16911 32419
rect 18046 32416 18052 32428
rect 18007 32388 18052 32416
rect 16853 32379 16911 32385
rect 18046 32376 18052 32388
rect 18104 32376 18110 32428
rect 18138 32376 18144 32428
rect 18196 32416 18202 32428
rect 19245 32419 19303 32425
rect 18196 32388 18241 32416
rect 18196 32376 18202 32388
rect 19245 32385 19257 32419
rect 19291 32416 19303 32419
rect 19334 32416 19340 32428
rect 19291 32388 19340 32416
rect 19291 32385 19303 32388
rect 19245 32379 19303 32385
rect 19334 32376 19340 32388
rect 19392 32376 19398 32428
rect 19981 32419 20039 32425
rect 19981 32385 19993 32419
rect 20027 32385 20039 32419
rect 19981 32379 20039 32385
rect 18325 32351 18383 32357
rect 18325 32317 18337 32351
rect 18371 32348 18383 32351
rect 18690 32348 18696 32360
rect 18371 32320 18696 32348
rect 18371 32317 18383 32320
rect 18325 32311 18383 32317
rect 18690 32308 18696 32320
rect 18748 32308 18754 32360
rect 18782 32308 18788 32360
rect 18840 32348 18846 32360
rect 19996 32348 20024 32379
rect 20070 32376 20076 32428
rect 20128 32416 20134 32428
rect 20272 32425 20300 32456
rect 20806 32444 20812 32456
rect 20864 32444 20870 32496
rect 24397 32487 24455 32493
rect 24397 32453 24409 32487
rect 24443 32484 24455 32487
rect 26418 32484 26424 32496
rect 24443 32456 26424 32484
rect 24443 32453 24455 32456
rect 24397 32447 24455 32453
rect 26418 32444 26424 32456
rect 26476 32444 26482 32496
rect 20257 32419 20315 32425
rect 20128 32388 20173 32416
rect 20128 32376 20134 32388
rect 20257 32385 20269 32419
rect 20303 32385 20315 32419
rect 20257 32379 20315 32385
rect 20346 32376 20352 32428
rect 20404 32416 20410 32428
rect 22005 32419 22063 32425
rect 20404 32388 20449 32416
rect 20404 32376 20410 32388
rect 22005 32385 22017 32419
rect 22051 32416 22063 32419
rect 22094 32416 22100 32428
rect 22051 32388 22100 32416
rect 22051 32385 22063 32388
rect 22005 32379 22063 32385
rect 22094 32376 22100 32388
rect 22152 32376 22158 32428
rect 22272 32419 22330 32425
rect 22272 32385 22284 32419
rect 22318 32416 22330 32419
rect 22646 32416 22652 32428
rect 22318 32388 22652 32416
rect 22318 32385 22330 32388
rect 22272 32379 22330 32385
rect 22646 32376 22652 32388
rect 22704 32376 22710 32428
rect 26510 32376 26516 32428
rect 26568 32416 26574 32428
rect 26605 32419 26663 32425
rect 26605 32416 26617 32419
rect 26568 32388 26617 32416
rect 26568 32376 26574 32388
rect 26605 32385 26617 32388
rect 26651 32385 26663 32419
rect 26605 32379 26663 32385
rect 27062 32376 27068 32428
rect 27120 32416 27126 32428
rect 27341 32419 27399 32425
rect 27341 32416 27353 32419
rect 27120 32388 27353 32416
rect 27120 32376 27126 32388
rect 27341 32385 27353 32388
rect 27387 32385 27399 32419
rect 27982 32416 27988 32428
rect 27943 32388 27988 32416
rect 27341 32379 27399 32385
rect 27982 32376 27988 32388
rect 28040 32376 28046 32428
rect 20162 32348 20168 32360
rect 18840 32320 18885 32348
rect 19996 32320 20168 32348
rect 18840 32308 18846 32320
rect 20162 32308 20168 32320
rect 20220 32348 20226 32360
rect 20990 32348 20996 32360
rect 20220 32320 20996 32348
rect 20220 32308 20226 32320
rect 20990 32308 20996 32320
rect 21048 32308 21054 32360
rect 24486 32308 24492 32360
rect 24544 32348 24550 32360
rect 24544 32320 24589 32348
rect 24544 32308 24550 32320
rect 16163 32252 16574 32280
rect 16163 32249 16175 32252
rect 16117 32243 16175 32249
rect 14921 32215 14979 32221
rect 14921 32181 14933 32215
rect 14967 32212 14979 32215
rect 15838 32212 15844 32224
rect 14967 32184 15844 32212
rect 14967 32181 14979 32184
rect 14921 32175 14979 32181
rect 15838 32172 15844 32184
rect 15896 32212 15902 32224
rect 15933 32215 15991 32221
rect 15933 32212 15945 32215
rect 15896 32184 15945 32212
rect 15896 32172 15902 32184
rect 15933 32181 15945 32184
rect 15979 32181 15991 32215
rect 17034 32212 17040 32224
rect 16995 32184 17040 32212
rect 15933 32175 15991 32181
rect 17034 32172 17040 32184
rect 17092 32172 17098 32224
rect 19058 32172 19064 32224
rect 19116 32212 19122 32224
rect 19429 32215 19487 32221
rect 19429 32212 19441 32215
rect 19116 32184 19441 32212
rect 19116 32172 19122 32184
rect 19429 32181 19441 32184
rect 19475 32181 19487 32215
rect 19429 32175 19487 32181
rect 21634 32172 21640 32224
rect 21692 32212 21698 32224
rect 23385 32215 23443 32221
rect 23385 32212 23397 32215
rect 21692 32184 23397 32212
rect 21692 32172 21698 32184
rect 23385 32181 23397 32184
rect 23431 32212 23443 32215
rect 23474 32212 23480 32224
rect 23431 32184 23480 32212
rect 23431 32181 23443 32184
rect 23385 32175 23443 32181
rect 23474 32172 23480 32184
rect 23532 32172 23538 32224
rect 23658 32172 23664 32224
rect 23716 32212 23722 32224
rect 23937 32215 23995 32221
rect 23937 32212 23949 32215
rect 23716 32184 23949 32212
rect 23716 32172 23722 32184
rect 23937 32181 23949 32184
rect 23983 32181 23995 32215
rect 23937 32175 23995 32181
rect 26694 32172 26700 32224
rect 26752 32212 26758 32224
rect 27433 32215 27491 32221
rect 27433 32212 27445 32215
rect 26752 32184 27445 32212
rect 26752 32172 26758 32184
rect 27433 32181 27445 32184
rect 27479 32181 27491 32215
rect 27433 32175 27491 32181
rect 1104 32122 28888 32144
rect 1104 32070 4423 32122
rect 4475 32070 4487 32122
rect 4539 32070 4551 32122
rect 4603 32070 4615 32122
rect 4667 32070 4679 32122
rect 4731 32070 11369 32122
rect 11421 32070 11433 32122
rect 11485 32070 11497 32122
rect 11549 32070 11561 32122
rect 11613 32070 11625 32122
rect 11677 32070 18315 32122
rect 18367 32070 18379 32122
rect 18431 32070 18443 32122
rect 18495 32070 18507 32122
rect 18559 32070 18571 32122
rect 18623 32070 25261 32122
rect 25313 32070 25325 32122
rect 25377 32070 25389 32122
rect 25441 32070 25453 32122
rect 25505 32070 25517 32122
rect 25569 32070 28888 32122
rect 1104 32048 28888 32070
rect 2038 32008 2044 32020
rect 1999 31980 2044 32008
rect 2038 31968 2044 31980
rect 2096 31968 2102 32020
rect 15930 31968 15936 32020
rect 15988 32008 15994 32020
rect 16209 32011 16267 32017
rect 16209 32008 16221 32011
rect 15988 31980 16221 32008
rect 15988 31968 15994 31980
rect 16209 31977 16221 31980
rect 16255 32008 16267 32011
rect 18230 32008 18236 32020
rect 16255 31980 18236 32008
rect 16255 31977 16267 31980
rect 16209 31971 16267 31977
rect 18230 31968 18236 31980
rect 18288 31968 18294 32020
rect 19521 32011 19579 32017
rect 19521 31977 19533 32011
rect 19567 32008 19579 32011
rect 19794 32008 19800 32020
rect 19567 31980 19800 32008
rect 19567 31977 19579 31980
rect 19521 31971 19579 31977
rect 19794 31968 19800 31980
rect 19852 31968 19858 32020
rect 20898 31968 20904 32020
rect 20956 32008 20962 32020
rect 21637 32011 21695 32017
rect 21637 32008 21649 32011
rect 20956 31980 21649 32008
rect 20956 31968 20962 31980
rect 21637 31977 21649 31980
rect 21683 31977 21695 32011
rect 21637 31971 21695 31977
rect 22097 32011 22155 32017
rect 22097 31977 22109 32011
rect 22143 32008 22155 32011
rect 22278 32008 22284 32020
rect 22143 31980 22284 32008
rect 22143 31977 22155 31980
rect 22097 31971 22155 31977
rect 21652 31940 21680 31971
rect 22278 31968 22284 31980
rect 22336 31968 22342 32020
rect 23293 32011 23351 32017
rect 23293 31977 23305 32011
rect 23339 32008 23351 32011
rect 23382 32008 23388 32020
rect 23339 31980 23388 32008
rect 23339 31977 23351 31980
rect 23293 31971 23351 31977
rect 23382 31968 23388 31980
rect 23440 31968 23446 32020
rect 25593 31943 25651 31949
rect 21652 31912 23520 31940
rect 16117 31875 16175 31881
rect 16117 31841 16129 31875
rect 16163 31872 16175 31875
rect 16574 31872 16580 31884
rect 16163 31844 16580 31872
rect 16163 31841 16175 31844
rect 16117 31835 16175 31841
rect 16574 31832 16580 31844
rect 16632 31832 16638 31884
rect 16850 31832 16856 31884
rect 16908 31872 16914 31884
rect 16945 31875 17003 31881
rect 16945 31872 16957 31875
rect 16908 31844 16957 31872
rect 16908 31832 16914 31844
rect 16945 31841 16957 31844
rect 16991 31841 17003 31875
rect 16945 31835 17003 31841
rect 20993 31875 21051 31881
rect 20993 31841 21005 31875
rect 21039 31872 21051 31875
rect 22738 31872 22744 31884
rect 21039 31844 22744 31872
rect 21039 31841 21051 31844
rect 20993 31835 21051 31841
rect 22738 31832 22744 31844
rect 22796 31832 22802 31884
rect 23492 31872 23520 31912
rect 25593 31909 25605 31943
rect 25639 31940 25651 31943
rect 25866 31940 25872 31952
rect 25639 31912 25872 31940
rect 25639 31909 25651 31912
rect 25593 31903 25651 31909
rect 25866 31900 25872 31912
rect 25924 31900 25930 31952
rect 27706 31940 27712 31952
rect 26206 31912 27712 31940
rect 26206 31872 26234 31912
rect 27706 31900 27712 31912
rect 27764 31900 27770 31952
rect 26694 31872 26700 31884
rect 23492 31844 26234 31872
rect 26655 31844 26700 31872
rect 2133 31807 2191 31813
rect 2133 31773 2145 31807
rect 2179 31804 2191 31807
rect 2590 31804 2596 31816
rect 2179 31776 2596 31804
rect 2179 31773 2191 31776
rect 2133 31767 2191 31773
rect 2590 31764 2596 31776
rect 2648 31804 2654 31816
rect 4154 31804 4160 31816
rect 2648 31776 4160 31804
rect 2648 31764 2654 31776
rect 4154 31764 4160 31776
rect 4212 31764 4218 31816
rect 15286 31764 15292 31816
rect 15344 31804 15350 31816
rect 16209 31807 16267 31813
rect 16209 31804 16221 31807
rect 15344 31776 16221 31804
rect 15344 31764 15350 31776
rect 16209 31773 16221 31776
rect 16255 31773 16267 31807
rect 16209 31767 16267 31773
rect 17034 31764 17040 31816
rect 17092 31804 17098 31816
rect 17201 31807 17259 31813
rect 17201 31804 17213 31807
rect 17092 31776 17213 31804
rect 17092 31764 17098 31776
rect 17201 31773 17213 31776
rect 17247 31773 17259 31807
rect 17201 31767 17259 31773
rect 18874 31764 18880 31816
rect 18932 31804 18938 31816
rect 19429 31807 19487 31813
rect 19429 31804 19441 31807
rect 18932 31776 19441 31804
rect 18932 31764 18938 31776
rect 19429 31773 19441 31776
rect 19475 31773 19487 31807
rect 19429 31767 19487 31773
rect 20717 31807 20775 31813
rect 20717 31773 20729 31807
rect 20763 31804 20775 31807
rect 20898 31804 20904 31816
rect 20763 31776 20904 31804
rect 20763 31773 20775 31776
rect 20717 31767 20775 31773
rect 20898 31764 20904 31776
rect 20956 31764 20962 31816
rect 21542 31804 21548 31816
rect 21503 31776 21548 31804
rect 21542 31764 21548 31776
rect 21600 31764 21606 31816
rect 21634 31764 21640 31816
rect 21692 31804 21698 31816
rect 23492 31813 23520 31844
rect 26694 31832 26700 31844
rect 26752 31832 26758 31884
rect 28350 31872 28356 31884
rect 28311 31844 28356 31872
rect 28350 31832 28356 31844
rect 28408 31832 28414 31884
rect 21821 31807 21879 31813
rect 21821 31804 21833 31807
rect 21692 31776 21833 31804
rect 21692 31764 21698 31776
rect 21821 31773 21833 31776
rect 21867 31773 21879 31807
rect 21821 31767 21879 31773
rect 23477 31807 23535 31813
rect 23477 31773 23489 31807
rect 23523 31773 23535 31807
rect 23658 31804 23664 31816
rect 23619 31776 23664 31804
rect 23477 31767 23535 31773
rect 23658 31764 23664 31776
rect 23716 31764 23722 31816
rect 25130 31764 25136 31816
rect 25188 31804 25194 31816
rect 25317 31807 25375 31813
rect 25317 31804 25329 31807
rect 25188 31776 25329 31804
rect 25188 31764 25194 31776
rect 25317 31773 25329 31776
rect 25363 31773 25375 31807
rect 25317 31767 25375 31773
rect 25409 31807 25467 31813
rect 25409 31773 25421 31807
rect 25455 31804 25467 31807
rect 25455 31776 26234 31804
rect 25455 31773 25467 31776
rect 25409 31767 25467 31773
rect 25590 31736 25596 31748
rect 25551 31708 25596 31736
rect 25590 31696 25596 31708
rect 25648 31696 25654 31748
rect 15841 31671 15899 31677
rect 15841 31637 15853 31671
rect 15887 31668 15899 31671
rect 16022 31668 16028 31680
rect 15887 31640 16028 31668
rect 15887 31637 15899 31640
rect 15841 31631 15899 31637
rect 16022 31628 16028 31640
rect 16080 31628 16086 31680
rect 18322 31668 18328 31680
rect 18283 31640 18328 31668
rect 18322 31628 18328 31640
rect 18380 31628 18386 31680
rect 26206 31668 26234 31776
rect 26326 31764 26332 31816
rect 26384 31804 26390 31816
rect 26513 31807 26571 31813
rect 26513 31804 26525 31807
rect 26384 31776 26525 31804
rect 26384 31764 26390 31776
rect 26513 31773 26525 31776
rect 26559 31773 26571 31807
rect 26513 31767 26571 31773
rect 26510 31668 26516 31680
rect 26206 31640 26516 31668
rect 26510 31628 26516 31640
rect 26568 31628 26574 31680
rect 1104 31578 29048 31600
rect 1104 31526 7896 31578
rect 7948 31526 7960 31578
rect 8012 31526 8024 31578
rect 8076 31526 8088 31578
rect 8140 31526 8152 31578
rect 8204 31526 14842 31578
rect 14894 31526 14906 31578
rect 14958 31526 14970 31578
rect 15022 31526 15034 31578
rect 15086 31526 15098 31578
rect 15150 31526 21788 31578
rect 21840 31526 21852 31578
rect 21904 31526 21916 31578
rect 21968 31526 21980 31578
rect 22032 31526 22044 31578
rect 22096 31526 28734 31578
rect 28786 31526 28798 31578
rect 28850 31526 28862 31578
rect 28914 31526 28926 31578
rect 28978 31526 28990 31578
rect 29042 31526 29048 31578
rect 1104 31504 29048 31526
rect 18230 31424 18236 31476
rect 18288 31464 18294 31476
rect 18417 31467 18475 31473
rect 18417 31464 18429 31467
rect 18288 31436 18429 31464
rect 18288 31424 18294 31436
rect 18417 31433 18429 31436
rect 18463 31433 18475 31467
rect 22646 31464 22652 31476
rect 22607 31436 22652 31464
rect 18417 31427 18475 31433
rect 22646 31424 22652 31436
rect 22704 31424 22710 31476
rect 24305 31467 24363 31473
rect 24305 31433 24317 31467
rect 24351 31464 24363 31467
rect 25038 31464 25044 31476
rect 24351 31436 25044 31464
rect 24351 31433 24363 31436
rect 24305 31427 24363 31433
rect 25038 31424 25044 31436
rect 25096 31424 25102 31476
rect 25590 31356 25596 31408
rect 25648 31396 25654 31408
rect 25648 31368 27568 31396
rect 25648 31356 25654 31368
rect 15838 31328 15844 31340
rect 15799 31300 15844 31328
rect 15838 31288 15844 31300
rect 15896 31288 15902 31340
rect 16025 31331 16083 31337
rect 16025 31297 16037 31331
rect 16071 31328 16083 31331
rect 16574 31328 16580 31340
rect 16071 31300 16580 31328
rect 16071 31297 16083 31300
rect 16025 31291 16083 31297
rect 16574 31288 16580 31300
rect 16632 31328 16638 31340
rect 17862 31328 17868 31340
rect 16632 31300 17868 31328
rect 16632 31288 16638 31300
rect 17862 31288 17868 31300
rect 17920 31288 17926 31340
rect 18322 31328 18328 31340
rect 18283 31300 18328 31328
rect 18322 31288 18328 31300
rect 18380 31288 18386 31340
rect 22557 31331 22615 31337
rect 22557 31297 22569 31331
rect 22603 31328 22615 31331
rect 22646 31328 22652 31340
rect 22603 31300 22652 31328
rect 22603 31297 22615 31300
rect 22557 31291 22615 31297
rect 22646 31288 22652 31300
rect 22704 31288 22710 31340
rect 22741 31331 22799 31337
rect 22741 31297 22753 31331
rect 22787 31297 22799 31331
rect 22741 31291 22799 31297
rect 22756 31260 22784 31291
rect 23474 31288 23480 31340
rect 23532 31328 23538 31340
rect 24213 31331 24271 31337
rect 24213 31328 24225 31331
rect 23532 31300 24225 31328
rect 23532 31288 23538 31300
rect 24213 31297 24225 31300
rect 24259 31297 24271 31331
rect 24394 31328 24400 31340
rect 24355 31300 24400 31328
rect 24213 31291 24271 31297
rect 24394 31288 24400 31300
rect 24452 31288 24458 31340
rect 26050 31288 26056 31340
rect 26108 31328 26114 31340
rect 26338 31331 26396 31337
rect 26338 31328 26350 31331
rect 26108 31300 26350 31328
rect 26108 31288 26114 31300
rect 26338 31297 26350 31300
rect 26384 31297 26396 31331
rect 26338 31291 26396 31297
rect 26510 31288 26516 31340
rect 26568 31328 26574 31340
rect 27540 31337 27568 31368
rect 27433 31331 27491 31337
rect 27433 31328 27445 31331
rect 26568 31300 27445 31328
rect 26568 31288 26574 31300
rect 27433 31297 27445 31300
rect 27479 31297 27491 31331
rect 27433 31291 27491 31297
rect 27525 31331 27583 31337
rect 27525 31297 27537 31331
rect 27571 31297 27583 31331
rect 27525 31291 27583 31297
rect 27617 31331 27675 31337
rect 27617 31297 27629 31331
rect 27663 31328 27675 31331
rect 27706 31328 27712 31340
rect 27663 31300 27712 31328
rect 27663 31297 27675 31300
rect 27617 31291 27675 31297
rect 27706 31288 27712 31300
rect 27764 31288 27770 31340
rect 28169 31331 28227 31337
rect 28169 31297 28181 31331
rect 28215 31328 28227 31331
rect 28350 31328 28356 31340
rect 28215 31300 28356 31328
rect 28215 31297 28227 31300
rect 28169 31291 28227 31297
rect 28350 31288 28356 31300
rect 28408 31288 28414 31340
rect 24486 31260 24492 31272
rect 22756 31232 24492 31260
rect 24486 31220 24492 31232
rect 24544 31220 24550 31272
rect 26605 31263 26663 31269
rect 26605 31229 26617 31263
rect 26651 31229 26663 31263
rect 27338 31260 27344 31272
rect 27299 31232 27344 31260
rect 26605 31223 26663 31229
rect 15930 31124 15936 31136
rect 15891 31096 15936 31124
rect 15930 31084 15936 31096
rect 15988 31084 15994 31136
rect 25225 31127 25283 31133
rect 25225 31093 25237 31127
rect 25271 31124 25283 31127
rect 25590 31124 25596 31136
rect 25271 31096 25596 31124
rect 25271 31093 25283 31096
rect 25225 31087 25283 31093
rect 25590 31084 25596 31096
rect 25648 31084 25654 31136
rect 25958 31084 25964 31136
rect 26016 31124 26022 31136
rect 26620 31124 26648 31223
rect 27338 31220 27344 31232
rect 27396 31220 27402 31272
rect 26016 31096 26648 31124
rect 26016 31084 26022 31096
rect 26694 31084 26700 31136
rect 26752 31124 26758 31136
rect 27157 31127 27215 31133
rect 27157 31124 27169 31127
rect 26752 31096 27169 31124
rect 26752 31084 26758 31096
rect 27157 31093 27169 31096
rect 27203 31093 27215 31127
rect 27157 31087 27215 31093
rect 28166 31084 28172 31136
rect 28224 31124 28230 31136
rect 28261 31127 28319 31133
rect 28261 31124 28273 31127
rect 28224 31096 28273 31124
rect 28224 31084 28230 31096
rect 28261 31093 28273 31096
rect 28307 31093 28319 31127
rect 28261 31087 28319 31093
rect 1104 31034 28888 31056
rect 1104 30982 4423 31034
rect 4475 30982 4487 31034
rect 4539 30982 4551 31034
rect 4603 30982 4615 31034
rect 4667 30982 4679 31034
rect 4731 30982 11369 31034
rect 11421 30982 11433 31034
rect 11485 30982 11497 31034
rect 11549 30982 11561 31034
rect 11613 30982 11625 31034
rect 11677 30982 18315 31034
rect 18367 30982 18379 31034
rect 18431 30982 18443 31034
rect 18495 30982 18507 31034
rect 18559 30982 18571 31034
rect 18623 30982 25261 31034
rect 25313 30982 25325 31034
rect 25377 30982 25389 31034
rect 25441 30982 25453 31034
rect 25505 30982 25517 31034
rect 25569 30982 28888 31034
rect 1104 30960 28888 30982
rect 16022 30920 16028 30932
rect 15983 30892 16028 30920
rect 16022 30880 16028 30892
rect 16080 30880 16086 30932
rect 17862 30920 17868 30932
rect 17823 30892 17868 30920
rect 17862 30880 17868 30892
rect 17920 30880 17926 30932
rect 25130 30880 25136 30932
rect 25188 30920 25194 30932
rect 25409 30923 25467 30929
rect 25409 30920 25421 30923
rect 25188 30892 25421 30920
rect 25188 30880 25194 30892
rect 25409 30889 25421 30892
rect 25455 30889 25467 30923
rect 26050 30920 26056 30932
rect 26011 30892 26056 30920
rect 25409 30883 25467 30889
rect 26050 30880 26056 30892
rect 26108 30880 26114 30932
rect 28350 30920 28356 30932
rect 26160 30892 28356 30920
rect 2130 30812 2136 30864
rect 2188 30852 2194 30864
rect 26160 30852 26188 30892
rect 28350 30880 28356 30892
rect 28408 30880 28414 30932
rect 2188 30824 26188 30852
rect 2188 30812 2194 30824
rect 28258 30812 28264 30864
rect 28316 30812 28322 30864
rect 8481 30787 8539 30793
rect 8481 30753 8493 30787
rect 8527 30784 8539 30787
rect 10781 30787 10839 30793
rect 10781 30784 10793 30787
rect 8527 30756 10793 30784
rect 8527 30753 8539 30756
rect 8481 30747 8539 30753
rect 10781 30753 10793 30756
rect 10827 30753 10839 30787
rect 27430 30784 27436 30796
rect 27391 30756 27436 30784
rect 10781 30747 10839 30753
rect 27430 30744 27436 30756
rect 27488 30744 27494 30796
rect 28166 30784 28172 30796
rect 28127 30756 28172 30784
rect 28166 30744 28172 30756
rect 28224 30744 28230 30796
rect 28276 30784 28304 30812
rect 28353 30787 28411 30793
rect 28353 30784 28365 30787
rect 28276 30756 28365 30784
rect 28353 30753 28365 30756
rect 28399 30753 28411 30787
rect 28353 30747 28411 30753
rect 8389 30719 8447 30725
rect 8389 30685 8401 30719
rect 8435 30685 8447 30719
rect 9122 30716 9128 30728
rect 9083 30688 9128 30716
rect 8389 30679 8447 30685
rect 8404 30648 8432 30679
rect 9122 30676 9128 30688
rect 9180 30676 9186 30728
rect 10965 30719 11023 30725
rect 10965 30685 10977 30719
rect 11011 30716 11023 30719
rect 12618 30716 12624 30728
rect 11011 30688 12624 30716
rect 11011 30685 11023 30688
rect 10965 30679 11023 30685
rect 12618 30676 12624 30688
rect 12676 30676 12682 30728
rect 17954 30716 17960 30728
rect 17915 30688 17960 30716
rect 17954 30676 17960 30688
rect 18012 30676 18018 30728
rect 24854 30716 24860 30728
rect 24815 30688 24860 30716
rect 24854 30676 24860 30688
rect 24912 30676 24918 30728
rect 25038 30716 25044 30728
rect 24999 30688 25044 30716
rect 25038 30676 25044 30688
rect 25096 30676 25102 30728
rect 25225 30719 25283 30725
rect 25225 30685 25237 30719
rect 25271 30685 25283 30719
rect 25866 30716 25872 30728
rect 25827 30688 25872 30716
rect 25225 30679 25283 30685
rect 9582 30648 9588 30660
rect 8404 30620 9588 30648
rect 9582 30608 9588 30620
rect 9640 30648 9646 30660
rect 9950 30648 9956 30660
rect 9640 30620 9956 30648
rect 9640 30608 9646 30620
rect 9950 30608 9956 30620
rect 10008 30608 10014 30660
rect 15838 30648 15844 30660
rect 15799 30620 15844 30648
rect 15838 30608 15844 30620
rect 15896 30608 15902 30660
rect 15930 30608 15936 30660
rect 15988 30648 15994 30660
rect 16041 30651 16099 30657
rect 16041 30648 16053 30651
rect 15988 30620 16053 30648
rect 15988 30608 15994 30620
rect 16041 30617 16053 30620
rect 16087 30617 16099 30651
rect 22554 30648 22560 30660
rect 22515 30620 22560 30648
rect 16041 30611 16099 30617
rect 22554 30608 22560 30620
rect 22612 30608 22618 30660
rect 24394 30608 24400 30660
rect 24452 30648 24458 30660
rect 25133 30651 25191 30657
rect 25133 30648 25145 30651
rect 24452 30620 25145 30648
rect 24452 30608 24458 30620
rect 25133 30617 25145 30620
rect 25179 30617 25191 30651
rect 25240 30648 25268 30679
rect 25866 30676 25872 30688
rect 25924 30676 25930 30728
rect 26053 30719 26111 30725
rect 26053 30685 26065 30719
rect 26099 30716 26111 30719
rect 26694 30716 26700 30728
rect 26099 30688 26700 30716
rect 26099 30685 26111 30688
rect 26053 30679 26111 30685
rect 26694 30676 26700 30688
rect 26752 30676 26758 30728
rect 25774 30648 25780 30660
rect 25240 30620 25780 30648
rect 25133 30611 25191 30617
rect 25774 30608 25780 30620
rect 25832 30608 25838 30660
rect 16206 30580 16212 30592
rect 16167 30552 16212 30580
rect 16206 30540 16212 30552
rect 16264 30540 16270 30592
rect 21269 30583 21327 30589
rect 21269 30549 21281 30583
rect 21315 30580 21327 30583
rect 22186 30580 22192 30592
rect 21315 30552 22192 30580
rect 21315 30549 21327 30552
rect 21269 30543 21327 30549
rect 22186 30540 22192 30552
rect 22244 30540 22250 30592
rect 1104 30490 29048 30512
rect 1104 30438 7896 30490
rect 7948 30438 7960 30490
rect 8012 30438 8024 30490
rect 8076 30438 8088 30490
rect 8140 30438 8152 30490
rect 8204 30438 14842 30490
rect 14894 30438 14906 30490
rect 14958 30438 14970 30490
rect 15022 30438 15034 30490
rect 15086 30438 15098 30490
rect 15150 30438 21788 30490
rect 21840 30438 21852 30490
rect 21904 30438 21916 30490
rect 21968 30438 21980 30490
rect 22032 30438 22044 30490
rect 22096 30438 28734 30490
rect 28786 30438 28798 30490
rect 28850 30438 28862 30490
rect 28914 30438 28926 30490
rect 28978 30438 28990 30490
rect 29042 30438 29048 30490
rect 1104 30416 29048 30438
rect 17954 30336 17960 30388
rect 18012 30376 18018 30388
rect 18233 30379 18291 30385
rect 18233 30376 18245 30379
rect 18012 30348 18245 30376
rect 18012 30336 18018 30348
rect 18233 30345 18245 30348
rect 18279 30345 18291 30379
rect 18233 30339 18291 30345
rect 19889 30311 19947 30317
rect 19889 30277 19901 30311
rect 19935 30308 19947 30311
rect 20530 30308 20536 30320
rect 19935 30280 20536 30308
rect 19935 30277 19947 30280
rect 19889 30271 19947 30277
rect 20530 30268 20536 30280
rect 20588 30268 20594 30320
rect 21174 30308 21180 30320
rect 20824 30280 21180 30308
rect 1578 30240 1584 30252
rect 1539 30212 1584 30240
rect 1578 30200 1584 30212
rect 1636 30200 1642 30252
rect 16117 30243 16175 30249
rect 16117 30209 16129 30243
rect 16163 30240 16175 30243
rect 16206 30240 16212 30252
rect 16163 30212 16212 30240
rect 16163 30209 16175 30212
rect 16117 30203 16175 30209
rect 16206 30200 16212 30212
rect 16264 30200 16270 30252
rect 16850 30240 16856 30252
rect 16811 30212 16856 30240
rect 16850 30200 16856 30212
rect 16908 30200 16914 30252
rect 20824 30249 20852 30280
rect 21174 30268 21180 30280
rect 21232 30308 21238 30320
rect 22646 30308 22652 30320
rect 21232 30280 22652 30308
rect 21232 30268 21238 30280
rect 22646 30268 22652 30280
rect 22704 30268 22710 30320
rect 17109 30243 17167 30249
rect 17109 30240 17121 30243
rect 16960 30212 17121 30240
rect 16960 30172 16988 30212
rect 17109 30209 17121 30212
rect 17155 30209 17167 30243
rect 17109 30203 17167 30209
rect 19981 30243 20039 30249
rect 19981 30209 19993 30243
rect 20027 30240 20039 30243
rect 20809 30243 20867 30249
rect 20027 30212 20760 30240
rect 20027 30209 20039 30212
rect 19981 30203 20039 30209
rect 20162 30172 20168 30184
rect 16316 30144 16988 30172
rect 20123 30144 20168 30172
rect 16316 30113 16344 30144
rect 20162 30132 20168 30144
rect 20220 30132 20226 30184
rect 20732 30172 20760 30212
rect 20809 30209 20821 30243
rect 20855 30209 20867 30243
rect 20990 30240 20996 30252
rect 20951 30212 20996 30240
rect 20809 30203 20867 30209
rect 20990 30200 20996 30212
rect 21048 30200 21054 30252
rect 26602 30240 26608 30252
rect 26563 30212 26608 30240
rect 26602 30200 26608 30212
rect 26660 30200 26666 30252
rect 22370 30172 22376 30184
rect 20732 30144 22376 30172
rect 22370 30132 22376 30144
rect 22428 30172 22434 30184
rect 24578 30172 24584 30184
rect 22428 30144 24584 30172
rect 22428 30132 22434 30144
rect 24578 30132 24584 30144
rect 24636 30132 24642 30184
rect 16301 30107 16359 30113
rect 16301 30073 16313 30107
rect 16347 30073 16359 30107
rect 26418 30104 26424 30116
rect 26379 30076 26424 30104
rect 16301 30067 16359 30073
rect 26418 30064 26424 30076
rect 26476 30064 26482 30116
rect 1765 30039 1823 30045
rect 1765 30005 1777 30039
rect 1811 30036 1823 30039
rect 1854 30036 1860 30048
rect 1811 30008 1860 30036
rect 1811 30005 1823 30008
rect 1765 29999 1823 30005
rect 1854 29996 1860 30008
rect 1912 29996 1918 30048
rect 19521 30039 19579 30045
rect 19521 30005 19533 30039
rect 19567 30036 19579 30039
rect 19610 30036 19616 30048
rect 19567 30008 19616 30036
rect 19567 30005 19579 30008
rect 19521 29999 19579 30005
rect 19610 29996 19616 30008
rect 19668 29996 19674 30048
rect 20806 29996 20812 30048
rect 20864 30036 20870 30048
rect 20993 30039 21051 30045
rect 20993 30036 21005 30039
rect 20864 30008 21005 30036
rect 20864 29996 20870 30008
rect 20993 30005 21005 30008
rect 21039 30005 21051 30039
rect 20993 29999 21051 30005
rect 27893 30039 27951 30045
rect 27893 30005 27905 30039
rect 27939 30036 27951 30039
rect 28350 30036 28356 30048
rect 27939 30008 28356 30036
rect 27939 30005 27951 30008
rect 27893 29999 27951 30005
rect 28350 29996 28356 30008
rect 28408 29996 28414 30048
rect 1104 29946 28888 29968
rect 1104 29894 4423 29946
rect 4475 29894 4487 29946
rect 4539 29894 4551 29946
rect 4603 29894 4615 29946
rect 4667 29894 4679 29946
rect 4731 29894 11369 29946
rect 11421 29894 11433 29946
rect 11485 29894 11497 29946
rect 11549 29894 11561 29946
rect 11613 29894 11625 29946
rect 11677 29894 18315 29946
rect 18367 29894 18379 29946
rect 18431 29894 18443 29946
rect 18495 29894 18507 29946
rect 18559 29894 18571 29946
rect 18623 29894 25261 29946
rect 25313 29894 25325 29946
rect 25377 29894 25389 29946
rect 25441 29894 25453 29946
rect 25505 29894 25517 29946
rect 25569 29894 28888 29946
rect 1104 29872 28888 29894
rect 16758 29792 16764 29844
rect 16816 29832 16822 29844
rect 17681 29835 17739 29841
rect 17681 29832 17693 29835
rect 16816 29804 17693 29832
rect 16816 29792 16822 29804
rect 17681 29801 17693 29804
rect 17727 29801 17739 29835
rect 17681 29795 17739 29801
rect 18230 29792 18236 29844
rect 18288 29832 18294 29844
rect 18325 29835 18383 29841
rect 18325 29832 18337 29835
rect 18288 29804 18337 29832
rect 18288 29792 18294 29804
rect 18325 29801 18337 29804
rect 18371 29801 18383 29835
rect 18325 29795 18383 29801
rect 18693 29835 18751 29841
rect 18693 29801 18705 29835
rect 18739 29832 18751 29835
rect 18782 29832 18788 29844
rect 18739 29804 18788 29832
rect 18739 29801 18751 29804
rect 18693 29795 18751 29801
rect 18782 29792 18788 29804
rect 18840 29792 18846 29844
rect 25133 29835 25191 29841
rect 25133 29801 25145 29835
rect 25179 29832 25191 29835
rect 25590 29832 25596 29844
rect 25179 29804 25596 29832
rect 25179 29801 25191 29804
rect 25133 29795 25191 29801
rect 25590 29792 25596 29804
rect 25648 29832 25654 29844
rect 26050 29832 26056 29844
rect 25648 29804 26056 29832
rect 25648 29792 25654 29804
rect 26050 29792 26056 29804
rect 26108 29792 26114 29844
rect 16666 29696 16672 29708
rect 16040 29668 16672 29696
rect 15841 29631 15899 29637
rect 15841 29597 15853 29631
rect 15887 29628 15899 29631
rect 15930 29628 15936 29640
rect 15887 29600 15936 29628
rect 15887 29597 15899 29600
rect 15841 29591 15899 29597
rect 15930 29588 15936 29600
rect 15988 29588 15994 29640
rect 16040 29637 16068 29668
rect 16666 29656 16672 29668
rect 16724 29696 16730 29708
rect 16776 29696 16804 29792
rect 23385 29767 23443 29773
rect 23385 29733 23397 29767
rect 23431 29733 23443 29767
rect 23385 29727 23443 29733
rect 16724 29668 16804 29696
rect 16724 29656 16730 29668
rect 18046 29656 18052 29708
rect 18104 29696 18110 29708
rect 18104 29668 18276 29696
rect 18104 29656 18110 29668
rect 16025 29631 16083 29637
rect 16025 29597 16037 29631
rect 16071 29597 16083 29631
rect 16574 29628 16580 29640
rect 16535 29600 16580 29628
rect 16025 29591 16083 29597
rect 16574 29588 16580 29600
rect 16632 29588 16638 29640
rect 17773 29631 17831 29637
rect 17773 29597 17785 29631
rect 17819 29628 17831 29631
rect 18138 29628 18144 29640
rect 17819 29600 18144 29628
rect 17819 29597 17831 29600
rect 17773 29591 17831 29597
rect 18138 29588 18144 29600
rect 18196 29588 18202 29640
rect 18248 29637 18276 29668
rect 19518 29656 19524 29708
rect 19576 29696 19582 29708
rect 20533 29699 20591 29705
rect 20533 29696 20545 29699
rect 19576 29668 20545 29696
rect 19576 29656 19582 29668
rect 20533 29665 20545 29668
rect 20579 29665 20591 29699
rect 20806 29696 20812 29708
rect 20767 29668 20812 29696
rect 20533 29659 20591 29665
rect 20806 29656 20812 29668
rect 20864 29656 20870 29708
rect 22646 29696 22652 29708
rect 22607 29668 22652 29696
rect 22646 29656 22652 29668
rect 22704 29656 22710 29708
rect 18233 29631 18291 29637
rect 18233 29597 18245 29631
rect 18279 29597 18291 29631
rect 18233 29591 18291 29597
rect 19429 29631 19487 29637
rect 19429 29597 19441 29631
rect 19475 29597 19487 29631
rect 19610 29628 19616 29640
rect 19571 29600 19616 29628
rect 19429 29591 19487 29597
rect 19444 29560 19472 29591
rect 19610 29588 19616 29600
rect 19668 29588 19674 29640
rect 21174 29628 21180 29640
rect 19720 29600 21180 29628
rect 19720 29560 19748 29600
rect 21174 29588 21180 29600
rect 21232 29588 21238 29640
rect 22830 29628 22836 29640
rect 22791 29600 22836 29628
rect 22830 29588 22836 29600
rect 22888 29588 22894 29640
rect 22925 29631 22983 29637
rect 22925 29597 22937 29631
rect 22971 29628 22983 29631
rect 23400 29628 23428 29727
rect 27522 29696 27528 29708
rect 27483 29668 27528 29696
rect 27522 29656 27528 29668
rect 27580 29656 27586 29708
rect 28350 29696 28356 29708
rect 28311 29668 28356 29696
rect 28350 29656 28356 29668
rect 28408 29656 28414 29708
rect 22971 29600 23428 29628
rect 23661 29631 23719 29637
rect 22971 29597 22983 29600
rect 22925 29591 22983 29597
rect 23661 29597 23673 29631
rect 23707 29628 23719 29631
rect 23934 29628 23940 29640
rect 23707 29600 23940 29628
rect 23707 29597 23719 29600
rect 23661 29591 23719 29597
rect 23934 29588 23940 29600
rect 23992 29588 23998 29640
rect 19444 29532 19748 29560
rect 23385 29563 23443 29569
rect 23385 29529 23397 29563
rect 23431 29560 23443 29563
rect 23474 29560 23480 29572
rect 23431 29532 23480 29560
rect 23431 29529 23443 29532
rect 23385 29523 23443 29529
rect 23474 29520 23480 29532
rect 23532 29520 23538 29572
rect 24854 29520 24860 29572
rect 24912 29560 24918 29572
rect 25317 29563 25375 29569
rect 24912 29532 25084 29560
rect 24912 29520 24918 29532
rect 15746 29452 15752 29504
rect 15804 29492 15810 29504
rect 15933 29495 15991 29501
rect 15933 29492 15945 29495
rect 15804 29464 15945 29492
rect 15804 29452 15810 29464
rect 15933 29461 15945 29464
rect 15979 29461 15991 29495
rect 16758 29492 16764 29504
rect 16719 29464 16764 29492
rect 15933 29455 15991 29461
rect 16758 29452 16764 29464
rect 16816 29452 16822 29504
rect 19518 29492 19524 29504
rect 19479 29464 19524 29492
rect 19518 29452 19524 29464
rect 19576 29452 19582 29504
rect 20898 29452 20904 29504
rect 20956 29492 20962 29504
rect 21913 29495 21971 29501
rect 21913 29492 21925 29495
rect 20956 29464 21925 29492
rect 20956 29452 20962 29464
rect 21913 29461 21925 29464
rect 21959 29461 21971 29495
rect 22922 29492 22928 29504
rect 22883 29464 22928 29492
rect 21913 29455 21971 29461
rect 22922 29452 22928 29464
rect 22980 29452 22986 29504
rect 23569 29495 23627 29501
rect 23569 29461 23581 29495
rect 23615 29492 23627 29495
rect 24946 29492 24952 29504
rect 23615 29464 24952 29492
rect 23615 29461 23627 29464
rect 23569 29455 23627 29461
rect 24946 29452 24952 29464
rect 25004 29452 25010 29504
rect 25056 29492 25084 29532
rect 25317 29529 25329 29563
rect 25363 29560 25375 29563
rect 26142 29560 26148 29572
rect 25363 29532 26148 29560
rect 25363 29529 25375 29532
rect 25317 29523 25375 29529
rect 26142 29520 26148 29532
rect 26200 29520 26206 29572
rect 27706 29520 27712 29572
rect 27764 29560 27770 29572
rect 28169 29563 28227 29569
rect 28169 29560 28181 29563
rect 27764 29532 28181 29560
rect 27764 29520 27770 29532
rect 28169 29529 28181 29532
rect 28215 29529 28227 29563
rect 28169 29523 28227 29529
rect 25117 29495 25175 29501
rect 25117 29492 25129 29495
rect 25056 29464 25129 29492
rect 25117 29461 25129 29464
rect 25163 29492 25175 29495
rect 25866 29492 25872 29504
rect 25163 29464 25872 29492
rect 25163 29461 25175 29464
rect 25117 29455 25175 29461
rect 25866 29452 25872 29464
rect 25924 29452 25930 29504
rect 1104 29402 29048 29424
rect 1104 29350 7896 29402
rect 7948 29350 7960 29402
rect 8012 29350 8024 29402
rect 8076 29350 8088 29402
rect 8140 29350 8152 29402
rect 8204 29350 14842 29402
rect 14894 29350 14906 29402
rect 14958 29350 14970 29402
rect 15022 29350 15034 29402
rect 15086 29350 15098 29402
rect 15150 29350 21788 29402
rect 21840 29350 21852 29402
rect 21904 29350 21916 29402
rect 21968 29350 21980 29402
rect 22032 29350 22044 29402
rect 22096 29350 28734 29402
rect 28786 29350 28798 29402
rect 28850 29350 28862 29402
rect 28914 29350 28926 29402
rect 28978 29350 28990 29402
rect 29042 29350 29048 29402
rect 1104 29328 29048 29350
rect 20990 29248 20996 29300
rect 21048 29288 21054 29300
rect 21170 29291 21228 29297
rect 21170 29288 21182 29291
rect 21048 29260 21182 29288
rect 21048 29248 21054 29260
rect 21170 29257 21182 29260
rect 21216 29257 21228 29291
rect 21170 29251 21228 29257
rect 22830 29248 22836 29300
rect 22888 29288 22894 29300
rect 23937 29291 23995 29297
rect 23937 29288 23949 29291
rect 22888 29260 23949 29288
rect 22888 29248 22894 29260
rect 23937 29257 23949 29260
rect 23983 29257 23995 29291
rect 27706 29288 27712 29300
rect 27667 29260 27712 29288
rect 23937 29251 23995 29257
rect 27706 29248 27712 29260
rect 27764 29248 27770 29300
rect 19981 29223 20039 29229
rect 19981 29189 19993 29223
rect 20027 29220 20039 29223
rect 22554 29220 22560 29232
rect 20027 29192 22560 29220
rect 20027 29189 20039 29192
rect 19981 29183 20039 29189
rect 22554 29180 22560 29192
rect 22612 29180 22618 29232
rect 24320 29192 24808 29220
rect 15841 29155 15899 29161
rect 15841 29121 15853 29155
rect 15887 29152 15899 29155
rect 15930 29152 15936 29164
rect 15887 29124 15936 29152
rect 15887 29121 15899 29124
rect 15841 29115 15899 29121
rect 15930 29112 15936 29124
rect 15988 29112 15994 29164
rect 16025 29155 16083 29161
rect 16025 29121 16037 29155
rect 16071 29152 16083 29155
rect 16666 29152 16672 29164
rect 16071 29124 16672 29152
rect 16071 29121 16083 29124
rect 16025 29115 16083 29121
rect 16666 29112 16672 29124
rect 16724 29112 16730 29164
rect 20898 29112 20904 29164
rect 20956 29152 20962 29164
rect 20993 29155 21051 29161
rect 20993 29152 21005 29155
rect 20956 29124 21005 29152
rect 20956 29112 20962 29124
rect 20993 29121 21005 29124
rect 21039 29121 21051 29155
rect 20993 29115 21051 29121
rect 21082 29112 21088 29164
rect 21140 29152 21146 29164
rect 21269 29155 21327 29161
rect 21140 29124 21185 29152
rect 21140 29112 21146 29124
rect 21269 29121 21281 29155
rect 21315 29152 21327 29155
rect 21315 29124 21680 29152
rect 21315 29121 21327 29124
rect 21269 29115 21327 29121
rect 21652 29096 21680 29124
rect 22094 29112 22100 29164
rect 22152 29152 22158 29164
rect 22364 29155 22422 29161
rect 22152 29124 22197 29152
rect 22152 29112 22158 29124
rect 22364 29121 22376 29155
rect 22410 29152 22422 29155
rect 22922 29152 22928 29164
rect 22410 29124 22928 29152
rect 22410 29121 22422 29124
rect 22364 29115 22422 29121
rect 22922 29112 22928 29124
rect 22980 29112 22986 29164
rect 23474 29112 23480 29164
rect 23532 29152 23538 29164
rect 24320 29161 24348 29192
rect 24213 29155 24271 29161
rect 24213 29152 24225 29155
rect 23532 29124 24225 29152
rect 23532 29112 23538 29124
rect 24213 29121 24225 29124
rect 24259 29121 24271 29155
rect 24213 29115 24271 29121
rect 24305 29155 24363 29161
rect 24305 29121 24317 29155
rect 24351 29121 24363 29155
rect 24305 29115 24363 29121
rect 24397 29155 24455 29161
rect 24397 29121 24409 29155
rect 24443 29121 24455 29155
rect 24578 29152 24584 29164
rect 24539 29124 24584 29152
rect 24397 29115 24455 29121
rect 16850 29044 16856 29096
rect 16908 29084 16914 29096
rect 18233 29087 18291 29093
rect 18233 29084 18245 29087
rect 16908 29056 18245 29084
rect 16908 29044 16914 29056
rect 18233 29053 18245 29056
rect 18279 29084 18291 29087
rect 19426 29084 19432 29096
rect 18279 29056 19432 29084
rect 18279 29053 18291 29056
rect 18233 29047 18291 29053
rect 19426 29044 19432 29056
rect 19484 29044 19490 29096
rect 21634 29044 21640 29096
rect 21692 29084 21698 29096
rect 21692 29056 22094 29084
rect 21692 29044 21698 29056
rect 22066 29016 22094 29056
rect 24026 29044 24032 29096
rect 24084 29084 24090 29096
rect 24320 29084 24348 29115
rect 24084 29056 24348 29084
rect 24412 29084 24440 29115
rect 24578 29112 24584 29124
rect 24636 29112 24642 29164
rect 24780 29152 24808 29192
rect 24946 29180 24952 29232
rect 25004 29220 25010 29232
rect 25409 29223 25467 29229
rect 25409 29220 25421 29223
rect 25004 29192 25421 29220
rect 25004 29180 25010 29192
rect 25409 29189 25421 29192
rect 25455 29189 25467 29223
rect 26142 29220 26148 29232
rect 26103 29192 26148 29220
rect 25409 29183 25467 29189
rect 26142 29180 26148 29192
rect 26200 29180 26206 29232
rect 25225 29155 25283 29161
rect 25225 29152 25237 29155
rect 24780 29124 25237 29152
rect 25225 29121 25237 29124
rect 25271 29121 25283 29155
rect 25866 29152 25872 29164
rect 25827 29124 25872 29152
rect 25225 29115 25283 29121
rect 25866 29112 25872 29124
rect 25924 29112 25930 29164
rect 25961 29155 26019 29161
rect 25961 29121 25973 29155
rect 26007 29152 26019 29155
rect 26050 29152 26056 29164
rect 26007 29124 26056 29152
rect 26007 29121 26019 29124
rect 25961 29115 26019 29121
rect 26050 29112 26056 29124
rect 26108 29152 26114 29164
rect 27617 29155 27675 29161
rect 26108 29124 26201 29152
rect 26108 29112 26114 29124
rect 25041 29087 25099 29093
rect 25041 29084 25053 29087
rect 24412 29056 25053 29084
rect 24084 29044 24090 29056
rect 25041 29053 25053 29056
rect 25087 29084 25099 29087
rect 25130 29084 25136 29096
rect 25087 29056 25136 29084
rect 25087 29053 25099 29056
rect 25041 29047 25099 29053
rect 25130 29044 25136 29056
rect 25188 29044 25194 29096
rect 23474 29016 23480 29028
rect 22066 28988 22140 29016
rect 23435 28988 23480 29016
rect 15930 28948 15936 28960
rect 15891 28920 15936 28948
rect 15930 28908 15936 28920
rect 15988 28908 15994 28960
rect 22112 28948 22140 28988
rect 23474 28976 23480 28988
rect 23532 28976 23538 29028
rect 26160 29016 26188 29124
rect 27617 29121 27629 29155
rect 27663 29152 27675 29155
rect 27890 29152 27896 29164
rect 27663 29124 27896 29152
rect 27663 29121 27675 29124
rect 27617 29115 27675 29121
rect 27890 29112 27896 29124
rect 27948 29112 27954 29164
rect 26160 28988 26280 29016
rect 26252 28960 26280 28988
rect 22278 28948 22284 28960
rect 22112 28920 22284 28948
rect 22278 28908 22284 28920
rect 22336 28908 22342 28960
rect 25590 28908 25596 28960
rect 25648 28948 25654 28960
rect 26145 28951 26203 28957
rect 26145 28948 26157 28951
rect 25648 28920 26157 28948
rect 25648 28908 25654 28920
rect 26145 28917 26157 28920
rect 26191 28917 26203 28951
rect 26145 28911 26203 28917
rect 26234 28908 26240 28960
rect 26292 28908 26298 28960
rect 1104 28858 28888 28880
rect 1104 28806 4423 28858
rect 4475 28806 4487 28858
rect 4539 28806 4551 28858
rect 4603 28806 4615 28858
rect 4667 28806 4679 28858
rect 4731 28806 11369 28858
rect 11421 28806 11433 28858
rect 11485 28806 11497 28858
rect 11549 28806 11561 28858
rect 11613 28806 11625 28858
rect 11677 28806 18315 28858
rect 18367 28806 18379 28858
rect 18431 28806 18443 28858
rect 18495 28806 18507 28858
rect 18559 28806 18571 28858
rect 18623 28806 25261 28858
rect 25313 28806 25325 28858
rect 25377 28806 25389 28858
rect 25441 28806 25453 28858
rect 25505 28806 25517 28858
rect 25569 28806 28888 28858
rect 1104 28784 28888 28806
rect 15838 28704 15844 28756
rect 15896 28744 15902 28756
rect 16117 28747 16175 28753
rect 16117 28744 16129 28747
rect 15896 28716 16129 28744
rect 15896 28704 15902 28716
rect 16117 28713 16129 28716
rect 16163 28713 16175 28747
rect 16117 28707 16175 28713
rect 16301 28747 16359 28753
rect 16301 28713 16313 28747
rect 16347 28744 16359 28747
rect 16574 28744 16580 28756
rect 16347 28716 16580 28744
rect 16347 28713 16359 28716
rect 16301 28707 16359 28713
rect 16132 28676 16160 28707
rect 16574 28704 16580 28716
rect 16632 28704 16638 28756
rect 18230 28744 18236 28756
rect 18191 28716 18236 28744
rect 18230 28704 18236 28716
rect 18288 28704 18294 28756
rect 20162 28704 20168 28756
rect 20220 28744 20226 28756
rect 20809 28747 20867 28753
rect 20809 28744 20821 28747
rect 20220 28716 20821 28744
rect 20220 28704 20226 28716
rect 20809 28713 20821 28716
rect 20855 28713 20867 28747
rect 20809 28707 20867 28713
rect 21542 28704 21548 28756
rect 21600 28744 21606 28756
rect 21637 28747 21695 28753
rect 21637 28744 21649 28747
rect 21600 28716 21649 28744
rect 21600 28704 21606 28716
rect 21637 28713 21649 28716
rect 21683 28713 21695 28747
rect 21637 28707 21695 28713
rect 23937 28747 23995 28753
rect 23937 28713 23949 28747
rect 23983 28744 23995 28747
rect 24578 28744 24584 28756
rect 23983 28716 24584 28744
rect 23983 28713 23995 28716
rect 23937 28707 23995 28713
rect 24578 28704 24584 28716
rect 24636 28704 24642 28756
rect 25130 28744 25136 28756
rect 25091 28716 25136 28744
rect 25130 28704 25136 28716
rect 25188 28704 25194 28756
rect 16666 28676 16672 28688
rect 16132 28648 16672 28676
rect 16666 28636 16672 28648
rect 16724 28636 16730 28688
rect 16850 28608 16856 28620
rect 16811 28580 16856 28608
rect 16850 28568 16856 28580
rect 16908 28568 16914 28620
rect 19426 28608 19432 28620
rect 19387 28580 19432 28608
rect 19426 28568 19432 28580
rect 19484 28568 19490 28620
rect 22094 28568 22100 28620
rect 22152 28608 22158 28620
rect 25958 28608 25964 28620
rect 22152 28580 25964 28608
rect 22152 28568 22158 28580
rect 25958 28568 25964 28580
rect 26016 28608 26022 28620
rect 26053 28611 26111 28617
rect 26053 28608 26065 28611
rect 26016 28580 26065 28608
rect 26016 28568 26022 28580
rect 26053 28577 26065 28580
rect 26099 28577 26111 28611
rect 26053 28571 26111 28577
rect 15746 28540 15752 28552
rect 15707 28512 15752 28540
rect 15746 28500 15752 28512
rect 15804 28500 15810 28552
rect 16758 28500 16764 28552
rect 16816 28540 16822 28552
rect 17109 28543 17167 28549
rect 17109 28540 17121 28543
rect 16816 28512 17121 28540
rect 16816 28500 16822 28512
rect 17109 28509 17121 28512
rect 17155 28509 17167 28543
rect 17109 28503 17167 28509
rect 19518 28500 19524 28552
rect 19576 28540 19582 28552
rect 19685 28543 19743 28549
rect 19685 28540 19697 28543
rect 19576 28512 19697 28540
rect 19576 28500 19582 28512
rect 19685 28509 19697 28512
rect 19731 28509 19743 28543
rect 19685 28503 19743 28509
rect 20530 28500 20536 28552
rect 20588 28540 20594 28552
rect 21453 28543 21511 28549
rect 21453 28540 21465 28543
rect 20588 28512 21465 28540
rect 20588 28500 20594 28512
rect 21453 28509 21465 28512
rect 21499 28509 21511 28543
rect 23658 28540 23664 28552
rect 23619 28512 23664 28540
rect 21453 28503 21511 28509
rect 23658 28500 23664 28512
rect 23716 28500 23722 28552
rect 23842 28500 23848 28552
rect 23900 28540 23906 28552
rect 23937 28543 23995 28549
rect 23937 28540 23949 28543
rect 23900 28512 23949 28540
rect 23900 28500 23906 28512
rect 23937 28509 23949 28512
rect 23983 28540 23995 28543
rect 24670 28540 24676 28552
rect 23983 28512 24676 28540
rect 23983 28509 23995 28512
rect 23937 28503 23995 28509
rect 24670 28500 24676 28512
rect 24728 28500 24734 28552
rect 24857 28543 24915 28549
rect 24857 28509 24869 28543
rect 24903 28509 24915 28543
rect 24857 28503 24915 28509
rect 15930 28432 15936 28484
rect 15988 28472 15994 28484
rect 16117 28475 16175 28481
rect 16117 28472 16129 28475
rect 15988 28444 16129 28472
rect 15988 28432 15994 28444
rect 16117 28441 16129 28444
rect 16163 28441 16175 28475
rect 16117 28435 16175 28441
rect 23382 28432 23388 28484
rect 23440 28472 23446 28484
rect 23753 28475 23811 28481
rect 23753 28472 23765 28475
rect 23440 28444 23765 28472
rect 23440 28432 23446 28444
rect 23753 28441 23765 28444
rect 23799 28472 23811 28475
rect 24394 28472 24400 28484
rect 23799 28444 24400 28472
rect 23799 28441 23811 28444
rect 23753 28435 23811 28441
rect 24394 28432 24400 28444
rect 24452 28432 24458 28484
rect 24872 28472 24900 28503
rect 24946 28500 24952 28552
rect 25004 28540 25010 28552
rect 25225 28543 25283 28549
rect 25004 28512 25049 28540
rect 25004 28500 25010 28512
rect 25225 28509 25237 28543
rect 25271 28540 25283 28543
rect 25590 28540 25596 28552
rect 25271 28512 25596 28540
rect 25271 28509 25283 28512
rect 25225 28503 25283 28509
rect 25590 28500 25596 28512
rect 25648 28500 25654 28552
rect 25038 28472 25044 28484
rect 24872 28444 25044 28472
rect 25038 28432 25044 28444
rect 25096 28432 25102 28484
rect 26142 28432 26148 28484
rect 26200 28472 26206 28484
rect 26298 28475 26356 28481
rect 26298 28472 26310 28475
rect 26200 28444 26310 28472
rect 26200 28432 26206 28444
rect 26298 28441 26310 28444
rect 26344 28441 26356 28475
rect 26298 28435 26356 28441
rect 18230 28364 18236 28416
rect 18288 28404 18294 28416
rect 19058 28404 19064 28416
rect 18288 28376 19064 28404
rect 18288 28364 18294 28376
rect 19058 28364 19064 28376
rect 19116 28364 19122 28416
rect 24857 28407 24915 28413
rect 24857 28373 24869 28407
rect 24903 28404 24915 28407
rect 25682 28404 25688 28416
rect 24903 28376 25688 28404
rect 24903 28373 24915 28376
rect 24857 28367 24915 28373
rect 25682 28364 25688 28376
rect 25740 28364 25746 28416
rect 26050 28364 26056 28416
rect 26108 28404 26114 28416
rect 27433 28407 27491 28413
rect 27433 28404 27445 28407
rect 26108 28376 27445 28404
rect 26108 28364 26114 28376
rect 27433 28373 27445 28376
rect 27479 28373 27491 28407
rect 27433 28367 27491 28373
rect 1104 28314 29048 28336
rect 1104 28262 7896 28314
rect 7948 28262 7960 28314
rect 8012 28262 8024 28314
rect 8076 28262 8088 28314
rect 8140 28262 8152 28314
rect 8204 28262 14842 28314
rect 14894 28262 14906 28314
rect 14958 28262 14970 28314
rect 15022 28262 15034 28314
rect 15086 28262 15098 28314
rect 15150 28262 21788 28314
rect 21840 28262 21852 28314
rect 21904 28262 21916 28314
rect 21968 28262 21980 28314
rect 22032 28262 22044 28314
rect 22096 28262 28734 28314
rect 28786 28262 28798 28314
rect 28850 28262 28862 28314
rect 28914 28262 28926 28314
rect 28978 28262 28990 28314
rect 29042 28262 29048 28314
rect 1104 28240 29048 28262
rect 19981 28203 20039 28209
rect 19981 28169 19993 28203
rect 20027 28200 20039 28203
rect 20346 28200 20352 28212
rect 20027 28172 20352 28200
rect 20027 28169 20039 28172
rect 19981 28163 20039 28169
rect 20346 28160 20352 28172
rect 20404 28160 20410 28212
rect 24486 28200 24492 28212
rect 24447 28172 24492 28200
rect 24486 28160 24492 28172
rect 24544 28160 24550 28212
rect 26142 28200 26148 28212
rect 26103 28172 26148 28200
rect 26142 28160 26148 28172
rect 26200 28160 26206 28212
rect 18230 28132 18236 28144
rect 18191 28104 18236 28132
rect 18230 28092 18236 28104
rect 18288 28092 18294 28144
rect 21082 28132 21088 28144
rect 18800 28104 21088 28132
rect 1578 28064 1584 28076
rect 1539 28036 1584 28064
rect 1578 28024 1584 28036
rect 1636 28024 1642 28076
rect 18800 28073 18828 28104
rect 21082 28092 21088 28104
rect 21140 28092 21146 28144
rect 25038 28092 25044 28144
rect 25096 28132 25102 28144
rect 26510 28132 26516 28144
rect 25096 28104 26516 28132
rect 25096 28092 25102 28104
rect 18049 28067 18107 28073
rect 18049 28033 18061 28067
rect 18095 28033 18107 28067
rect 18049 28027 18107 28033
rect 18325 28067 18383 28073
rect 18325 28033 18337 28067
rect 18371 28033 18383 28067
rect 18325 28027 18383 28033
rect 18785 28067 18843 28073
rect 18785 28033 18797 28067
rect 18831 28033 18843 28067
rect 18785 28027 18843 28033
rect 18064 27928 18092 28027
rect 18340 27996 18368 28027
rect 18874 28024 18880 28076
rect 18932 28064 18938 28076
rect 19058 28064 19064 28076
rect 18932 28036 18977 28064
rect 19019 28036 19064 28064
rect 18932 28024 18938 28036
rect 19058 28024 19064 28036
rect 19116 28024 19122 28076
rect 19150 28024 19156 28076
rect 19208 28064 19214 28076
rect 19886 28064 19892 28076
rect 19208 28036 19253 28064
rect 19847 28036 19892 28064
rect 19208 28024 19214 28036
rect 19886 28024 19892 28036
rect 19944 28024 19950 28076
rect 23382 28064 23388 28076
rect 23343 28036 23388 28064
rect 23382 28024 23388 28036
rect 23440 28024 23446 28076
rect 23474 28024 23480 28076
rect 23532 28064 23538 28076
rect 23661 28067 23719 28073
rect 23661 28064 23673 28067
rect 23532 28036 23673 28064
rect 23532 28024 23538 28036
rect 23661 28033 23673 28036
rect 23707 28033 23719 28067
rect 23661 28027 23719 28033
rect 24121 28067 24179 28073
rect 24121 28033 24133 28067
rect 24167 28064 24179 28067
rect 24167 28036 24808 28064
rect 24167 28033 24179 28036
rect 24121 28027 24179 28033
rect 19168 27996 19196 28024
rect 18340 27968 19196 27996
rect 23676 27996 23704 28027
rect 24213 27999 24271 28005
rect 24213 27996 24225 27999
rect 23676 27968 24225 27996
rect 24213 27965 24225 27968
rect 24259 27965 24271 27999
rect 24213 27959 24271 27965
rect 18874 27928 18880 27940
rect 18064 27900 18880 27928
rect 18874 27888 18880 27900
rect 18932 27888 18938 27940
rect 23569 27931 23627 27937
rect 23569 27897 23581 27931
rect 23615 27928 23627 27931
rect 23658 27928 23664 27940
rect 23615 27900 23664 27928
rect 23615 27897 23627 27900
rect 23569 27891 23627 27897
rect 23658 27888 23664 27900
rect 23716 27928 23722 27940
rect 24320 27928 24348 28036
rect 24780 27996 24808 28036
rect 25130 28024 25136 28076
rect 25188 28064 25194 28076
rect 25501 28067 25559 28073
rect 25501 28064 25513 28067
rect 25188 28036 25513 28064
rect 25188 28024 25194 28036
rect 25501 28033 25513 28036
rect 25547 28033 25559 28067
rect 25682 28064 25688 28076
rect 25643 28036 25688 28064
rect 25501 28027 25559 28033
rect 25682 28024 25688 28036
rect 25740 28024 25746 28076
rect 25792 28073 25820 28104
rect 26510 28092 26516 28104
rect 26568 28092 26574 28144
rect 25777 28067 25835 28073
rect 25777 28033 25789 28067
rect 25823 28033 25835 28067
rect 25777 28027 25835 28033
rect 25869 28067 25927 28073
rect 25869 28033 25881 28067
rect 25915 28064 25927 28067
rect 26050 28064 26056 28076
rect 25915 28036 26056 28064
rect 25915 28033 25927 28036
rect 25869 28027 25927 28033
rect 26050 28024 26056 28036
rect 26108 28064 26114 28076
rect 27341 28067 27399 28073
rect 27341 28064 27353 28067
rect 26108 28036 27353 28064
rect 26108 28024 26114 28036
rect 27341 28033 27353 28036
rect 27387 28033 27399 28067
rect 27341 28027 27399 28033
rect 27525 28067 27583 28073
rect 27525 28033 27537 28067
rect 27571 28033 27583 28067
rect 27525 28027 27583 28033
rect 24780 27968 25728 27996
rect 23716 27900 24348 27928
rect 23716 27888 23722 27900
rect 25700 27872 25728 27968
rect 26602 27956 26608 28008
rect 26660 27996 26666 28008
rect 27540 27996 27568 28027
rect 26660 27968 27568 27996
rect 26660 27956 26666 27968
rect 26142 27888 26148 27940
rect 26200 27928 26206 27940
rect 26200 27900 27384 27928
rect 26200 27888 26206 27900
rect 1762 27860 1768 27872
rect 1723 27832 1768 27860
rect 1762 27820 1768 27832
rect 1820 27820 1826 27872
rect 17865 27863 17923 27869
rect 17865 27829 17877 27863
rect 17911 27860 17923 27863
rect 18782 27860 18788 27872
rect 17911 27832 18788 27860
rect 17911 27829 17923 27832
rect 17865 27823 17923 27829
rect 18782 27820 18788 27832
rect 18840 27820 18846 27872
rect 19337 27863 19395 27869
rect 19337 27829 19349 27863
rect 19383 27860 19395 27863
rect 20530 27860 20536 27872
rect 19383 27832 20536 27860
rect 19383 27829 19395 27832
rect 19337 27823 19395 27829
rect 20530 27820 20536 27832
rect 20588 27820 20594 27872
rect 23014 27820 23020 27872
rect 23072 27860 23078 27872
rect 23201 27863 23259 27869
rect 23201 27860 23213 27863
rect 23072 27832 23213 27860
rect 23072 27820 23078 27832
rect 23201 27829 23213 27832
rect 23247 27829 23259 27863
rect 23201 27823 23259 27829
rect 24305 27863 24363 27869
rect 24305 27829 24317 27863
rect 24351 27860 24363 27863
rect 24854 27860 24860 27872
rect 24351 27832 24860 27860
rect 24351 27829 24363 27832
rect 24305 27823 24363 27829
rect 24854 27820 24860 27832
rect 24912 27820 24918 27872
rect 25682 27820 25688 27872
rect 25740 27860 25746 27872
rect 27356 27869 27384 27900
rect 27157 27863 27215 27869
rect 27157 27860 27169 27863
rect 25740 27832 27169 27860
rect 25740 27820 25746 27832
rect 27157 27829 27169 27832
rect 27203 27829 27215 27863
rect 27157 27823 27215 27829
rect 27341 27863 27399 27869
rect 27341 27829 27353 27863
rect 27387 27829 27399 27863
rect 28166 27860 28172 27872
rect 28127 27832 28172 27860
rect 27341 27823 27399 27829
rect 28166 27820 28172 27832
rect 28224 27820 28230 27872
rect 1104 27770 28888 27792
rect 1104 27718 4423 27770
rect 4475 27718 4487 27770
rect 4539 27718 4551 27770
rect 4603 27718 4615 27770
rect 4667 27718 4679 27770
rect 4731 27718 11369 27770
rect 11421 27718 11433 27770
rect 11485 27718 11497 27770
rect 11549 27718 11561 27770
rect 11613 27718 11625 27770
rect 11677 27718 18315 27770
rect 18367 27718 18379 27770
rect 18431 27718 18443 27770
rect 18495 27718 18507 27770
rect 18559 27718 18571 27770
rect 18623 27718 25261 27770
rect 25313 27718 25325 27770
rect 25377 27718 25389 27770
rect 25441 27718 25453 27770
rect 25505 27718 25517 27770
rect 25569 27718 28888 27770
rect 1104 27696 28888 27718
rect 24946 27616 24952 27668
rect 25004 27656 25010 27668
rect 25133 27659 25191 27665
rect 25133 27656 25145 27659
rect 25004 27628 25145 27656
rect 25004 27616 25010 27628
rect 25133 27625 25145 27628
rect 25179 27625 25191 27659
rect 25133 27619 25191 27625
rect 18046 27588 18052 27600
rect 18007 27560 18052 27588
rect 18046 27548 18052 27560
rect 18104 27548 18110 27600
rect 21450 27548 21456 27600
rect 21508 27588 21514 27600
rect 22097 27591 22155 27597
rect 22097 27588 22109 27591
rect 21508 27560 22109 27588
rect 21508 27548 21514 27560
rect 22097 27557 22109 27560
rect 22143 27557 22155 27591
rect 22097 27551 22155 27557
rect 15378 27520 15384 27532
rect 15339 27492 15384 27520
rect 15378 27480 15384 27492
rect 15436 27480 15442 27532
rect 16669 27455 16727 27461
rect 16669 27421 16681 27455
rect 16715 27452 16727 27455
rect 16758 27452 16764 27464
rect 16715 27424 16764 27452
rect 16715 27421 16727 27424
rect 16669 27415 16727 27421
rect 16758 27412 16764 27424
rect 16816 27412 16822 27464
rect 18064 27452 18092 27548
rect 19426 27480 19432 27532
rect 19484 27520 19490 27532
rect 19981 27523 20039 27529
rect 19981 27520 19993 27523
rect 19484 27492 19993 27520
rect 19484 27480 19490 27492
rect 19981 27489 19993 27492
rect 20027 27489 20039 27523
rect 27522 27520 27528 27532
rect 27483 27492 27528 27520
rect 19981 27483 20039 27489
rect 27522 27480 27528 27492
rect 27580 27480 27586 27532
rect 28166 27480 28172 27532
rect 28224 27520 28230 27532
rect 28353 27523 28411 27529
rect 28353 27520 28365 27523
rect 28224 27492 28365 27520
rect 28224 27480 28230 27492
rect 28353 27489 28365 27492
rect 28399 27489 28411 27523
rect 28353 27483 28411 27489
rect 16868 27424 18092 27452
rect 1762 27344 1768 27396
rect 1820 27384 1826 27396
rect 15473 27387 15531 27393
rect 15473 27384 15485 27387
rect 1820 27356 15485 27384
rect 1820 27344 1826 27356
rect 15473 27353 15485 27356
rect 15519 27353 15531 27387
rect 15473 27347 15531 27353
rect 15565 27387 15623 27393
rect 15565 27353 15577 27387
rect 15611 27384 15623 27387
rect 16868 27384 16896 27424
rect 18782 27412 18788 27464
rect 18840 27452 18846 27464
rect 21821 27455 21879 27461
rect 21821 27452 21833 27455
rect 18840 27424 21833 27452
rect 18840 27412 18846 27424
rect 21821 27421 21833 27424
rect 21867 27421 21879 27455
rect 21821 27415 21879 27421
rect 22097 27455 22155 27461
rect 22097 27421 22109 27455
rect 22143 27452 22155 27455
rect 23014 27452 23020 27464
rect 22143 27424 23020 27452
rect 22143 27421 22155 27424
rect 22097 27415 22155 27421
rect 23014 27412 23020 27424
rect 23072 27412 23078 27464
rect 23842 27452 23848 27464
rect 23803 27424 23848 27452
rect 23842 27412 23848 27424
rect 23900 27412 23906 27464
rect 24026 27452 24032 27464
rect 23987 27424 24032 27452
rect 24026 27412 24032 27424
rect 24084 27412 24090 27464
rect 24854 27412 24860 27464
rect 24912 27452 24918 27464
rect 25317 27455 25375 27461
rect 25317 27452 25329 27455
rect 24912 27424 25329 27452
rect 24912 27412 24918 27424
rect 25317 27421 25329 27424
rect 25363 27452 25375 27455
rect 25593 27455 25651 27461
rect 25363 27424 25452 27452
rect 25363 27421 25375 27424
rect 25317 27415 25375 27421
rect 15611 27356 16896 27384
rect 16936 27387 16994 27393
rect 15611 27353 15623 27356
rect 15565 27347 15623 27353
rect 16936 27353 16948 27387
rect 16982 27384 16994 27387
rect 17034 27384 17040 27396
rect 16982 27356 17040 27384
rect 16982 27353 16994 27356
rect 16936 27347 16994 27353
rect 17034 27344 17040 27356
rect 17092 27344 17098 27396
rect 20248 27387 20306 27393
rect 20248 27353 20260 27387
rect 20294 27384 20306 27387
rect 20806 27384 20812 27396
rect 20294 27356 20812 27384
rect 20294 27353 20306 27356
rect 20248 27347 20306 27353
rect 20806 27344 20812 27356
rect 20864 27344 20870 27396
rect 21913 27387 21971 27393
rect 21913 27353 21925 27387
rect 21959 27384 21971 27387
rect 22370 27384 22376 27396
rect 21959 27356 22376 27384
rect 21959 27353 21971 27356
rect 21913 27347 21971 27353
rect 22370 27344 22376 27356
rect 22428 27344 22434 27396
rect 15654 27276 15660 27328
rect 15712 27316 15718 27328
rect 15933 27319 15991 27325
rect 15933 27316 15945 27319
rect 15712 27288 15945 27316
rect 15712 27276 15718 27288
rect 15933 27285 15945 27288
rect 15979 27285 15991 27319
rect 21358 27316 21364 27328
rect 21319 27288 21364 27316
rect 15933 27279 15991 27285
rect 21358 27276 21364 27288
rect 21416 27276 21422 27328
rect 23934 27316 23940 27328
rect 23895 27288 23940 27316
rect 23934 27276 23940 27288
rect 23992 27276 23998 27328
rect 25424 27316 25452 27424
rect 25593 27421 25605 27455
rect 25639 27452 25651 27455
rect 25866 27452 25872 27464
rect 25639 27424 25872 27452
rect 25639 27421 25651 27424
rect 25593 27415 25651 27421
rect 25866 27412 25872 27424
rect 25924 27412 25930 27464
rect 25501 27387 25559 27393
rect 25501 27353 25513 27387
rect 25547 27384 25559 27387
rect 25682 27384 25688 27396
rect 25547 27356 25688 27384
rect 25547 27353 25559 27356
rect 25501 27347 25559 27353
rect 25682 27344 25688 27356
rect 25740 27344 25746 27396
rect 27890 27344 27896 27396
rect 27948 27384 27954 27396
rect 28169 27387 28227 27393
rect 28169 27384 28181 27387
rect 27948 27356 28181 27384
rect 27948 27344 27954 27356
rect 28169 27353 28181 27356
rect 28215 27353 28227 27387
rect 28169 27347 28227 27353
rect 25590 27316 25596 27328
rect 25424 27288 25596 27316
rect 25590 27276 25596 27288
rect 25648 27276 25654 27328
rect 1104 27226 29048 27248
rect 1104 27174 7896 27226
rect 7948 27174 7960 27226
rect 8012 27174 8024 27226
rect 8076 27174 8088 27226
rect 8140 27174 8152 27226
rect 8204 27174 14842 27226
rect 14894 27174 14906 27226
rect 14958 27174 14970 27226
rect 15022 27174 15034 27226
rect 15086 27174 15098 27226
rect 15150 27174 21788 27226
rect 21840 27174 21852 27226
rect 21904 27174 21916 27226
rect 21968 27174 21980 27226
rect 22032 27174 22044 27226
rect 22096 27174 28734 27226
rect 28786 27174 28798 27226
rect 28850 27174 28862 27226
rect 28914 27174 28926 27226
rect 28978 27174 28990 27226
rect 29042 27174 29048 27226
rect 1104 27152 29048 27174
rect 17034 27112 17040 27124
rect 16995 27084 17040 27112
rect 17034 27072 17040 27084
rect 17092 27072 17098 27124
rect 20714 27112 20720 27124
rect 18524 27084 20720 27112
rect 15565 27047 15623 27053
rect 15565 27013 15577 27047
rect 15611 27044 15623 27047
rect 15654 27044 15660 27056
rect 15611 27016 15660 27044
rect 15611 27013 15623 27016
rect 15565 27007 15623 27013
rect 15654 27004 15660 27016
rect 15712 27004 15718 27056
rect 15749 27047 15807 27053
rect 15749 27013 15761 27047
rect 15795 27044 15807 27047
rect 16206 27044 16212 27056
rect 15795 27016 16212 27044
rect 15795 27013 15807 27016
rect 15749 27007 15807 27013
rect 16206 27004 16212 27016
rect 16264 27044 16270 27056
rect 18524 27053 18552 27084
rect 20714 27072 20720 27084
rect 20772 27072 20778 27124
rect 22462 27112 22468 27124
rect 22066 27084 22468 27112
rect 18509 27047 18567 27053
rect 18509 27044 18521 27047
rect 16264 27016 18521 27044
rect 16264 27004 16270 27016
rect 18509 27013 18521 27016
rect 18555 27013 18567 27047
rect 18509 27007 18567 27013
rect 18693 27047 18751 27053
rect 18693 27013 18705 27047
rect 18739 27044 18751 27047
rect 22066 27044 22094 27084
rect 22462 27072 22468 27084
rect 22520 27072 22526 27124
rect 25866 27112 25872 27124
rect 25827 27084 25872 27112
rect 25866 27072 25872 27084
rect 25924 27072 25930 27124
rect 27890 27112 27896 27124
rect 27851 27084 27896 27112
rect 27890 27072 27896 27084
rect 27948 27072 27954 27124
rect 22189 27047 22247 27053
rect 22189 27044 22201 27047
rect 18739 27016 22201 27044
rect 18739 27013 18751 27016
rect 18693 27007 18751 27013
rect 22189 27013 22201 27016
rect 22235 27013 22247 27047
rect 22189 27007 22247 27013
rect 22278 27004 22284 27056
rect 22336 27044 22342 27056
rect 22373 27047 22431 27053
rect 22373 27044 22385 27047
rect 22336 27016 22385 27044
rect 22336 27004 22342 27016
rect 22373 27013 22385 27016
rect 22419 27044 22431 27047
rect 22738 27044 22744 27056
rect 22419 27016 22744 27044
rect 22419 27013 22431 27016
rect 22373 27007 22431 27013
rect 22738 27004 22744 27016
rect 22796 27004 22802 27056
rect 15933 26979 15991 26985
rect 15933 26945 15945 26979
rect 15979 26976 15991 26979
rect 16853 26979 16911 26985
rect 16853 26976 16865 26979
rect 15979 26948 16865 26976
rect 15979 26945 15991 26948
rect 15933 26939 15991 26945
rect 16853 26945 16865 26948
rect 16899 26945 16911 26979
rect 18782 26976 18788 26988
rect 18743 26948 18788 26976
rect 16853 26939 16911 26945
rect 18782 26936 18788 26948
rect 18840 26936 18846 26988
rect 20990 26936 20996 26988
rect 21048 26976 21054 26988
rect 21174 26976 21180 26988
rect 21048 26948 21180 26976
rect 21048 26936 21054 26948
rect 21174 26936 21180 26948
rect 21232 26976 21238 26988
rect 21269 26979 21327 26985
rect 21269 26976 21281 26979
rect 21232 26948 21281 26976
rect 21232 26936 21238 26948
rect 21269 26945 21281 26948
rect 21315 26945 21327 26979
rect 21450 26976 21456 26988
rect 21411 26948 21456 26976
rect 21269 26939 21327 26945
rect 21450 26936 21456 26948
rect 21508 26936 21514 26988
rect 26142 26976 26148 26988
rect 26103 26948 26148 26976
rect 26142 26936 26148 26948
rect 26200 26936 26206 26988
rect 27614 26936 27620 26988
rect 27672 26976 27678 26988
rect 27801 26979 27859 26985
rect 27801 26976 27813 26979
rect 27672 26948 27813 26976
rect 27672 26936 27678 26948
rect 27801 26945 27813 26948
rect 27847 26945 27859 26979
rect 27801 26939 27859 26945
rect 25869 26911 25927 26917
rect 25869 26877 25881 26911
rect 25915 26908 25927 26911
rect 26050 26908 26056 26920
rect 25915 26880 26056 26908
rect 25915 26877 25927 26880
rect 25869 26871 25927 26877
rect 26050 26868 26056 26880
rect 26108 26868 26114 26920
rect 21542 26800 21548 26852
rect 21600 26840 21606 26852
rect 22005 26843 22063 26849
rect 22005 26840 22017 26843
rect 21600 26812 22017 26840
rect 21600 26800 21606 26812
rect 22005 26809 22017 26812
rect 22051 26809 22063 26843
rect 26602 26840 26608 26852
rect 22005 26803 22063 26809
rect 26068 26812 26608 26840
rect 17034 26732 17040 26784
rect 17092 26772 17098 26784
rect 18509 26775 18567 26781
rect 18509 26772 18521 26775
rect 17092 26744 18521 26772
rect 17092 26732 17098 26744
rect 18509 26741 18521 26744
rect 18555 26741 18567 26775
rect 18509 26735 18567 26741
rect 21453 26775 21511 26781
rect 21453 26741 21465 26775
rect 21499 26772 21511 26775
rect 21726 26772 21732 26784
rect 21499 26744 21732 26772
rect 21499 26741 21511 26744
rect 21453 26735 21511 26741
rect 21726 26732 21732 26744
rect 21784 26732 21790 26784
rect 26068 26781 26096 26812
rect 26602 26800 26608 26812
rect 26660 26800 26666 26852
rect 26053 26775 26111 26781
rect 26053 26741 26065 26775
rect 26099 26741 26111 26775
rect 26053 26735 26111 26741
rect 26510 26732 26516 26784
rect 26568 26772 26574 26784
rect 27157 26775 27215 26781
rect 27157 26772 27169 26775
rect 26568 26744 27169 26772
rect 26568 26732 26574 26744
rect 27157 26741 27169 26744
rect 27203 26741 27215 26775
rect 27157 26735 27215 26741
rect 1104 26682 28888 26704
rect 1104 26630 4423 26682
rect 4475 26630 4487 26682
rect 4539 26630 4551 26682
rect 4603 26630 4615 26682
rect 4667 26630 4679 26682
rect 4731 26630 11369 26682
rect 11421 26630 11433 26682
rect 11485 26630 11497 26682
rect 11549 26630 11561 26682
rect 11613 26630 11625 26682
rect 11677 26630 18315 26682
rect 18367 26630 18379 26682
rect 18431 26630 18443 26682
rect 18495 26630 18507 26682
rect 18559 26630 18571 26682
rect 18623 26630 25261 26682
rect 25313 26630 25325 26682
rect 25377 26630 25389 26682
rect 25441 26630 25453 26682
rect 25505 26630 25517 26682
rect 25569 26630 28888 26682
rect 1104 26608 28888 26630
rect 19521 26571 19579 26577
rect 19521 26537 19533 26571
rect 19567 26568 19579 26571
rect 20070 26568 20076 26580
rect 19567 26540 20076 26568
rect 19567 26537 19579 26540
rect 19521 26531 19579 26537
rect 20070 26528 20076 26540
rect 20128 26528 20134 26580
rect 22186 26568 22192 26580
rect 21928 26540 22192 26568
rect 16666 26460 16672 26512
rect 16724 26500 16730 26512
rect 17037 26503 17095 26509
rect 17037 26500 17049 26503
rect 16724 26472 17049 26500
rect 16724 26460 16730 26472
rect 17037 26469 17049 26472
rect 17083 26500 17095 26503
rect 17402 26500 17408 26512
rect 17083 26472 17408 26500
rect 17083 26469 17095 26472
rect 17037 26463 17095 26469
rect 17402 26460 17408 26472
rect 17460 26460 17466 26512
rect 20993 26435 21051 26441
rect 20993 26401 21005 26435
rect 21039 26432 21051 26435
rect 21358 26432 21364 26444
rect 21039 26404 21364 26432
rect 21039 26401 21051 26404
rect 20993 26395 21051 26401
rect 21358 26392 21364 26404
rect 21416 26392 21422 26444
rect 21928 26441 21956 26540
rect 22186 26528 22192 26540
rect 22244 26528 22250 26580
rect 23293 26571 23351 26577
rect 23293 26537 23305 26571
rect 23339 26568 23351 26571
rect 23382 26568 23388 26580
rect 23339 26540 23388 26568
rect 23339 26537 23351 26540
rect 23293 26531 23351 26537
rect 23382 26528 23388 26540
rect 23440 26528 23446 26580
rect 21913 26435 21971 26441
rect 21913 26401 21925 26435
rect 21959 26401 21971 26435
rect 26510 26432 26516 26444
rect 26471 26404 26516 26432
rect 21913 26395 21971 26401
rect 26510 26392 26516 26404
rect 26568 26392 26574 26444
rect 28350 26432 28356 26444
rect 28311 26404 28356 26432
rect 28350 26392 28356 26404
rect 28408 26392 28414 26444
rect 1670 26324 1676 26376
rect 1728 26364 1734 26376
rect 1765 26367 1823 26373
rect 1765 26364 1777 26367
rect 1728 26336 1777 26364
rect 1728 26324 1734 26336
rect 1765 26333 1777 26336
rect 1811 26333 1823 26367
rect 1765 26327 1823 26333
rect 16853 26367 16911 26373
rect 16853 26333 16865 26367
rect 16899 26364 16911 26367
rect 17034 26364 17040 26376
rect 16899 26336 17040 26364
rect 16899 26333 16911 26336
rect 16853 26327 16911 26333
rect 17034 26324 17040 26336
rect 17092 26324 17098 26376
rect 19426 26364 19432 26376
rect 19387 26336 19432 26364
rect 19426 26324 19432 26336
rect 19484 26324 19490 26376
rect 21453 26367 21511 26373
rect 21453 26333 21465 26367
rect 21499 26364 21511 26367
rect 21542 26364 21548 26376
rect 21499 26336 21548 26364
rect 21499 26333 21511 26336
rect 21453 26327 21511 26333
rect 21542 26324 21548 26336
rect 21600 26324 21606 26376
rect 21726 26324 21732 26376
rect 21784 26364 21790 26376
rect 22169 26367 22227 26373
rect 22169 26364 22181 26367
rect 21784 26336 22181 26364
rect 21784 26324 21790 26336
rect 22169 26333 22181 26336
rect 22215 26333 22227 26367
rect 22169 26327 22227 26333
rect 24486 26324 24492 26376
rect 24544 26364 24550 26376
rect 24581 26367 24639 26373
rect 24581 26364 24593 26367
rect 24544 26336 24593 26364
rect 24544 26324 24550 26336
rect 24581 26333 24593 26336
rect 24627 26333 24639 26367
rect 24581 26327 24639 26333
rect 21361 26299 21419 26305
rect 21361 26265 21373 26299
rect 21407 26296 21419 26299
rect 21634 26296 21640 26308
rect 21407 26268 21640 26296
rect 21407 26265 21419 26268
rect 21361 26259 21419 26265
rect 21634 26256 21640 26268
rect 21692 26256 21698 26308
rect 26694 26296 26700 26308
rect 26655 26268 26700 26296
rect 26694 26256 26700 26268
rect 26752 26256 26758 26308
rect 21266 26228 21272 26240
rect 21227 26200 21272 26228
rect 21266 26188 21272 26200
rect 21324 26188 21330 26240
rect 24670 26228 24676 26240
rect 24631 26200 24676 26228
rect 24670 26188 24676 26200
rect 24728 26188 24734 26240
rect 1104 26138 29048 26160
rect 1104 26086 7896 26138
rect 7948 26086 7960 26138
rect 8012 26086 8024 26138
rect 8076 26086 8088 26138
rect 8140 26086 8152 26138
rect 8204 26086 14842 26138
rect 14894 26086 14906 26138
rect 14958 26086 14970 26138
rect 15022 26086 15034 26138
rect 15086 26086 15098 26138
rect 15150 26086 21788 26138
rect 21840 26086 21852 26138
rect 21904 26086 21916 26138
rect 21968 26086 21980 26138
rect 22032 26086 22044 26138
rect 22096 26086 28734 26138
rect 28786 26086 28798 26138
rect 28850 26086 28862 26138
rect 28914 26086 28926 26138
rect 28978 26086 28990 26138
rect 29042 26086 29048 26138
rect 1104 26064 29048 26086
rect 15933 26027 15991 26033
rect 15933 25993 15945 26027
rect 15979 26024 15991 26027
rect 18233 26027 18291 26033
rect 18233 26024 18245 26027
rect 15979 25996 18245 26024
rect 15979 25993 15991 25996
rect 15933 25987 15991 25993
rect 18233 25993 18245 25996
rect 18279 26024 18291 26027
rect 19886 26024 19892 26036
rect 18279 25996 19892 26024
rect 18279 25993 18291 25996
rect 18233 25987 18291 25993
rect 19886 25984 19892 25996
rect 19944 25984 19950 26036
rect 21085 26027 21143 26033
rect 21085 25993 21097 26027
rect 21131 26024 21143 26027
rect 21358 26024 21364 26036
rect 21131 25996 21364 26024
rect 21131 25993 21143 25996
rect 21085 25987 21143 25993
rect 21358 25984 21364 25996
rect 21416 25984 21422 26036
rect 23842 25984 23848 26036
rect 23900 26024 23906 26036
rect 24578 26024 24584 26036
rect 23900 25996 24584 26024
rect 23900 25984 23906 25996
rect 24578 25984 24584 25996
rect 24636 26024 24642 26036
rect 24636 25996 24900 26024
rect 24636 25984 24642 25996
rect 23937 25959 23995 25965
rect 16868 25928 18828 25956
rect 1670 25888 1676 25900
rect 1631 25860 1676 25888
rect 1670 25848 1676 25860
rect 1728 25848 1734 25900
rect 16758 25848 16764 25900
rect 16816 25888 16822 25900
rect 16868 25897 16896 25928
rect 17126 25897 17132 25900
rect 16853 25891 16911 25897
rect 16853 25888 16865 25891
rect 16816 25860 16865 25888
rect 16816 25848 16822 25860
rect 16853 25857 16865 25860
rect 16899 25857 16911 25891
rect 16853 25851 16911 25857
rect 17120 25851 17132 25897
rect 17184 25888 17190 25900
rect 18800 25897 18828 25928
rect 23937 25925 23949 25959
rect 23983 25956 23995 25959
rect 24762 25956 24768 25968
rect 23983 25928 24768 25956
rect 23983 25925 23995 25928
rect 23937 25919 23995 25925
rect 24762 25916 24768 25928
rect 24820 25916 24826 25968
rect 18785 25891 18843 25897
rect 17184 25860 17220 25888
rect 17126 25848 17132 25851
rect 17184 25848 17190 25860
rect 18785 25857 18797 25891
rect 18831 25857 18843 25891
rect 18785 25851 18843 25857
rect 18874 25848 18880 25900
rect 18932 25888 18938 25900
rect 19041 25891 19099 25897
rect 19041 25888 19053 25891
rect 18932 25860 19053 25888
rect 18932 25848 18938 25860
rect 19041 25857 19053 25860
rect 19087 25857 19099 25891
rect 19041 25851 19099 25857
rect 20162 25848 20168 25900
rect 20220 25888 20226 25900
rect 20993 25891 21051 25897
rect 20993 25888 21005 25891
rect 20220 25860 21005 25888
rect 20220 25848 20226 25860
rect 20993 25857 21005 25860
rect 21039 25857 21051 25891
rect 24670 25888 24676 25900
rect 24631 25860 24676 25888
rect 20993 25851 21051 25857
rect 24670 25848 24676 25860
rect 24728 25848 24734 25900
rect 24872 25897 24900 25996
rect 26694 25984 26700 26036
rect 26752 26024 26758 26036
rect 27249 26027 27307 26033
rect 27249 26024 27261 26027
rect 26752 25996 27261 26024
rect 26752 25984 26758 25996
rect 27249 25993 27261 25996
rect 27295 25993 27307 26027
rect 27249 25987 27307 25993
rect 26513 25959 26571 25965
rect 26513 25956 26525 25959
rect 25700 25928 26525 25956
rect 25700 25897 25728 25928
rect 26513 25925 26525 25928
rect 26559 25925 26571 25959
rect 26513 25919 26571 25925
rect 24857 25891 24915 25897
rect 24857 25857 24869 25891
rect 24903 25857 24915 25891
rect 25685 25891 25743 25897
rect 25685 25888 25697 25891
rect 24857 25851 24915 25857
rect 24964 25860 25697 25888
rect 1857 25823 1915 25829
rect 1857 25789 1869 25823
rect 1903 25820 1915 25823
rect 2406 25820 2412 25832
rect 1903 25792 2412 25820
rect 1903 25789 1915 25792
rect 1857 25783 1915 25789
rect 2406 25780 2412 25792
rect 2464 25780 2470 25832
rect 2774 25820 2780 25832
rect 2735 25792 2780 25820
rect 2774 25780 2780 25792
rect 2832 25780 2838 25832
rect 15562 25780 15568 25832
rect 15620 25820 15626 25832
rect 15657 25823 15715 25829
rect 15657 25820 15669 25823
rect 15620 25792 15669 25820
rect 15620 25780 15626 25792
rect 15657 25789 15669 25792
rect 15703 25789 15715 25823
rect 15838 25820 15844 25832
rect 15799 25792 15844 25820
rect 15657 25783 15715 25789
rect 15838 25780 15844 25792
rect 15896 25780 15902 25832
rect 19978 25780 19984 25832
rect 20036 25820 20042 25832
rect 20898 25820 20904 25832
rect 20036 25792 20904 25820
rect 20036 25780 20042 25792
rect 20898 25780 20904 25792
rect 20956 25820 20962 25832
rect 21177 25823 21235 25829
rect 21177 25820 21189 25823
rect 20956 25792 21189 25820
rect 20956 25780 20962 25792
rect 21177 25789 21189 25792
rect 21223 25789 21235 25823
rect 21177 25783 21235 25789
rect 23382 25780 23388 25832
rect 23440 25820 23446 25832
rect 24964 25820 24992 25860
rect 25685 25857 25697 25860
rect 25731 25857 25743 25891
rect 25685 25851 25743 25857
rect 25774 25848 25780 25900
rect 25832 25888 25838 25900
rect 26329 25891 26387 25897
rect 26329 25888 26341 25891
rect 25832 25860 26341 25888
rect 25832 25848 25838 25860
rect 26329 25857 26341 25860
rect 26375 25857 26387 25891
rect 26329 25851 26387 25857
rect 26602 25848 26608 25900
rect 26660 25888 26666 25900
rect 26660 25860 26705 25888
rect 26660 25848 26666 25860
rect 26878 25848 26884 25900
rect 26936 25888 26942 25900
rect 27157 25891 27215 25897
rect 27157 25888 27169 25891
rect 26936 25860 27169 25888
rect 26936 25848 26942 25860
rect 27157 25857 27169 25860
rect 27203 25857 27215 25891
rect 27157 25851 27215 25857
rect 23440 25792 24992 25820
rect 23440 25780 23446 25792
rect 25038 25780 25044 25832
rect 25096 25820 25102 25832
rect 25133 25823 25191 25829
rect 25133 25820 25145 25823
rect 25096 25792 25145 25820
rect 25096 25780 25102 25792
rect 25133 25789 25145 25792
rect 25179 25820 25191 25823
rect 26142 25820 26148 25832
rect 25179 25792 26148 25820
rect 25179 25789 25191 25792
rect 25133 25783 25191 25789
rect 26142 25780 26148 25792
rect 26200 25780 26206 25832
rect 26329 25755 26387 25761
rect 26329 25721 26341 25755
rect 26375 25752 26387 25755
rect 27338 25752 27344 25764
rect 26375 25724 27344 25752
rect 26375 25721 26387 25724
rect 26329 25715 26387 25721
rect 27338 25712 27344 25724
rect 27396 25712 27402 25764
rect 16114 25644 16120 25696
rect 16172 25684 16178 25696
rect 16301 25687 16359 25693
rect 16301 25684 16313 25687
rect 16172 25656 16313 25684
rect 16172 25644 16178 25656
rect 16301 25653 16313 25656
rect 16347 25653 16359 25687
rect 20162 25684 20168 25696
rect 20123 25656 20168 25684
rect 16301 25647 16359 25653
rect 20162 25644 20168 25656
rect 20220 25644 20226 25696
rect 20622 25684 20628 25696
rect 20583 25656 20628 25684
rect 20622 25644 20628 25656
rect 20680 25644 20686 25696
rect 22465 25687 22523 25693
rect 22465 25653 22477 25687
rect 22511 25684 22523 25687
rect 22554 25684 22560 25696
rect 22511 25656 22560 25684
rect 22511 25653 22523 25656
rect 22465 25647 22523 25653
rect 22554 25644 22560 25656
rect 22612 25644 22618 25696
rect 24026 25644 24032 25696
rect 24084 25684 24090 25696
rect 24670 25684 24676 25696
rect 24084 25656 24676 25684
rect 24084 25644 24090 25656
rect 24670 25644 24676 25656
rect 24728 25644 24734 25696
rect 25590 25644 25596 25696
rect 25648 25684 25654 25696
rect 25869 25687 25927 25693
rect 25869 25684 25881 25687
rect 25648 25656 25881 25684
rect 25648 25644 25654 25656
rect 25869 25653 25881 25656
rect 25915 25684 25927 25687
rect 26050 25684 26056 25696
rect 25915 25656 26056 25684
rect 25915 25653 25927 25656
rect 25869 25647 25927 25653
rect 26050 25644 26056 25656
rect 26108 25644 26114 25696
rect 27985 25687 28043 25693
rect 27985 25653 27997 25687
rect 28031 25684 28043 25687
rect 28350 25684 28356 25696
rect 28031 25656 28356 25684
rect 28031 25653 28043 25656
rect 27985 25647 28043 25653
rect 28350 25644 28356 25656
rect 28408 25644 28414 25696
rect 1104 25594 28888 25616
rect 1104 25542 4423 25594
rect 4475 25542 4487 25594
rect 4539 25542 4551 25594
rect 4603 25542 4615 25594
rect 4667 25542 4679 25594
rect 4731 25542 11369 25594
rect 11421 25542 11433 25594
rect 11485 25542 11497 25594
rect 11549 25542 11561 25594
rect 11613 25542 11625 25594
rect 11677 25542 18315 25594
rect 18367 25542 18379 25594
rect 18431 25542 18443 25594
rect 18495 25542 18507 25594
rect 18559 25542 18571 25594
rect 18623 25542 25261 25594
rect 25313 25542 25325 25594
rect 25377 25542 25389 25594
rect 25441 25542 25453 25594
rect 25505 25542 25517 25594
rect 25569 25542 28888 25594
rect 1104 25520 28888 25542
rect 2406 25480 2412 25492
rect 2367 25452 2412 25480
rect 2406 25440 2412 25452
rect 2464 25440 2470 25492
rect 17126 25480 17132 25492
rect 17087 25452 17132 25480
rect 17126 25440 17132 25452
rect 17184 25440 17190 25492
rect 18874 25480 18880 25492
rect 18835 25452 18880 25480
rect 18874 25440 18880 25452
rect 18932 25440 18938 25492
rect 20806 25480 20812 25492
rect 20767 25452 20812 25480
rect 20806 25440 20812 25452
rect 20864 25440 20870 25492
rect 23382 25480 23388 25492
rect 23343 25452 23388 25480
rect 23382 25440 23388 25452
rect 23440 25440 23446 25492
rect 24578 25440 24584 25492
rect 24636 25480 24642 25492
rect 24673 25483 24731 25489
rect 24673 25480 24685 25483
rect 24636 25452 24685 25480
rect 24636 25440 24642 25452
rect 24673 25449 24685 25452
rect 24719 25449 24731 25483
rect 24673 25443 24731 25449
rect 25685 25483 25743 25489
rect 25685 25449 25697 25483
rect 25731 25480 25743 25483
rect 25774 25480 25780 25492
rect 25731 25452 25780 25480
rect 25731 25449 25743 25452
rect 25685 25443 25743 25449
rect 25774 25440 25780 25452
rect 25832 25440 25838 25492
rect 20622 25344 20628 25356
rect 19628 25316 20628 25344
rect 1578 25276 1584 25288
rect 1539 25248 1584 25276
rect 1578 25236 1584 25248
rect 1636 25236 1642 25288
rect 2501 25279 2559 25285
rect 2501 25245 2513 25279
rect 2547 25276 2559 25279
rect 4246 25276 4252 25288
rect 2547 25248 4252 25276
rect 2547 25245 2559 25248
rect 2501 25239 2559 25245
rect 4246 25236 4252 25248
rect 4304 25236 4310 25288
rect 16114 25276 16120 25288
rect 16075 25248 16120 25276
rect 16114 25236 16120 25248
rect 16172 25236 16178 25288
rect 19628 25285 19656 25316
rect 20622 25304 20628 25316
rect 20680 25304 20686 25356
rect 21266 25344 21272 25356
rect 21227 25316 21272 25344
rect 21266 25304 21272 25316
rect 21324 25304 21330 25356
rect 22462 25304 22468 25356
rect 22520 25344 22526 25356
rect 23293 25347 23351 25353
rect 23293 25344 23305 25347
rect 22520 25316 23305 25344
rect 22520 25304 22526 25316
rect 23293 25313 23305 25316
rect 23339 25313 23351 25347
rect 24762 25344 24768 25356
rect 24723 25316 24768 25344
rect 23293 25307 23351 25313
rect 24762 25304 24768 25316
rect 24820 25304 24826 25356
rect 24946 25304 24952 25356
rect 25004 25344 25010 25356
rect 25958 25344 25964 25356
rect 25004 25316 25964 25344
rect 25004 25304 25010 25316
rect 16485 25279 16543 25285
rect 16485 25245 16497 25279
rect 16531 25276 16543 25279
rect 16945 25279 17003 25285
rect 16945 25276 16957 25279
rect 16531 25248 16957 25276
rect 16531 25245 16543 25248
rect 16485 25239 16543 25245
rect 16945 25245 16957 25248
rect 16991 25245 17003 25279
rect 16945 25239 17003 25245
rect 18693 25279 18751 25285
rect 18693 25245 18705 25279
rect 18739 25276 18751 25279
rect 19429 25279 19487 25285
rect 19429 25276 19441 25279
rect 18739 25248 19441 25276
rect 18739 25245 18751 25248
rect 18693 25239 18751 25245
rect 19429 25245 19441 25248
rect 19475 25245 19487 25279
rect 19429 25239 19487 25245
rect 19613 25279 19671 25285
rect 19613 25245 19625 25279
rect 19659 25245 19671 25279
rect 19613 25239 19671 25245
rect 19702 25236 19708 25288
rect 19760 25276 19766 25288
rect 20990 25276 20996 25288
rect 19760 25248 19805 25276
rect 20951 25248 20996 25276
rect 19760 25236 19766 25248
rect 20990 25236 20996 25248
rect 21048 25236 21054 25288
rect 21177 25279 21235 25285
rect 21177 25245 21189 25279
rect 21223 25276 21235 25279
rect 22370 25276 22376 25288
rect 21223 25248 22376 25276
rect 21223 25245 21235 25248
rect 21177 25239 21235 25245
rect 22370 25236 22376 25248
rect 22428 25236 22434 25288
rect 23569 25279 23627 25285
rect 23569 25245 23581 25279
rect 23615 25276 23627 25279
rect 24486 25276 24492 25288
rect 23615 25248 24492 25276
rect 23615 25245 23627 25248
rect 23569 25239 23627 25245
rect 24486 25236 24492 25248
rect 24544 25236 24550 25288
rect 24673 25279 24731 25285
rect 24673 25245 24685 25279
rect 24719 25245 24731 25279
rect 24673 25239 24731 25245
rect 16301 25211 16359 25217
rect 16301 25177 16313 25211
rect 16347 25208 16359 25211
rect 17126 25208 17132 25220
rect 16347 25180 17132 25208
rect 16347 25177 16359 25180
rect 16301 25171 16359 25177
rect 17126 25168 17132 25180
rect 17184 25168 17190 25220
rect 24688 25208 24716 25239
rect 24854 25236 24860 25288
rect 24912 25276 24918 25288
rect 25700 25285 25728 25316
rect 25958 25304 25964 25316
rect 26016 25304 26022 25356
rect 27522 25344 27528 25356
rect 27483 25316 27528 25344
rect 27522 25304 27528 25316
rect 27580 25304 27586 25356
rect 28350 25344 28356 25356
rect 28311 25316 28356 25344
rect 28350 25304 28356 25316
rect 28408 25304 28414 25356
rect 25501 25279 25559 25285
rect 25501 25276 25513 25279
rect 24912 25248 25513 25276
rect 24912 25236 24918 25248
rect 25501 25245 25513 25248
rect 25547 25245 25559 25279
rect 25501 25239 25559 25245
rect 25685 25279 25743 25285
rect 25685 25245 25697 25279
rect 25731 25245 25743 25279
rect 25685 25239 25743 25245
rect 25222 25208 25228 25220
rect 24688 25180 25228 25208
rect 25222 25168 25228 25180
rect 25280 25168 25286 25220
rect 28166 25208 28172 25220
rect 28127 25180 28172 25208
rect 28166 25168 28172 25180
rect 28224 25168 28230 25220
rect 1762 25140 1768 25152
rect 1723 25112 1768 25140
rect 1762 25100 1768 25112
rect 1820 25100 1826 25152
rect 23753 25143 23811 25149
rect 23753 25109 23765 25143
rect 23799 25140 23811 25143
rect 23842 25140 23848 25152
rect 23799 25112 23848 25140
rect 23799 25109 23811 25112
rect 23753 25103 23811 25109
rect 23842 25100 23848 25112
rect 23900 25100 23906 25152
rect 25038 25140 25044 25152
rect 24999 25112 25044 25140
rect 25038 25100 25044 25112
rect 25096 25100 25102 25152
rect 1104 25050 29048 25072
rect 1104 24998 7896 25050
rect 7948 24998 7960 25050
rect 8012 24998 8024 25050
rect 8076 24998 8088 25050
rect 8140 24998 8152 25050
rect 8204 24998 14842 25050
rect 14894 24998 14906 25050
rect 14958 24998 14970 25050
rect 15022 24998 15034 25050
rect 15086 24998 15098 25050
rect 15150 24998 21788 25050
rect 21840 24998 21852 25050
rect 21904 24998 21916 25050
rect 21968 24998 21980 25050
rect 22032 24998 22044 25050
rect 22096 24998 28734 25050
rect 28786 24998 28798 25050
rect 28850 24998 28862 25050
rect 28914 24998 28926 25050
rect 28978 24998 28990 25050
rect 29042 24998 29048 25050
rect 1104 24976 29048 24998
rect 1762 24896 1768 24948
rect 1820 24936 1826 24948
rect 15838 24936 15844 24948
rect 1820 24908 15844 24936
rect 1820 24896 1826 24908
rect 15838 24896 15844 24908
rect 15896 24896 15902 24948
rect 22370 24936 22376 24948
rect 22331 24908 22376 24936
rect 22370 24896 22376 24908
rect 22428 24896 22434 24948
rect 28166 24936 28172 24948
rect 28127 24908 28172 24936
rect 28166 24896 28172 24908
rect 28224 24896 28230 24948
rect 17126 24828 17132 24880
rect 17184 24868 17190 24880
rect 20898 24868 20904 24880
rect 17184 24840 20904 24868
rect 17184 24828 17190 24840
rect 20898 24828 20904 24840
rect 20956 24828 20962 24880
rect 22738 24868 22744 24880
rect 22511 24837 22569 24843
rect 22699 24840 22744 24868
rect 22511 24834 22523 24837
rect 17037 24803 17095 24809
rect 17037 24769 17049 24803
rect 17083 24800 17095 24803
rect 17218 24800 17224 24812
rect 17083 24772 17224 24800
rect 17083 24769 17095 24772
rect 17037 24763 17095 24769
rect 17218 24760 17224 24772
rect 17276 24760 17282 24812
rect 21634 24760 21640 24812
rect 21692 24800 21698 24812
rect 21818 24800 21824 24812
rect 21692 24772 21824 24800
rect 21692 24760 21698 24772
rect 21818 24760 21824 24772
rect 21876 24800 21882 24812
rect 22388 24806 22523 24834
rect 22388 24800 22416 24806
rect 21876 24772 22416 24800
rect 22511 24803 22523 24806
rect 22557 24803 22569 24837
rect 22738 24828 22744 24840
rect 22796 24828 22802 24880
rect 23382 24828 23388 24880
rect 23440 24868 23446 24880
rect 25593 24871 25651 24877
rect 25593 24868 25605 24871
rect 23440 24840 23520 24868
rect 23440 24828 23446 24840
rect 23492 24809 23520 24840
rect 24504 24840 25605 24868
rect 22511 24797 22569 24803
rect 23477 24803 23535 24809
rect 21876 24760 21882 24772
rect 23477 24769 23489 24803
rect 23523 24769 23535 24803
rect 23477 24763 23535 24769
rect 23492 24732 23520 24763
rect 23750 24760 23756 24812
rect 23808 24800 23814 24812
rect 24213 24803 24271 24809
rect 23808 24772 23853 24800
rect 23808 24760 23814 24772
rect 24213 24769 24225 24803
rect 24259 24769 24271 24803
rect 24394 24800 24400 24812
rect 24355 24772 24400 24800
rect 24213 24763 24271 24769
rect 24228 24732 24256 24763
rect 24394 24760 24400 24772
rect 24452 24760 24458 24812
rect 24504 24732 24532 24840
rect 25593 24837 25605 24840
rect 25639 24837 25651 24871
rect 25593 24831 25651 24837
rect 25222 24800 25228 24812
rect 25183 24772 25228 24800
rect 25222 24760 25228 24772
rect 25280 24760 25286 24812
rect 25409 24803 25467 24809
rect 25409 24800 25421 24803
rect 25332 24772 25421 24800
rect 23492 24704 24532 24732
rect 23566 24664 23572 24676
rect 22572 24636 23572 24664
rect 16850 24596 16856 24608
rect 16811 24568 16856 24596
rect 16850 24556 16856 24568
rect 16908 24556 16914 24608
rect 22572 24605 22600 24636
rect 23566 24624 23572 24636
rect 23624 24624 23630 24676
rect 24578 24664 24584 24676
rect 23676 24636 24584 24664
rect 22557 24599 22615 24605
rect 22557 24565 22569 24599
rect 22603 24565 22615 24599
rect 22557 24559 22615 24565
rect 23201 24599 23259 24605
rect 23201 24565 23213 24599
rect 23247 24596 23259 24599
rect 23290 24596 23296 24608
rect 23247 24568 23296 24596
rect 23247 24565 23259 24568
rect 23201 24559 23259 24565
rect 23290 24556 23296 24568
rect 23348 24556 23354 24608
rect 23676 24605 23704 24636
rect 24578 24624 24584 24636
rect 24636 24624 24642 24676
rect 25332 24664 25360 24772
rect 25409 24769 25421 24772
rect 25455 24769 25467 24803
rect 25409 24763 25467 24769
rect 25498 24760 25504 24812
rect 25556 24800 25562 24812
rect 25774 24809 25780 24812
rect 25731 24803 25780 24809
rect 25556 24772 25601 24800
rect 25556 24760 25562 24772
rect 25731 24769 25743 24803
rect 25777 24769 25780 24803
rect 25731 24763 25780 24769
rect 25774 24760 25780 24763
rect 25832 24760 25838 24812
rect 25866 24760 25872 24812
rect 25924 24800 25930 24812
rect 26605 24803 26663 24809
rect 25924 24772 25969 24800
rect 25924 24760 25930 24772
rect 26605 24769 26617 24803
rect 26651 24800 26663 24803
rect 27430 24800 27436 24812
rect 26651 24772 26740 24800
rect 27391 24772 27436 24800
rect 26651 24769 26663 24772
rect 26605 24763 26663 24769
rect 26712 24744 26740 24772
rect 27430 24760 27436 24772
rect 27488 24760 27494 24812
rect 28074 24800 28080 24812
rect 28035 24772 28080 24800
rect 28074 24760 28080 24772
rect 28132 24760 28138 24812
rect 26329 24735 26387 24741
rect 26329 24701 26341 24735
rect 26375 24732 26387 24735
rect 26418 24732 26424 24744
rect 26375 24704 26424 24732
rect 26375 24701 26387 24704
rect 26329 24695 26387 24701
rect 26418 24692 26424 24704
rect 26476 24692 26482 24744
rect 26694 24732 26700 24744
rect 26607 24704 26700 24732
rect 26694 24692 26700 24704
rect 26752 24724 26758 24744
rect 27157 24735 27215 24741
rect 27157 24732 27169 24735
rect 26988 24724 27169 24732
rect 26752 24704 27169 24724
rect 26752 24696 27016 24704
rect 27157 24701 27169 24704
rect 27203 24701 27215 24735
rect 26752 24692 26758 24696
rect 27157 24695 27215 24701
rect 26234 24664 26240 24676
rect 25332 24636 26240 24664
rect 26234 24624 26240 24636
rect 26292 24624 26298 24676
rect 26602 24624 26608 24676
rect 26660 24664 26666 24676
rect 27617 24667 27675 24673
rect 27617 24664 27629 24667
rect 26660 24636 27629 24664
rect 26660 24624 26666 24636
rect 27617 24633 27629 24636
rect 27663 24633 27675 24667
rect 27617 24627 27675 24633
rect 23661 24599 23719 24605
rect 23661 24565 23673 24599
rect 23707 24565 23719 24599
rect 23661 24559 23719 24565
rect 24489 24599 24547 24605
rect 24489 24565 24501 24599
rect 24535 24596 24547 24599
rect 24670 24596 24676 24608
rect 24535 24568 24676 24596
rect 24535 24565 24547 24568
rect 24489 24559 24547 24565
rect 24670 24556 24676 24568
rect 24728 24556 24734 24608
rect 25682 24556 25688 24608
rect 25740 24596 25746 24608
rect 26421 24599 26479 24605
rect 26421 24596 26433 24599
rect 25740 24568 26433 24596
rect 25740 24556 25746 24568
rect 26421 24565 26433 24568
rect 26467 24565 26479 24599
rect 26421 24559 26479 24565
rect 26510 24556 26516 24608
rect 26568 24596 26574 24608
rect 27249 24599 27307 24605
rect 27249 24596 27261 24599
rect 26568 24568 27261 24596
rect 26568 24556 26574 24568
rect 27249 24565 27261 24568
rect 27295 24565 27307 24599
rect 27249 24559 27307 24565
rect 1104 24506 28888 24528
rect 1104 24454 4423 24506
rect 4475 24454 4487 24506
rect 4539 24454 4551 24506
rect 4603 24454 4615 24506
rect 4667 24454 4679 24506
rect 4731 24454 11369 24506
rect 11421 24454 11433 24506
rect 11485 24454 11497 24506
rect 11549 24454 11561 24506
rect 11613 24454 11625 24506
rect 11677 24454 18315 24506
rect 18367 24454 18379 24506
rect 18431 24454 18443 24506
rect 18495 24454 18507 24506
rect 18559 24454 18571 24506
rect 18623 24454 25261 24506
rect 25313 24454 25325 24506
rect 25377 24454 25389 24506
rect 25441 24454 25453 24506
rect 25505 24454 25517 24506
rect 25569 24454 28888 24506
rect 1104 24432 28888 24454
rect 18141 24395 18199 24401
rect 18141 24392 18153 24395
rect 15948 24364 18153 24392
rect 15562 24216 15568 24268
rect 15620 24256 15626 24268
rect 15657 24259 15715 24265
rect 15657 24256 15669 24259
rect 15620 24228 15669 24256
rect 15620 24216 15626 24228
rect 15657 24225 15669 24228
rect 15703 24225 15715 24259
rect 15657 24219 15715 24225
rect 15948 24197 15976 24364
rect 18141 24361 18153 24364
rect 18187 24392 18199 24395
rect 19426 24392 19432 24404
rect 18187 24364 19432 24392
rect 18187 24361 18199 24364
rect 18141 24355 18199 24361
rect 19426 24352 19432 24364
rect 19484 24352 19490 24404
rect 22738 24352 22744 24404
rect 22796 24392 22802 24404
rect 24394 24392 24400 24404
rect 22796 24364 24400 24392
rect 22796 24352 22802 24364
rect 24394 24352 24400 24364
rect 24452 24352 24458 24404
rect 26418 24352 26424 24404
rect 26476 24392 26482 24404
rect 27430 24392 27436 24404
rect 26476 24364 27436 24392
rect 26476 24352 26482 24364
rect 27430 24352 27436 24364
rect 27488 24352 27494 24404
rect 26513 24259 26571 24265
rect 26513 24225 26525 24259
rect 26559 24256 26571 24259
rect 27890 24256 27896 24268
rect 26559 24228 27896 24256
rect 26559 24225 26571 24228
rect 26513 24219 26571 24225
rect 27890 24216 27896 24228
rect 27948 24216 27954 24268
rect 28350 24256 28356 24268
rect 28311 24228 28356 24256
rect 28350 24216 28356 24228
rect 28408 24216 28414 24268
rect 15933 24191 15991 24197
rect 15933 24157 15945 24191
rect 15979 24157 15991 24191
rect 16758 24188 16764 24200
rect 16719 24160 16764 24188
rect 15933 24151 15991 24157
rect 16758 24148 16764 24160
rect 16816 24148 16822 24200
rect 16850 24148 16856 24200
rect 16908 24188 16914 24200
rect 17017 24191 17075 24197
rect 17017 24188 17029 24191
rect 16908 24160 17029 24188
rect 16908 24148 16914 24160
rect 17017 24157 17029 24160
rect 17063 24157 17075 24191
rect 18782 24188 18788 24200
rect 18743 24160 18788 24188
rect 17017 24151 17075 24157
rect 18782 24148 18788 24160
rect 18840 24148 18846 24200
rect 20070 24148 20076 24200
rect 20128 24188 20134 24200
rect 21177 24191 21235 24197
rect 21177 24188 21189 24191
rect 20128 24160 21189 24188
rect 20128 24148 20134 24160
rect 21177 24157 21189 24160
rect 21223 24157 21235 24191
rect 21177 24151 21235 24157
rect 21542 24148 21548 24200
rect 21600 24188 21606 24200
rect 21637 24191 21695 24197
rect 21637 24188 21649 24191
rect 21600 24160 21649 24188
rect 21600 24148 21606 24160
rect 21637 24157 21649 24160
rect 21683 24157 21695 24191
rect 21637 24151 21695 24157
rect 21726 24148 21732 24200
rect 21784 24188 21790 24200
rect 22557 24191 22615 24197
rect 22557 24188 22569 24191
rect 21784 24160 22569 24188
rect 21784 24148 21790 24160
rect 22557 24157 22569 24160
rect 22603 24157 22615 24191
rect 22557 24151 22615 24157
rect 21358 24080 21364 24132
rect 21416 24120 21422 24132
rect 22830 24129 22836 24132
rect 21416 24092 21588 24120
rect 21416 24080 21422 24092
rect 9398 24012 9404 24064
rect 9456 24052 9462 24064
rect 15841 24055 15899 24061
rect 15841 24052 15853 24055
rect 9456 24024 15853 24052
rect 9456 24012 9462 24024
rect 15841 24021 15853 24024
rect 15887 24021 15899 24055
rect 15841 24015 15899 24021
rect 16301 24055 16359 24061
rect 16301 24021 16313 24055
rect 16347 24052 16359 24055
rect 16850 24052 16856 24064
rect 16347 24024 16856 24052
rect 16347 24021 16359 24024
rect 16301 24015 16359 24021
rect 16850 24012 16856 24024
rect 16908 24012 16914 24064
rect 18598 24052 18604 24064
rect 18559 24024 18604 24052
rect 18598 24012 18604 24024
rect 18656 24012 18662 24064
rect 21450 24052 21456 24064
rect 21411 24024 21456 24052
rect 21450 24012 21456 24024
rect 21508 24012 21514 24064
rect 21560 24061 21588 24092
rect 22824 24083 22836 24129
rect 22888 24120 22894 24132
rect 26697 24123 26755 24129
rect 22888 24092 22924 24120
rect 22830 24080 22836 24083
rect 22888 24080 22894 24092
rect 26697 24089 26709 24123
rect 26743 24120 26755 24123
rect 27338 24120 27344 24132
rect 26743 24092 27344 24120
rect 26743 24089 26755 24092
rect 26697 24083 26755 24089
rect 27338 24080 27344 24092
rect 27396 24080 27402 24132
rect 21545 24055 21603 24061
rect 21545 24021 21557 24055
rect 21591 24052 21603 24055
rect 21818 24052 21824 24064
rect 21591 24024 21824 24052
rect 21591 24021 21603 24024
rect 21545 24015 21603 24021
rect 21818 24012 21824 24024
rect 21876 24012 21882 24064
rect 23750 24012 23756 24064
rect 23808 24052 23814 24064
rect 23937 24055 23995 24061
rect 23937 24052 23949 24055
rect 23808 24024 23949 24052
rect 23808 24012 23814 24024
rect 23937 24021 23949 24024
rect 23983 24052 23995 24055
rect 24210 24052 24216 24064
rect 23983 24024 24216 24052
rect 23983 24021 23995 24024
rect 23937 24015 23995 24021
rect 24210 24012 24216 24024
rect 24268 24012 24274 24064
rect 1104 23962 29048 23984
rect 1104 23910 7896 23962
rect 7948 23910 7960 23962
rect 8012 23910 8024 23962
rect 8076 23910 8088 23962
rect 8140 23910 8152 23962
rect 8204 23910 14842 23962
rect 14894 23910 14906 23962
rect 14958 23910 14970 23962
rect 15022 23910 15034 23962
rect 15086 23910 15098 23962
rect 15150 23910 21788 23962
rect 21840 23910 21852 23962
rect 21904 23910 21916 23962
rect 21968 23910 21980 23962
rect 22032 23910 22044 23962
rect 22096 23910 28734 23962
rect 28786 23910 28798 23962
rect 28850 23910 28862 23962
rect 28914 23910 28926 23962
rect 28978 23910 28990 23962
rect 29042 23910 29048 23962
rect 1104 23888 29048 23910
rect 17218 23848 17224 23860
rect 17179 23820 17224 23848
rect 17218 23808 17224 23820
rect 17276 23808 17282 23860
rect 20070 23848 20076 23860
rect 20031 23820 20076 23848
rect 20070 23808 20076 23820
rect 20128 23808 20134 23860
rect 22830 23848 22836 23860
rect 22791 23820 22836 23848
rect 22830 23808 22836 23820
rect 22888 23808 22894 23860
rect 24946 23848 24952 23860
rect 24907 23820 24952 23848
rect 24946 23808 24952 23820
rect 25004 23808 25010 23860
rect 25774 23848 25780 23860
rect 25735 23820 25780 23848
rect 25774 23808 25780 23820
rect 25832 23808 25838 23860
rect 26234 23848 26240 23860
rect 26195 23820 26240 23848
rect 26234 23808 26240 23820
rect 26292 23808 26298 23860
rect 16850 23780 16856 23792
rect 16811 23752 16856 23780
rect 16850 23740 16856 23752
rect 16908 23740 16914 23792
rect 17037 23783 17095 23789
rect 17037 23749 17049 23783
rect 17083 23780 17095 23783
rect 17126 23780 17132 23792
rect 17083 23752 17132 23780
rect 17083 23749 17095 23752
rect 17037 23743 17095 23749
rect 17126 23740 17132 23752
rect 17184 23740 17190 23792
rect 18500 23783 18558 23789
rect 18500 23749 18512 23783
rect 18546 23780 18558 23783
rect 18598 23780 18604 23792
rect 18546 23752 18604 23780
rect 18546 23749 18558 23752
rect 18500 23743 18558 23749
rect 18598 23740 18604 23752
rect 18656 23740 18662 23792
rect 21358 23740 21364 23792
rect 21416 23780 21422 23792
rect 22157 23783 22215 23789
rect 22157 23780 22169 23783
rect 21416 23752 22169 23780
rect 21416 23740 21422 23752
rect 22157 23749 22169 23752
rect 22203 23749 22215 23783
rect 22370 23780 22376 23792
rect 22283 23752 22376 23780
rect 22157 23743 22215 23749
rect 22370 23740 22376 23752
rect 22428 23780 22434 23792
rect 22738 23780 22744 23792
rect 22428 23752 22744 23780
rect 22428 23740 22434 23752
rect 22738 23740 22744 23752
rect 22796 23740 22802 23792
rect 24210 23780 24216 23792
rect 23124 23752 24216 23780
rect 21174 23712 21180 23724
rect 21232 23721 21238 23724
rect 23124 23721 23152 23752
rect 24210 23740 24216 23752
rect 24268 23740 24274 23792
rect 25130 23780 25136 23792
rect 24596 23752 25136 23780
rect 21144 23684 21180 23712
rect 21174 23672 21180 23684
rect 21232 23675 21244 23721
rect 23109 23715 23167 23721
rect 23109 23681 23121 23715
rect 23155 23681 23167 23715
rect 23109 23675 23167 23681
rect 23201 23715 23259 23721
rect 23201 23681 23213 23715
rect 23247 23681 23259 23715
rect 23201 23675 23259 23681
rect 21232 23672 21238 23675
rect 16758 23604 16764 23656
rect 16816 23644 16822 23656
rect 18233 23647 18291 23653
rect 18233 23644 18245 23647
rect 16816 23616 18245 23644
rect 16816 23604 16822 23616
rect 18233 23613 18245 23616
rect 18279 23613 18291 23647
rect 18233 23607 18291 23613
rect 21453 23647 21511 23653
rect 21453 23613 21465 23647
rect 21499 23644 21511 23647
rect 21634 23644 21640 23656
rect 21499 23616 21640 23644
rect 21499 23613 21511 23616
rect 21453 23607 21511 23613
rect 21634 23604 21640 23616
rect 21692 23604 21698 23656
rect 23216 23644 23244 23675
rect 23290 23672 23296 23724
rect 23348 23712 23354 23724
rect 23477 23715 23535 23721
rect 23348 23684 23393 23712
rect 23348 23672 23354 23684
rect 23477 23681 23489 23715
rect 23523 23712 23535 23715
rect 24596 23712 24624 23752
rect 25130 23740 25136 23752
rect 25188 23740 25194 23792
rect 23523 23684 24624 23712
rect 23523 23681 23535 23684
rect 23477 23675 23535 23681
rect 24762 23672 24768 23724
rect 24820 23712 24826 23724
rect 25409 23715 25467 23721
rect 25409 23712 25421 23715
rect 24820 23684 25421 23712
rect 24820 23672 24826 23684
rect 25409 23681 25421 23684
rect 25455 23681 25467 23715
rect 25409 23675 25467 23681
rect 25593 23715 25651 23721
rect 25593 23681 25605 23715
rect 25639 23712 25651 23715
rect 26418 23712 26424 23724
rect 25639 23684 26424 23712
rect 25639 23681 25651 23684
rect 25593 23675 25651 23681
rect 23934 23644 23940 23656
rect 23216 23616 23940 23644
rect 23934 23604 23940 23616
rect 23992 23604 23998 23656
rect 24302 23604 24308 23656
rect 24360 23644 24366 23656
rect 24581 23647 24639 23653
rect 24581 23644 24593 23647
rect 24360 23616 24593 23644
rect 24360 23604 24366 23616
rect 24581 23613 24593 23616
rect 24627 23644 24639 23647
rect 25608 23644 25636 23675
rect 26418 23672 26424 23684
rect 26476 23672 26482 23724
rect 26510 23672 26516 23724
rect 26568 23712 26574 23724
rect 26605 23715 26663 23721
rect 26605 23712 26617 23715
rect 26568 23684 26617 23712
rect 26568 23672 26574 23684
rect 26605 23681 26617 23684
rect 26651 23681 26663 23715
rect 26605 23675 26663 23681
rect 26786 23672 26792 23724
rect 26844 23712 26850 23724
rect 27062 23712 27068 23724
rect 26844 23684 27068 23712
rect 26844 23672 26850 23684
rect 27062 23672 27068 23684
rect 27120 23712 27126 23724
rect 27249 23715 27307 23721
rect 27249 23712 27261 23715
rect 27120 23684 27261 23712
rect 27120 23672 27126 23684
rect 27249 23681 27261 23684
rect 27295 23681 27307 23715
rect 27249 23675 27307 23681
rect 24627 23616 25636 23644
rect 24627 23613 24639 23616
rect 24581 23607 24639 23613
rect 23658 23536 23664 23588
rect 23716 23576 23722 23588
rect 26528 23576 26556 23672
rect 26694 23604 26700 23656
rect 26752 23604 26758 23656
rect 26712 23576 26740 23604
rect 23716 23548 26556 23576
rect 26620 23548 26740 23576
rect 23716 23536 23722 23548
rect 19610 23508 19616 23520
rect 19571 23480 19616 23508
rect 19610 23468 19616 23480
rect 19668 23468 19674 23520
rect 22002 23508 22008 23520
rect 21963 23480 22008 23508
rect 22002 23468 22008 23480
rect 22060 23468 22066 23520
rect 22189 23511 22247 23517
rect 22189 23477 22201 23511
rect 22235 23508 22247 23511
rect 24394 23508 24400 23520
rect 22235 23480 24400 23508
rect 22235 23477 22247 23480
rect 22189 23471 22247 23477
rect 24394 23468 24400 23480
rect 24452 23508 24458 23520
rect 26620 23517 26648 23548
rect 26605 23511 26663 23517
rect 26605 23508 26617 23511
rect 24452 23480 26617 23508
rect 24452 23468 24458 23480
rect 26605 23477 26617 23480
rect 26651 23477 26663 23511
rect 26605 23471 26663 23477
rect 26694 23468 26700 23520
rect 26752 23508 26758 23520
rect 27341 23511 27399 23517
rect 27341 23508 27353 23511
rect 26752 23480 27353 23508
rect 26752 23468 26758 23480
rect 27341 23477 27353 23480
rect 27387 23477 27399 23511
rect 27341 23471 27399 23477
rect 27430 23468 27436 23520
rect 27488 23508 27494 23520
rect 27893 23511 27951 23517
rect 27893 23508 27905 23511
rect 27488 23480 27905 23508
rect 27488 23468 27494 23480
rect 27893 23477 27905 23480
rect 27939 23477 27951 23511
rect 27893 23471 27951 23477
rect 1104 23418 28888 23440
rect 1104 23366 4423 23418
rect 4475 23366 4487 23418
rect 4539 23366 4551 23418
rect 4603 23366 4615 23418
rect 4667 23366 4679 23418
rect 4731 23366 11369 23418
rect 11421 23366 11433 23418
rect 11485 23366 11497 23418
rect 11549 23366 11561 23418
rect 11613 23366 11625 23418
rect 11677 23366 18315 23418
rect 18367 23366 18379 23418
rect 18431 23366 18443 23418
rect 18495 23366 18507 23418
rect 18559 23366 18571 23418
rect 18623 23366 25261 23418
rect 25313 23366 25325 23418
rect 25377 23366 25389 23418
rect 25441 23366 25453 23418
rect 25505 23366 25517 23418
rect 25569 23366 28888 23418
rect 1104 23344 28888 23366
rect 18782 23304 18788 23316
rect 18743 23276 18788 23304
rect 18782 23264 18788 23276
rect 18840 23264 18846 23316
rect 20993 23307 21051 23313
rect 20993 23273 21005 23307
rect 21039 23304 21051 23307
rect 21174 23304 21180 23316
rect 21039 23276 21180 23304
rect 21039 23273 21051 23276
rect 20993 23267 21051 23273
rect 21174 23264 21180 23276
rect 21232 23264 21238 23316
rect 21361 23307 21419 23313
rect 21361 23273 21373 23307
rect 21407 23304 21419 23307
rect 22002 23304 22008 23316
rect 21407 23276 22008 23304
rect 21407 23273 21419 23276
rect 21361 23267 21419 23273
rect 22002 23264 22008 23276
rect 22060 23264 22066 23316
rect 19429 23239 19487 23245
rect 19429 23205 19441 23239
rect 19475 23205 19487 23239
rect 19429 23199 19487 23205
rect 16390 23100 16396 23112
rect 16351 23072 16396 23100
rect 16390 23060 16396 23072
rect 16448 23060 16454 23112
rect 18509 23103 18567 23109
rect 18509 23069 18521 23103
rect 18555 23069 18567 23103
rect 18509 23063 18567 23069
rect 18601 23103 18659 23109
rect 18601 23069 18613 23103
rect 18647 23100 18659 23103
rect 19444 23100 19472 23199
rect 25222 23196 25228 23248
rect 25280 23236 25286 23248
rect 26142 23236 26148 23248
rect 25280 23208 26148 23236
rect 25280 23196 25286 23208
rect 19978 23168 19984 23180
rect 19939 23140 19984 23168
rect 19978 23128 19984 23140
rect 20036 23128 20042 23180
rect 21450 23168 21456 23180
rect 21411 23140 21456 23168
rect 21450 23128 21456 23140
rect 21508 23128 21514 23180
rect 25038 23128 25044 23180
rect 25096 23168 25102 23180
rect 25096 23140 25452 23168
rect 25096 23128 25102 23140
rect 18647 23072 19472 23100
rect 18647 23069 18659 23072
rect 18601 23063 18659 23069
rect 18524 23032 18552 23063
rect 19610 23060 19616 23112
rect 19668 23100 19674 23112
rect 19797 23103 19855 23109
rect 19797 23100 19809 23103
rect 19668 23072 19809 23100
rect 19668 23060 19674 23072
rect 19797 23069 19809 23072
rect 19843 23069 19855 23103
rect 19797 23063 19855 23069
rect 19889 23103 19947 23109
rect 19889 23069 19901 23103
rect 19935 23100 19947 23103
rect 20070 23100 20076 23112
rect 19935 23072 20076 23100
rect 19935 23069 19947 23072
rect 19889 23063 19947 23069
rect 20070 23060 20076 23072
rect 20128 23060 20134 23112
rect 20990 23060 20996 23112
rect 21048 23100 21054 23112
rect 21177 23103 21235 23109
rect 21177 23100 21189 23103
rect 21048 23072 21189 23100
rect 21048 23060 21054 23072
rect 21177 23069 21189 23072
rect 21223 23069 21235 23103
rect 21177 23063 21235 23069
rect 25130 23060 25136 23112
rect 25188 23100 25194 23112
rect 25424 23109 25452 23140
rect 25516 23109 25544 23208
rect 26142 23196 26148 23208
rect 26200 23196 26206 23248
rect 27430 23236 27436 23248
rect 26528 23208 27436 23236
rect 26528 23177 26556 23208
rect 27430 23196 27436 23208
rect 27488 23196 27494 23248
rect 26513 23171 26571 23177
rect 26513 23137 26525 23171
rect 26559 23137 26571 23171
rect 26694 23168 26700 23180
rect 26655 23140 26700 23168
rect 26513 23131 26571 23137
rect 26694 23128 26700 23140
rect 26752 23128 26758 23180
rect 28353 23171 28411 23177
rect 28353 23137 28365 23171
rect 28399 23168 28411 23171
rect 29914 23168 29920 23180
rect 28399 23140 29920 23168
rect 28399 23137 28411 23140
rect 28353 23131 28411 23137
rect 29914 23128 29920 23140
rect 29972 23128 29978 23180
rect 25225 23103 25283 23109
rect 25225 23100 25237 23103
rect 25188 23072 25237 23100
rect 25188 23060 25194 23072
rect 25225 23069 25237 23072
rect 25271 23069 25283 23103
rect 25225 23063 25283 23069
rect 25409 23103 25467 23109
rect 25409 23069 25421 23103
rect 25455 23069 25467 23103
rect 25409 23063 25467 23069
rect 25501 23103 25559 23109
rect 25501 23069 25513 23103
rect 25547 23069 25559 23103
rect 25501 23063 25559 23069
rect 25593 23103 25651 23109
rect 25593 23069 25605 23103
rect 25639 23069 25651 23103
rect 25593 23063 25651 23069
rect 18782 23032 18788 23044
rect 18524 23004 18788 23032
rect 18782 22992 18788 23004
rect 18840 23032 18846 23044
rect 19702 23032 19708 23044
rect 18840 23004 19708 23032
rect 18840 22992 18846 23004
rect 19702 22992 19708 23004
rect 19760 22992 19766 23044
rect 24302 22992 24308 23044
rect 24360 23032 24366 23044
rect 25608 23032 25636 23063
rect 24360 23004 25636 23032
rect 24360 22992 24366 23004
rect 16574 22964 16580 22976
rect 16535 22936 16580 22964
rect 16574 22924 16580 22936
rect 16632 22924 16638 22976
rect 25866 22964 25872 22976
rect 25827 22936 25872 22964
rect 25866 22924 25872 22936
rect 25924 22924 25930 22976
rect 1104 22874 29048 22896
rect 1104 22822 7896 22874
rect 7948 22822 7960 22874
rect 8012 22822 8024 22874
rect 8076 22822 8088 22874
rect 8140 22822 8152 22874
rect 8204 22822 14842 22874
rect 14894 22822 14906 22874
rect 14958 22822 14970 22874
rect 15022 22822 15034 22874
rect 15086 22822 15098 22874
rect 15150 22822 21788 22874
rect 21840 22822 21852 22874
rect 21904 22822 21916 22874
rect 21968 22822 21980 22874
rect 22032 22822 22044 22874
rect 22096 22822 28734 22874
rect 28786 22822 28798 22874
rect 28850 22822 28862 22874
rect 28914 22822 28926 22874
rect 28978 22822 28990 22874
rect 29042 22822 29048 22874
rect 1104 22800 29048 22822
rect 15749 22763 15807 22769
rect 15749 22729 15761 22763
rect 15795 22760 15807 22763
rect 18138 22760 18144 22772
rect 15795 22732 18144 22760
rect 15795 22729 15807 22732
rect 15749 22723 15807 22729
rect 18138 22720 18144 22732
rect 18196 22760 18202 22772
rect 18233 22763 18291 22769
rect 18233 22760 18245 22763
rect 18196 22732 18245 22760
rect 18196 22720 18202 22732
rect 18233 22729 18245 22732
rect 18279 22729 18291 22763
rect 18233 22723 18291 22729
rect 20530 22720 20536 22772
rect 20588 22760 20594 22772
rect 22173 22763 22231 22769
rect 22173 22760 22185 22763
rect 20588 22732 22185 22760
rect 20588 22720 20594 22732
rect 22173 22729 22185 22732
rect 22219 22760 22231 22763
rect 24026 22760 24032 22772
rect 22219 22732 24032 22760
rect 22219 22729 22231 22732
rect 22173 22723 22231 22729
rect 24026 22720 24032 22732
rect 24084 22720 24090 22772
rect 24581 22763 24639 22769
rect 24581 22729 24593 22763
rect 24627 22760 24639 22763
rect 24762 22760 24768 22772
rect 24627 22732 24768 22760
rect 24627 22729 24639 22732
rect 24581 22723 24639 22729
rect 24762 22720 24768 22732
rect 24820 22720 24826 22772
rect 26418 22720 26424 22772
rect 26476 22760 26482 22772
rect 26605 22763 26663 22769
rect 26605 22760 26617 22763
rect 26476 22732 26617 22760
rect 26476 22720 26482 22732
rect 26605 22729 26617 22732
rect 26651 22729 26663 22763
rect 27338 22760 27344 22772
rect 27299 22732 27344 22760
rect 26605 22723 26663 22729
rect 27338 22720 27344 22732
rect 27396 22720 27402 22772
rect 16574 22652 16580 22704
rect 16632 22692 16638 22704
rect 17098 22695 17156 22701
rect 17098 22692 17110 22695
rect 16632 22664 17110 22692
rect 16632 22652 16638 22664
rect 17098 22661 17110 22664
rect 17144 22661 17156 22695
rect 22370 22692 22376 22704
rect 22331 22664 22376 22692
rect 17098 22655 17156 22661
rect 22370 22652 22376 22664
rect 22428 22652 22434 22704
rect 24210 22692 24216 22704
rect 24171 22664 24216 22692
rect 24210 22652 24216 22664
rect 24268 22652 24274 22704
rect 24413 22695 24471 22701
rect 24413 22692 24425 22695
rect 24412 22661 24425 22692
rect 24459 22661 24471 22695
rect 24412 22655 24471 22661
rect 25492 22695 25550 22701
rect 25492 22661 25504 22695
rect 25538 22692 25550 22695
rect 25866 22692 25872 22704
rect 25538 22664 25872 22692
rect 25538 22661 25550 22664
rect 25492 22655 25550 22661
rect 15657 22627 15715 22633
rect 15657 22624 15669 22627
rect 6886 22596 15669 22624
rect 1854 22516 1860 22568
rect 1912 22556 1918 22568
rect 6886 22556 6914 22596
rect 15657 22593 15669 22596
rect 15703 22593 15715 22627
rect 15657 22587 15715 22593
rect 23658 22584 23664 22636
rect 23716 22624 23722 22636
rect 24412 22624 24440 22655
rect 25866 22652 25872 22664
rect 25924 22652 25930 22704
rect 23716 22596 24440 22624
rect 23716 22584 23722 22596
rect 27246 22584 27252 22636
rect 27304 22624 27310 22636
rect 27433 22627 27491 22633
rect 27433 22624 27445 22627
rect 27304 22596 27445 22624
rect 27304 22584 27310 22596
rect 27433 22593 27445 22596
rect 27479 22593 27491 22627
rect 27890 22624 27896 22636
rect 27851 22596 27896 22624
rect 27433 22587 27491 22593
rect 27890 22584 27896 22596
rect 27948 22584 27954 22636
rect 1912 22528 6914 22556
rect 1912 22516 1918 22528
rect 15378 22516 15384 22568
rect 15436 22556 15442 22568
rect 15473 22559 15531 22565
rect 15473 22556 15485 22559
rect 15436 22528 15485 22556
rect 15436 22516 15442 22528
rect 15473 22525 15485 22528
rect 15519 22556 15531 22559
rect 16666 22556 16672 22568
rect 15519 22528 16672 22556
rect 15519 22525 15531 22528
rect 15473 22519 15531 22525
rect 16666 22516 16672 22528
rect 16724 22516 16730 22568
rect 16758 22516 16764 22568
rect 16816 22556 16822 22568
rect 16853 22559 16911 22565
rect 16853 22556 16865 22559
rect 16816 22528 16865 22556
rect 16816 22516 16822 22528
rect 16853 22525 16865 22528
rect 16899 22525 16911 22559
rect 16853 22519 16911 22525
rect 25038 22516 25044 22568
rect 25096 22556 25102 22568
rect 25225 22559 25283 22565
rect 25225 22556 25237 22559
rect 25096 22528 25237 22556
rect 25096 22516 25102 22528
rect 25225 22525 25237 22528
rect 25271 22525 25283 22559
rect 25225 22519 25283 22525
rect 23934 22448 23940 22500
rect 23992 22488 23998 22500
rect 23992 22460 24440 22488
rect 23992 22448 23998 22460
rect 24412 22432 24440 22460
rect 16114 22420 16120 22432
rect 16075 22392 16120 22420
rect 16114 22380 16120 22392
rect 16172 22380 16178 22432
rect 21266 22380 21272 22432
rect 21324 22420 21330 22432
rect 22005 22423 22063 22429
rect 22005 22420 22017 22423
rect 21324 22392 22017 22420
rect 21324 22380 21330 22392
rect 22005 22389 22017 22392
rect 22051 22389 22063 22423
rect 22005 22383 22063 22389
rect 22189 22423 22247 22429
rect 22189 22389 22201 22423
rect 22235 22420 22247 22423
rect 24302 22420 24308 22432
rect 22235 22392 24308 22420
rect 22235 22389 22247 22392
rect 22189 22383 22247 22389
rect 24302 22380 24308 22392
rect 24360 22380 24366 22432
rect 24394 22380 24400 22432
rect 24452 22420 24458 22432
rect 24452 22392 24497 22420
rect 24452 22380 24458 22392
rect 1104 22330 28888 22352
rect 1104 22278 4423 22330
rect 4475 22278 4487 22330
rect 4539 22278 4551 22330
rect 4603 22278 4615 22330
rect 4667 22278 4679 22330
rect 4731 22278 11369 22330
rect 11421 22278 11433 22330
rect 11485 22278 11497 22330
rect 11549 22278 11561 22330
rect 11613 22278 11625 22330
rect 11677 22278 18315 22330
rect 18367 22278 18379 22330
rect 18431 22278 18443 22330
rect 18495 22278 18507 22330
rect 18559 22278 18571 22330
rect 18623 22278 25261 22330
rect 25313 22278 25325 22330
rect 25377 22278 25389 22330
rect 25441 22278 25453 22330
rect 25505 22278 25517 22330
rect 25569 22278 28888 22330
rect 1104 22256 28888 22278
rect 15749 22219 15807 22225
rect 15749 22185 15761 22219
rect 15795 22216 15807 22219
rect 16390 22216 16396 22228
rect 15795 22188 16396 22216
rect 15795 22185 15807 22188
rect 15749 22179 15807 22185
rect 16390 22176 16396 22188
rect 16448 22176 16454 22228
rect 22370 22176 22376 22228
rect 22428 22216 22434 22228
rect 22925 22219 22983 22225
rect 22925 22216 22937 22219
rect 22428 22188 22937 22216
rect 22428 22176 22434 22188
rect 22925 22185 22937 22188
rect 22971 22185 22983 22219
rect 22925 22179 22983 22185
rect 23937 22219 23995 22225
rect 23937 22185 23949 22219
rect 23983 22216 23995 22219
rect 23983 22188 24992 22216
rect 23983 22185 23995 22188
rect 23937 22179 23995 22185
rect 24964 22157 24992 22188
rect 24949 22151 25007 22157
rect 24949 22117 24961 22151
rect 24995 22117 25007 22151
rect 24949 22111 25007 22117
rect 24854 22080 24860 22092
rect 24815 22052 24860 22080
rect 24854 22040 24860 22052
rect 24912 22040 24918 22092
rect 25958 22080 25964 22092
rect 24964 22052 25964 22080
rect 16114 22012 16120 22024
rect 16075 21984 16120 22012
rect 16114 21972 16120 21984
rect 16172 21972 16178 22024
rect 16574 22012 16580 22024
rect 16535 21984 16580 22012
rect 16574 21972 16580 21984
rect 16632 21972 16638 22024
rect 19702 21972 19708 22024
rect 19760 22012 19766 22024
rect 20901 22015 20959 22021
rect 20901 22012 20913 22015
rect 19760 21984 20913 22012
rect 19760 21972 19766 21984
rect 20901 21981 20913 21984
rect 20947 21981 20959 22015
rect 20901 21975 20959 21981
rect 21361 22015 21419 22021
rect 21361 21981 21373 22015
rect 21407 22012 21419 22015
rect 21450 22012 21456 22024
rect 21407 21984 21456 22012
rect 21407 21981 21419 21984
rect 21361 21975 21419 21981
rect 21450 21972 21456 21984
rect 21508 21972 21514 22024
rect 23658 22012 23664 22024
rect 23619 21984 23664 22012
rect 23658 21972 23664 21984
rect 23716 21972 23722 22024
rect 24578 22012 24584 22024
rect 24539 21984 24584 22012
rect 24578 21972 24584 21984
rect 24636 21972 24642 22024
rect 24765 22015 24823 22021
rect 24765 22012 24777 22015
rect 24688 21984 24777 22012
rect 15933 21947 15991 21953
rect 15933 21913 15945 21947
rect 15979 21944 15991 21947
rect 16206 21944 16212 21956
rect 15979 21916 16212 21944
rect 15979 21913 15991 21916
rect 15933 21907 15991 21913
rect 16206 21904 16212 21916
rect 16264 21904 16270 21956
rect 22893 21947 22951 21953
rect 22893 21944 22905 21947
rect 22296 21916 22905 21944
rect 22296 21888 22324 21916
rect 22893 21913 22905 21916
rect 22939 21913 22951 21947
rect 22893 21907 22951 21913
rect 23109 21947 23167 21953
rect 23109 21913 23121 21947
rect 23155 21913 23167 21947
rect 23934 21944 23940 21956
rect 23895 21916 23940 21944
rect 23109 21907 23167 21913
rect 16761 21879 16819 21885
rect 16761 21845 16773 21879
rect 16807 21876 16819 21879
rect 16942 21876 16948 21888
rect 16807 21848 16948 21876
rect 16807 21845 16819 21848
rect 16761 21839 16819 21845
rect 16942 21836 16948 21848
rect 17000 21836 17006 21888
rect 21174 21876 21180 21888
rect 21135 21848 21180 21876
rect 21174 21836 21180 21848
rect 21232 21836 21238 21888
rect 21269 21879 21327 21885
rect 21269 21845 21281 21879
rect 21315 21876 21327 21879
rect 21358 21876 21364 21888
rect 21315 21848 21364 21876
rect 21315 21845 21327 21848
rect 21269 21839 21327 21845
rect 21358 21836 21364 21848
rect 21416 21876 21422 21888
rect 22278 21876 22284 21888
rect 21416 21848 22284 21876
rect 21416 21836 21422 21848
rect 22278 21836 22284 21848
rect 22336 21836 22342 21888
rect 22738 21876 22744 21888
rect 22699 21848 22744 21876
rect 22738 21836 22744 21848
rect 22796 21836 22802 21888
rect 23124 21876 23152 21907
rect 23934 21904 23940 21916
rect 23992 21904 23998 21956
rect 24486 21904 24492 21956
rect 24544 21944 24550 21956
rect 24688 21944 24716 21984
rect 24765 21981 24777 21984
rect 24811 22012 24823 22015
rect 24964 22012 24992 22052
rect 25958 22040 25964 22052
rect 26016 22040 26022 22092
rect 27522 22080 27528 22092
rect 27483 22052 27528 22080
rect 27522 22040 27528 22052
rect 27580 22040 27586 22092
rect 24811 21984 24992 22012
rect 25041 22015 25099 22021
rect 24811 21981 24823 21984
rect 24765 21975 24823 21981
rect 25041 21981 25053 22015
rect 25087 21981 25099 22015
rect 25041 21975 25099 21981
rect 25056 21944 25084 21975
rect 28350 21972 28356 22024
rect 28408 22012 28414 22024
rect 28408 21984 28453 22012
rect 28408 21972 28414 21984
rect 28166 21944 28172 21956
rect 24544 21916 24716 21944
rect 24780 21916 25084 21944
rect 28127 21916 28172 21944
rect 24544 21904 24550 21916
rect 24780 21888 24808 21916
rect 28166 21904 28172 21916
rect 28224 21904 28230 21956
rect 23750 21876 23756 21888
rect 23124 21848 23756 21876
rect 23750 21836 23756 21848
rect 23808 21876 23814 21888
rect 24210 21876 24216 21888
rect 23808 21848 24216 21876
rect 23808 21836 23814 21848
rect 24210 21836 24216 21848
rect 24268 21836 24274 21888
rect 24762 21836 24768 21888
rect 24820 21836 24826 21888
rect 25130 21836 25136 21888
rect 25188 21876 25194 21888
rect 25225 21879 25283 21885
rect 25225 21876 25237 21879
rect 25188 21848 25237 21876
rect 25188 21836 25194 21848
rect 25225 21845 25237 21848
rect 25271 21845 25283 21879
rect 25225 21839 25283 21845
rect 1104 21786 29048 21808
rect 1104 21734 7896 21786
rect 7948 21734 7960 21786
rect 8012 21734 8024 21786
rect 8076 21734 8088 21786
rect 8140 21734 8152 21786
rect 8204 21734 14842 21786
rect 14894 21734 14906 21786
rect 14958 21734 14970 21786
rect 15022 21734 15034 21786
rect 15086 21734 15098 21786
rect 15150 21734 21788 21786
rect 21840 21734 21852 21786
rect 21904 21734 21916 21786
rect 21968 21734 21980 21786
rect 22032 21734 22044 21786
rect 22096 21734 28734 21786
rect 28786 21734 28798 21786
rect 28850 21734 28862 21786
rect 28914 21734 28926 21786
rect 28978 21734 28990 21786
rect 29042 21734 29048 21786
rect 1104 21712 29048 21734
rect 15933 21675 15991 21681
rect 15933 21641 15945 21675
rect 15979 21672 15991 21675
rect 18233 21675 18291 21681
rect 18233 21672 18245 21675
rect 15979 21644 18245 21672
rect 15979 21641 15991 21644
rect 15933 21635 15991 21641
rect 18233 21641 18245 21644
rect 18279 21672 18291 21675
rect 19058 21672 19064 21684
rect 18279 21644 19064 21672
rect 18279 21641 18291 21644
rect 18233 21635 18291 21641
rect 19058 21632 19064 21644
rect 19116 21632 19122 21684
rect 28166 21672 28172 21684
rect 28127 21644 28172 21672
rect 28166 21632 28172 21644
rect 28224 21632 28230 21684
rect 21082 21604 21088 21616
rect 16868 21576 21088 21604
rect 15194 21496 15200 21548
rect 15252 21536 15258 21548
rect 15841 21539 15899 21545
rect 15841 21536 15853 21539
rect 15252 21508 15853 21536
rect 15252 21496 15258 21508
rect 15841 21505 15853 21508
rect 15887 21505 15899 21539
rect 15841 21499 15899 21505
rect 16758 21496 16764 21548
rect 16816 21536 16822 21548
rect 16868 21545 16896 21576
rect 16853 21539 16911 21545
rect 16853 21536 16865 21539
rect 16816 21508 16865 21536
rect 16816 21496 16822 21508
rect 16853 21505 16865 21508
rect 16899 21505 16911 21539
rect 16853 21499 16911 21505
rect 16942 21496 16948 21548
rect 17000 21536 17006 21548
rect 18708 21545 18736 21576
rect 21082 21564 21088 21576
rect 21140 21564 21146 21616
rect 28350 21604 28356 21616
rect 27632 21576 28356 21604
rect 18966 21545 18972 21548
rect 17109 21539 17167 21545
rect 17109 21536 17121 21539
rect 17000 21508 17121 21536
rect 17000 21496 17006 21508
rect 17109 21505 17121 21508
rect 17155 21505 17167 21539
rect 17109 21499 17167 21505
rect 18693 21539 18751 21545
rect 18693 21505 18705 21539
rect 18739 21505 18751 21539
rect 18693 21499 18751 21505
rect 18960 21499 18972 21545
rect 19024 21536 19030 21548
rect 20990 21536 20996 21548
rect 19024 21508 19060 21536
rect 20951 21508 20996 21536
rect 18966 21496 18972 21499
rect 19024 21496 19030 21508
rect 20990 21496 20996 21508
rect 21048 21496 21054 21548
rect 21174 21496 21180 21548
rect 21232 21536 21238 21548
rect 21269 21539 21327 21545
rect 21269 21536 21281 21539
rect 21232 21508 21281 21536
rect 21232 21496 21238 21508
rect 21269 21505 21281 21508
rect 21315 21505 21327 21539
rect 21269 21499 21327 21505
rect 22557 21539 22615 21545
rect 22557 21505 22569 21539
rect 22603 21505 22615 21539
rect 22738 21536 22744 21548
rect 22699 21508 22744 21536
rect 22557 21499 22615 21505
rect 15654 21428 15660 21480
rect 15712 21468 15718 21480
rect 15749 21471 15807 21477
rect 15749 21468 15761 21471
rect 15712 21440 15761 21468
rect 15712 21428 15718 21440
rect 15749 21437 15761 21440
rect 15795 21437 15807 21471
rect 21008 21468 21036 21496
rect 21008 21440 22094 21468
rect 15749 21431 15807 21437
rect 15764 21400 15792 21431
rect 16850 21400 16856 21412
rect 15764 21372 16856 21400
rect 16850 21360 16856 21372
rect 16908 21360 16914 21412
rect 21177 21403 21235 21409
rect 21177 21369 21189 21403
rect 21223 21400 21235 21403
rect 21266 21400 21272 21412
rect 21223 21372 21272 21400
rect 21223 21369 21235 21372
rect 21177 21363 21235 21369
rect 21266 21360 21272 21372
rect 21324 21360 21330 21412
rect 22066 21400 22094 21440
rect 22572 21400 22600 21499
rect 22738 21496 22744 21508
rect 22796 21496 22802 21548
rect 25130 21536 25136 21548
rect 25091 21508 25136 21536
rect 25130 21496 25136 21508
rect 25188 21496 25194 21548
rect 25222 21496 25228 21548
rect 25280 21536 25286 21548
rect 25317 21539 25375 21545
rect 25317 21536 25329 21539
rect 25280 21508 25329 21536
rect 25280 21496 25286 21508
rect 25317 21505 25329 21508
rect 25363 21536 25375 21539
rect 25682 21536 25688 21548
rect 25363 21508 25688 21536
rect 25363 21505 25375 21508
rect 25317 21499 25375 21505
rect 25682 21496 25688 21508
rect 25740 21496 25746 21548
rect 27632 21545 27660 21576
rect 28350 21564 28356 21576
rect 28408 21564 28414 21616
rect 27617 21539 27675 21545
rect 27617 21505 27629 21539
rect 27663 21505 27675 21539
rect 27617 21499 27675 21505
rect 28077 21539 28135 21545
rect 28077 21505 28089 21539
rect 28123 21536 28135 21539
rect 28258 21536 28264 21548
rect 28123 21508 28264 21536
rect 28123 21505 28135 21508
rect 28077 21499 28135 21505
rect 22830 21468 22836 21480
rect 22791 21440 22836 21468
rect 22830 21428 22836 21440
rect 22888 21428 22894 21480
rect 28092 21468 28120 21499
rect 28258 21496 28264 21508
rect 28316 21496 28322 21548
rect 27632 21440 28120 21468
rect 27632 21412 27660 21440
rect 24946 21400 24952 21412
rect 22066 21372 24952 21400
rect 24946 21360 24952 21372
rect 25004 21360 25010 21412
rect 27614 21360 27620 21412
rect 27672 21360 27678 21412
rect 16298 21332 16304 21344
rect 16259 21304 16304 21332
rect 16298 21292 16304 21304
rect 16356 21292 16362 21344
rect 20070 21332 20076 21344
rect 20031 21304 20076 21332
rect 20070 21292 20076 21304
rect 20128 21292 20134 21344
rect 20806 21332 20812 21344
rect 20767 21304 20812 21332
rect 20806 21292 20812 21304
rect 20864 21292 20870 21344
rect 22370 21332 22376 21344
rect 22331 21304 22376 21332
rect 22370 21292 22376 21304
rect 22428 21292 22434 21344
rect 25225 21335 25283 21341
rect 25225 21301 25237 21335
rect 25271 21332 25283 21335
rect 25590 21332 25596 21344
rect 25271 21304 25596 21332
rect 25271 21301 25283 21304
rect 25225 21295 25283 21301
rect 25590 21292 25596 21304
rect 25648 21292 25654 21344
rect 1104 21242 28888 21264
rect 1104 21190 4423 21242
rect 4475 21190 4487 21242
rect 4539 21190 4551 21242
rect 4603 21190 4615 21242
rect 4667 21190 4679 21242
rect 4731 21190 11369 21242
rect 11421 21190 11433 21242
rect 11485 21190 11497 21242
rect 11549 21190 11561 21242
rect 11613 21190 11625 21242
rect 11677 21190 18315 21242
rect 18367 21190 18379 21242
rect 18431 21190 18443 21242
rect 18495 21190 18507 21242
rect 18559 21190 18571 21242
rect 18623 21190 25261 21242
rect 25313 21190 25325 21242
rect 25377 21190 25389 21242
rect 25441 21190 25453 21242
rect 25505 21190 25517 21242
rect 25569 21190 28888 21242
rect 1104 21168 28888 21190
rect 14734 21088 14740 21140
rect 14792 21128 14798 21140
rect 15013 21131 15071 21137
rect 15013 21128 15025 21131
rect 14792 21100 15025 21128
rect 14792 21088 14798 21100
rect 15013 21097 15025 21100
rect 15059 21097 15071 21131
rect 15013 21091 15071 21097
rect 15933 21131 15991 21137
rect 15933 21097 15945 21131
rect 15979 21128 15991 21131
rect 16574 21128 16580 21140
rect 15979 21100 16580 21128
rect 15979 21097 15991 21100
rect 15933 21091 15991 21097
rect 16574 21088 16580 21100
rect 16632 21088 16638 21140
rect 19702 21128 19708 21140
rect 19663 21100 19708 21128
rect 19702 21088 19708 21100
rect 19760 21088 19766 21140
rect 18509 20995 18567 21001
rect 18509 20961 18521 20995
rect 18555 20992 18567 20995
rect 18782 20992 18788 21004
rect 18555 20964 18788 20992
rect 18555 20961 18567 20964
rect 18509 20955 18567 20961
rect 18782 20952 18788 20964
rect 18840 20952 18846 21004
rect 21082 20992 21088 21004
rect 21043 20964 21088 20992
rect 21082 20952 21088 20964
rect 21140 20952 21146 21004
rect 21634 20952 21640 21004
rect 21692 20992 21698 21004
rect 21821 20995 21879 21001
rect 21821 20992 21833 20995
rect 21692 20964 21833 20992
rect 21692 20952 21698 20964
rect 21821 20961 21833 20964
rect 21867 20961 21879 20995
rect 27522 20992 27528 21004
rect 27483 20964 27528 20992
rect 21821 20955 21879 20961
rect 27522 20952 27528 20964
rect 27580 20952 27586 21004
rect 16298 20924 16304 20936
rect 16259 20896 16304 20924
rect 16298 20884 16304 20896
rect 16356 20884 16362 20936
rect 18693 20927 18751 20933
rect 18693 20893 18705 20927
rect 18739 20924 18751 20927
rect 19518 20924 19524 20936
rect 18739 20896 19524 20924
rect 18739 20893 18751 20896
rect 18693 20887 18751 20893
rect 19518 20884 19524 20896
rect 19576 20884 19582 20936
rect 20806 20884 20812 20936
rect 20864 20933 20870 20936
rect 20864 20924 20876 20933
rect 22088 20927 22146 20933
rect 20864 20896 20909 20924
rect 20864 20887 20876 20896
rect 22088 20893 22100 20927
rect 22134 20924 22146 20927
rect 22370 20924 22376 20936
rect 22134 20896 22376 20924
rect 22134 20893 22146 20896
rect 22088 20887 22146 20893
rect 20864 20884 20870 20887
rect 22370 20884 22376 20896
rect 22428 20884 22434 20936
rect 24946 20884 24952 20936
rect 25004 20924 25010 20936
rect 25409 20927 25467 20933
rect 25409 20924 25421 20927
rect 25004 20896 25421 20924
rect 25004 20884 25010 20896
rect 25409 20893 25421 20896
rect 25455 20893 25467 20927
rect 25590 20924 25596 20936
rect 25551 20896 25596 20924
rect 25409 20887 25467 20893
rect 25590 20884 25596 20896
rect 25648 20884 25654 20936
rect 25682 20884 25688 20936
rect 25740 20924 25746 20936
rect 25823 20927 25881 20933
rect 25740 20896 25785 20924
rect 25740 20884 25746 20896
rect 25823 20893 25835 20927
rect 25869 20924 25881 20927
rect 25958 20924 25964 20936
rect 25869 20896 25964 20924
rect 25869 20893 25881 20896
rect 25823 20887 25881 20893
rect 25958 20884 25964 20896
rect 26016 20884 26022 20936
rect 28350 20884 28356 20936
rect 28408 20924 28414 20936
rect 28408 20896 28453 20924
rect 28408 20884 28414 20896
rect 14734 20816 14740 20868
rect 14792 20856 14798 20868
rect 15197 20859 15255 20865
rect 15197 20856 15209 20859
rect 14792 20828 15209 20856
rect 14792 20816 14798 20828
rect 15197 20825 15209 20828
rect 15243 20825 15255 20859
rect 15378 20856 15384 20868
rect 15339 20828 15384 20856
rect 15197 20819 15255 20825
rect 15378 20816 15384 20828
rect 15436 20816 15442 20868
rect 16117 20859 16175 20865
rect 16117 20825 16129 20859
rect 16163 20856 16175 20859
rect 16206 20856 16212 20868
rect 16163 20828 16212 20856
rect 16163 20825 16175 20828
rect 16117 20819 16175 20825
rect 16206 20816 16212 20828
rect 16264 20816 16270 20868
rect 28166 20856 28172 20868
rect 28127 20828 28172 20856
rect 28166 20816 28172 20828
rect 28224 20816 28230 20868
rect 18690 20748 18696 20800
rect 18748 20788 18754 20800
rect 18877 20791 18935 20797
rect 18877 20788 18889 20791
rect 18748 20760 18889 20788
rect 18748 20748 18754 20760
rect 18877 20757 18889 20760
rect 18923 20757 18935 20791
rect 18877 20751 18935 20757
rect 22462 20748 22468 20800
rect 22520 20788 22526 20800
rect 23201 20791 23259 20797
rect 23201 20788 23213 20791
rect 22520 20760 23213 20788
rect 22520 20748 22526 20760
rect 23201 20757 23213 20760
rect 23247 20757 23259 20791
rect 26050 20788 26056 20800
rect 26011 20760 26056 20788
rect 23201 20751 23259 20757
rect 26050 20748 26056 20760
rect 26108 20748 26114 20800
rect 1104 20698 29048 20720
rect 1104 20646 7896 20698
rect 7948 20646 7960 20698
rect 8012 20646 8024 20698
rect 8076 20646 8088 20698
rect 8140 20646 8152 20698
rect 8204 20646 14842 20698
rect 14894 20646 14906 20698
rect 14958 20646 14970 20698
rect 15022 20646 15034 20698
rect 15086 20646 15098 20698
rect 15150 20646 21788 20698
rect 21840 20646 21852 20698
rect 21904 20646 21916 20698
rect 21968 20646 21980 20698
rect 22032 20646 22044 20698
rect 22096 20646 28734 20698
rect 28786 20646 28798 20698
rect 28850 20646 28862 20698
rect 28914 20646 28926 20698
rect 28978 20646 28990 20698
rect 29042 20646 29048 20698
rect 1104 20624 29048 20646
rect 12618 20584 12624 20596
rect 12579 20556 12624 20584
rect 12618 20544 12624 20556
rect 12676 20544 12682 20596
rect 18877 20587 18935 20593
rect 18877 20553 18889 20587
rect 18923 20584 18935 20587
rect 18966 20584 18972 20596
rect 18923 20556 18972 20584
rect 18923 20553 18935 20556
rect 18877 20547 18935 20553
rect 18966 20544 18972 20556
rect 19024 20544 19030 20596
rect 19518 20584 19524 20596
rect 19479 20556 19524 20584
rect 19518 20544 19524 20556
rect 19576 20544 19582 20596
rect 19794 20544 19800 20596
rect 19852 20584 19858 20596
rect 19889 20587 19947 20593
rect 19889 20584 19901 20587
rect 19852 20556 19901 20584
rect 19852 20544 19858 20556
rect 19889 20553 19901 20556
rect 19935 20584 19947 20587
rect 20070 20584 20076 20596
rect 19935 20556 20076 20584
rect 19935 20553 19947 20556
rect 19889 20547 19947 20553
rect 20070 20544 20076 20556
rect 20128 20544 20134 20596
rect 22465 20587 22523 20593
rect 22465 20553 22477 20587
rect 22511 20584 22523 20587
rect 22830 20584 22836 20596
rect 22511 20556 22836 20584
rect 22511 20553 22523 20556
rect 22465 20547 22523 20553
rect 22830 20544 22836 20556
rect 22888 20544 22894 20596
rect 24670 20544 24676 20596
rect 24728 20584 24734 20596
rect 28166 20584 28172 20596
rect 24728 20556 25820 20584
rect 28127 20556 28172 20584
rect 24728 20544 24734 20556
rect 14458 20476 14464 20528
rect 14516 20516 14522 20528
rect 14737 20519 14795 20525
rect 14737 20516 14749 20519
rect 14516 20488 14749 20516
rect 14516 20476 14522 20488
rect 14737 20485 14749 20488
rect 14783 20485 14795 20519
rect 14737 20479 14795 20485
rect 19702 20476 19708 20528
rect 19760 20516 19766 20528
rect 19981 20519 20039 20525
rect 19981 20516 19993 20519
rect 19760 20488 19993 20516
rect 19760 20476 19766 20488
rect 19981 20485 19993 20488
rect 20027 20485 20039 20519
rect 23658 20516 23664 20528
rect 23571 20488 23664 20516
rect 19981 20479 20039 20485
rect 23658 20476 23664 20488
rect 23716 20516 23722 20528
rect 24688 20516 24716 20544
rect 23716 20488 24716 20516
rect 23716 20476 23722 20488
rect 24946 20476 24952 20528
rect 25004 20516 25010 20528
rect 25682 20516 25688 20528
rect 25004 20488 25084 20516
rect 25004 20476 25010 20488
rect 2498 20448 2504 20460
rect 2459 20420 2504 20448
rect 2498 20408 2504 20420
rect 2556 20408 2562 20460
rect 12805 20451 12863 20457
rect 12805 20417 12817 20451
rect 12851 20417 12863 20451
rect 12986 20448 12992 20460
rect 12947 20420 12992 20448
rect 12805 20411 12863 20417
rect 12820 20380 12848 20411
rect 12986 20408 12992 20420
rect 13044 20408 13050 20460
rect 13078 20408 13084 20460
rect 13136 20448 13142 20460
rect 14642 20448 14648 20460
rect 13136 20420 13181 20448
rect 14603 20420 14648 20448
rect 13136 20408 13142 20420
rect 14642 20408 14648 20420
rect 14700 20408 14706 20460
rect 14826 20408 14832 20460
rect 14884 20448 14890 20460
rect 14921 20451 14979 20457
rect 14921 20448 14933 20451
rect 14884 20420 14933 20448
rect 14884 20408 14890 20420
rect 14921 20417 14933 20420
rect 14967 20417 14979 20451
rect 18690 20448 18696 20460
rect 18651 20420 18696 20448
rect 14921 20411 14979 20417
rect 18690 20408 18696 20420
rect 18748 20408 18754 20460
rect 21450 20408 21456 20460
rect 21508 20448 21514 20460
rect 22281 20451 22339 20457
rect 22281 20448 22293 20451
rect 21508 20420 22293 20448
rect 21508 20408 21514 20420
rect 22281 20417 22293 20420
rect 22327 20417 22339 20451
rect 22281 20411 22339 20417
rect 22370 20408 22376 20460
rect 22428 20448 22434 20460
rect 22428 20420 22473 20448
rect 22428 20408 22434 20420
rect 13814 20380 13820 20392
rect 12820 20352 13820 20380
rect 13814 20340 13820 20352
rect 13872 20380 13878 20392
rect 14844 20380 14872 20408
rect 13872 20352 14872 20380
rect 13872 20340 13878 20352
rect 19978 20340 19984 20392
rect 20036 20380 20042 20392
rect 20073 20383 20131 20389
rect 20073 20380 20085 20383
rect 20036 20352 20085 20380
rect 20036 20340 20042 20352
rect 20073 20349 20085 20352
rect 20119 20349 20131 20383
rect 20073 20343 20131 20349
rect 22462 20340 22468 20392
rect 22520 20380 22526 20392
rect 23676 20389 23704 20476
rect 23753 20451 23811 20457
rect 23753 20417 23765 20451
rect 23799 20448 23811 20451
rect 23934 20448 23940 20460
rect 23799 20420 23940 20448
rect 23799 20417 23811 20420
rect 23753 20411 23811 20417
rect 23934 20408 23940 20420
rect 23992 20448 23998 20460
rect 25056 20457 25084 20488
rect 25332 20488 25688 20516
rect 25041 20451 25099 20457
rect 23992 20420 24992 20448
rect 23992 20408 23998 20420
rect 22741 20383 22799 20389
rect 22741 20380 22753 20383
rect 22520 20352 22753 20380
rect 22520 20340 22526 20352
rect 22741 20349 22753 20352
rect 22787 20349 22799 20383
rect 22741 20343 22799 20349
rect 23661 20383 23719 20389
rect 23661 20349 23673 20383
rect 23707 20349 23719 20383
rect 23661 20343 23719 20349
rect 24121 20383 24179 20389
rect 24121 20349 24133 20383
rect 24167 20380 24179 20383
rect 24578 20380 24584 20392
rect 24167 20352 24584 20380
rect 24167 20349 24179 20352
rect 24121 20343 24179 20349
rect 24578 20340 24584 20352
rect 24636 20340 24642 20392
rect 24964 20380 24992 20420
rect 25041 20417 25053 20451
rect 25087 20417 25099 20451
rect 25041 20411 25099 20417
rect 25130 20408 25136 20460
rect 25188 20448 25194 20460
rect 25332 20457 25360 20488
rect 25682 20476 25688 20488
rect 25740 20476 25746 20528
rect 25225 20451 25283 20457
rect 25225 20448 25237 20451
rect 25188 20420 25237 20448
rect 25188 20408 25194 20420
rect 25225 20417 25237 20420
rect 25271 20417 25283 20451
rect 25225 20411 25283 20417
rect 25317 20451 25375 20457
rect 25317 20417 25329 20451
rect 25363 20417 25375 20451
rect 25317 20411 25375 20417
rect 25409 20451 25467 20457
rect 25409 20417 25421 20451
rect 25455 20448 25467 20451
rect 25792 20448 25820 20556
rect 28166 20544 28172 20556
rect 28224 20544 28230 20596
rect 28074 20448 28080 20460
rect 25455 20420 25820 20448
rect 28035 20420 28080 20448
rect 25455 20417 25467 20420
rect 25409 20411 25467 20417
rect 28074 20408 28080 20420
rect 28132 20408 28138 20460
rect 25958 20380 25964 20392
rect 24964 20352 25964 20380
rect 25958 20340 25964 20352
rect 26016 20340 26022 20392
rect 27617 20383 27675 20389
rect 27617 20349 27629 20383
rect 27663 20380 27675 20383
rect 28350 20380 28356 20392
rect 27663 20352 28356 20380
rect 27663 20349 27675 20352
rect 27617 20343 27675 20349
rect 28350 20340 28356 20352
rect 28408 20340 28414 20392
rect 15105 20315 15163 20321
rect 15105 20281 15117 20315
rect 15151 20312 15163 20315
rect 26326 20312 26332 20324
rect 15151 20284 26332 20312
rect 15151 20281 15163 20284
rect 15105 20275 15163 20281
rect 26326 20272 26332 20284
rect 26384 20272 26390 20324
rect 1578 20204 1584 20256
rect 1636 20244 1642 20256
rect 1673 20247 1731 20253
rect 1673 20244 1685 20247
rect 1636 20216 1685 20244
rect 1636 20204 1642 20216
rect 1673 20213 1685 20216
rect 1719 20213 1731 20247
rect 1673 20207 1731 20213
rect 1762 20204 1768 20256
rect 1820 20244 1826 20256
rect 2409 20247 2467 20253
rect 2409 20244 2421 20247
rect 1820 20216 2421 20244
rect 1820 20204 1826 20216
rect 2409 20213 2421 20216
rect 2455 20213 2467 20247
rect 25682 20244 25688 20256
rect 25643 20216 25688 20244
rect 2409 20207 2467 20213
rect 25682 20204 25688 20216
rect 25740 20204 25746 20256
rect 1104 20154 28888 20176
rect 1104 20102 4423 20154
rect 4475 20102 4487 20154
rect 4539 20102 4551 20154
rect 4603 20102 4615 20154
rect 4667 20102 4679 20154
rect 4731 20102 11369 20154
rect 11421 20102 11433 20154
rect 11485 20102 11497 20154
rect 11549 20102 11561 20154
rect 11613 20102 11625 20154
rect 11677 20102 18315 20154
rect 18367 20102 18379 20154
rect 18431 20102 18443 20154
rect 18495 20102 18507 20154
rect 18559 20102 18571 20154
rect 18623 20102 25261 20154
rect 25313 20102 25325 20154
rect 25377 20102 25389 20154
rect 25441 20102 25453 20154
rect 25505 20102 25517 20154
rect 25569 20102 28888 20154
rect 1104 20080 28888 20102
rect 13078 20000 13084 20052
rect 13136 20040 13142 20052
rect 13357 20043 13415 20049
rect 13357 20040 13369 20043
rect 13136 20012 13369 20040
rect 13136 20000 13142 20012
rect 13357 20009 13369 20012
rect 13403 20009 13415 20043
rect 14642 20040 14648 20052
rect 14603 20012 14648 20040
rect 13357 20003 13415 20009
rect 14642 20000 14648 20012
rect 14700 20000 14706 20052
rect 14734 20000 14740 20052
rect 14792 20040 14798 20052
rect 14829 20043 14887 20049
rect 14829 20040 14841 20043
rect 14792 20012 14841 20040
rect 14792 20000 14798 20012
rect 14829 20009 14841 20012
rect 14875 20009 14887 20043
rect 14829 20003 14887 20009
rect 15378 20000 15384 20052
rect 15436 20040 15442 20052
rect 15841 20043 15899 20049
rect 15841 20040 15853 20043
rect 15436 20012 15853 20040
rect 15436 20000 15442 20012
rect 15841 20009 15853 20012
rect 15887 20009 15899 20043
rect 25130 20040 25136 20052
rect 25091 20012 25136 20040
rect 15841 20003 15899 20009
rect 25130 20000 25136 20012
rect 25188 20000 25194 20052
rect 25958 20000 25964 20052
rect 26016 20040 26022 20052
rect 27157 20043 27215 20049
rect 27157 20040 27169 20043
rect 26016 20012 27169 20040
rect 26016 20000 26022 20012
rect 27157 20009 27169 20012
rect 27203 20009 27215 20043
rect 27157 20003 27215 20009
rect 1578 19904 1584 19916
rect 1539 19876 1584 19904
rect 1578 19864 1584 19876
rect 1636 19864 1642 19916
rect 1762 19904 1768 19916
rect 1723 19876 1768 19904
rect 1762 19864 1768 19876
rect 1820 19864 1826 19916
rect 2774 19904 2780 19916
rect 2735 19876 2780 19904
rect 2774 19864 2780 19876
rect 2832 19864 2838 19916
rect 23934 19864 23940 19916
rect 23992 19904 23998 19916
rect 24486 19904 24492 19916
rect 23992 19876 24492 19904
rect 23992 19864 23998 19876
rect 24486 19864 24492 19876
rect 24544 19904 24550 19916
rect 24673 19907 24731 19913
rect 24673 19904 24685 19907
rect 24544 19876 24685 19904
rect 24544 19864 24550 19876
rect 24673 19873 24685 19876
rect 24719 19873 24731 19907
rect 24673 19867 24731 19873
rect 24762 19864 24768 19916
rect 24820 19904 24826 19916
rect 24820 19876 24992 19904
rect 24820 19864 24826 19876
rect 13541 19839 13599 19845
rect 13541 19805 13553 19839
rect 13587 19836 13599 19839
rect 13722 19836 13728 19848
rect 13587 19808 13728 19836
rect 13587 19805 13599 19808
rect 13541 19799 13599 19805
rect 13722 19796 13728 19808
rect 13780 19836 13786 19848
rect 14550 19836 14556 19848
rect 13780 19808 14556 19836
rect 13780 19796 13786 19808
rect 14550 19796 14556 19808
rect 14608 19796 14614 19848
rect 14642 19796 14648 19848
rect 14700 19836 14706 19848
rect 15105 19839 15163 19845
rect 15105 19836 15117 19839
rect 14700 19808 15117 19836
rect 14700 19796 14706 19808
rect 15105 19805 15117 19808
rect 15151 19836 15163 19839
rect 15565 19839 15623 19845
rect 15565 19836 15577 19839
rect 15151 19808 15577 19836
rect 15151 19805 15163 19808
rect 15105 19799 15163 19805
rect 15565 19805 15577 19808
rect 15611 19805 15623 19839
rect 15565 19799 15623 19805
rect 16574 19796 16580 19848
rect 16632 19836 16638 19848
rect 16761 19839 16819 19845
rect 16761 19836 16773 19839
rect 16632 19808 16773 19836
rect 16632 19796 16638 19808
rect 16761 19805 16773 19808
rect 16807 19805 16819 19839
rect 16761 19799 16819 19805
rect 24581 19839 24639 19845
rect 24581 19805 24593 19839
rect 24627 19805 24639 19839
rect 24854 19836 24860 19848
rect 24815 19808 24860 19836
rect 24581 19799 24639 19805
rect 13265 19771 13323 19777
rect 13265 19737 13277 19771
rect 13311 19737 13323 19771
rect 13265 19731 13323 19737
rect 13449 19771 13507 19777
rect 13449 19737 13461 19771
rect 13495 19768 13507 19771
rect 13998 19768 14004 19780
rect 13495 19740 14004 19768
rect 13495 19737 13507 19740
rect 13449 19731 13507 19737
rect 13280 19700 13308 19731
rect 13998 19728 14004 19740
rect 14056 19728 14062 19780
rect 15841 19771 15899 19777
rect 15841 19737 15853 19771
rect 15887 19768 15899 19771
rect 15930 19768 15936 19780
rect 15887 19740 15936 19768
rect 15887 19737 15899 19740
rect 15841 19731 15899 19737
rect 15930 19728 15936 19740
rect 15988 19728 15994 19780
rect 24596 19768 24624 19799
rect 24854 19796 24860 19808
rect 24912 19796 24918 19848
rect 24964 19845 24992 19876
rect 25038 19864 25044 19916
rect 25096 19904 25102 19916
rect 25777 19907 25835 19913
rect 25777 19904 25789 19907
rect 25096 19876 25789 19904
rect 25096 19864 25102 19876
rect 25777 19873 25789 19876
rect 25823 19873 25835 19907
rect 25777 19867 25835 19873
rect 24949 19839 25007 19845
rect 24949 19805 24961 19839
rect 24995 19805 25007 19839
rect 24949 19799 25007 19805
rect 25133 19839 25191 19845
rect 25133 19805 25145 19839
rect 25179 19836 25191 19839
rect 25590 19836 25596 19848
rect 25179 19808 25596 19836
rect 25179 19805 25191 19808
rect 25133 19799 25191 19805
rect 25590 19796 25596 19808
rect 25648 19796 25654 19848
rect 26050 19845 26056 19848
rect 26044 19836 26056 19845
rect 26011 19808 26056 19836
rect 26044 19799 26056 19808
rect 26050 19796 26056 19799
rect 26108 19796 26114 19848
rect 27890 19836 27896 19848
rect 27851 19808 27896 19836
rect 27890 19796 27896 19808
rect 27948 19796 27954 19848
rect 24670 19768 24676 19780
rect 24596 19740 24676 19768
rect 24670 19728 24676 19740
rect 24728 19728 24734 19780
rect 14274 19700 14280 19712
rect 13280 19672 14280 19700
rect 14274 19660 14280 19672
rect 14332 19660 14338 19712
rect 14734 19660 14740 19712
rect 14792 19700 14798 19712
rect 15657 19703 15715 19709
rect 15657 19700 15669 19703
rect 14792 19672 15669 19700
rect 14792 19660 14798 19672
rect 15657 19669 15669 19672
rect 15703 19669 15715 19703
rect 15657 19663 15715 19669
rect 16945 19703 17003 19709
rect 16945 19669 16957 19703
rect 16991 19700 17003 19703
rect 17218 19700 17224 19712
rect 16991 19672 17224 19700
rect 16991 19669 17003 19672
rect 16945 19663 17003 19669
rect 17218 19660 17224 19672
rect 17276 19660 17282 19712
rect 1104 19610 29048 19632
rect 1104 19558 7896 19610
rect 7948 19558 7960 19610
rect 8012 19558 8024 19610
rect 8076 19558 8088 19610
rect 8140 19558 8152 19610
rect 8204 19558 14842 19610
rect 14894 19558 14906 19610
rect 14958 19558 14970 19610
rect 15022 19558 15034 19610
rect 15086 19558 15098 19610
rect 15150 19558 21788 19610
rect 21840 19558 21852 19610
rect 21904 19558 21916 19610
rect 21968 19558 21980 19610
rect 22032 19558 22044 19610
rect 22096 19558 28734 19610
rect 28786 19558 28798 19610
rect 28850 19558 28862 19610
rect 28914 19558 28926 19610
rect 28978 19558 28990 19610
rect 29042 19558 29048 19610
rect 1104 19536 29048 19558
rect 12897 19499 12955 19505
rect 12897 19465 12909 19499
rect 12943 19496 12955 19499
rect 13814 19496 13820 19508
rect 12943 19468 13820 19496
rect 12943 19465 12955 19468
rect 12897 19459 12955 19465
rect 13814 19456 13820 19468
rect 13872 19496 13878 19508
rect 14090 19496 14096 19508
rect 13872 19468 14096 19496
rect 13872 19456 13878 19468
rect 14090 19456 14096 19468
rect 14148 19456 14154 19508
rect 14458 19496 14464 19508
rect 14419 19468 14464 19496
rect 14458 19456 14464 19468
rect 14516 19456 14522 19508
rect 14734 19456 14740 19508
rect 14792 19496 14798 19508
rect 15013 19499 15071 19505
rect 15013 19496 15025 19499
rect 14792 19468 15025 19496
rect 14792 19456 14798 19468
rect 15013 19465 15025 19468
rect 15059 19465 15071 19499
rect 15013 19459 15071 19465
rect 16301 19499 16359 19505
rect 16301 19465 16313 19499
rect 16347 19496 16359 19499
rect 16942 19496 16948 19508
rect 16347 19468 16948 19496
rect 16347 19465 16359 19468
rect 16301 19459 16359 19465
rect 16942 19456 16948 19468
rect 17000 19456 17006 19508
rect 19245 19499 19303 19505
rect 19245 19496 19257 19499
rect 17052 19468 19257 19496
rect 12802 19428 12808 19440
rect 12715 19400 12808 19428
rect 12728 19369 12756 19400
rect 12802 19388 12808 19400
rect 12860 19428 12866 19440
rect 12860 19400 14412 19428
rect 12860 19388 12866 19400
rect 12713 19363 12771 19369
rect 12713 19329 12725 19363
rect 12759 19329 12771 19363
rect 13722 19360 13728 19372
rect 13683 19332 13728 19360
rect 12713 19323 12771 19329
rect 13722 19320 13728 19332
rect 13780 19320 13786 19372
rect 13909 19364 13967 19369
rect 13998 19364 14004 19372
rect 13909 19363 14004 19364
rect 13909 19329 13921 19363
rect 13955 19336 14004 19363
rect 13955 19329 13967 19336
rect 13909 19323 13967 19329
rect 13998 19320 14004 19336
rect 14056 19320 14062 19372
rect 14384 19369 14412 19400
rect 14550 19388 14556 19440
rect 14608 19428 14614 19440
rect 15657 19431 15715 19437
rect 15657 19428 15669 19431
rect 14608 19400 15669 19428
rect 14608 19388 14614 19400
rect 15657 19397 15669 19400
rect 15703 19428 15715 19431
rect 17052 19428 17080 19468
rect 19245 19465 19257 19468
rect 19291 19465 19303 19499
rect 19610 19496 19616 19508
rect 19571 19468 19616 19496
rect 19245 19459 19303 19465
rect 19610 19456 19616 19468
rect 19668 19456 19674 19508
rect 17218 19437 17224 19440
rect 17212 19428 17224 19437
rect 15703 19400 17080 19428
rect 17179 19400 17224 19428
rect 15703 19397 15715 19400
rect 15657 19391 15715 19397
rect 17212 19391 17224 19400
rect 17218 19388 17224 19391
rect 17276 19388 17282 19440
rect 14369 19363 14427 19369
rect 14369 19329 14381 19363
rect 14415 19358 14427 19363
rect 15930 19360 15936 19372
rect 14568 19358 15936 19360
rect 14415 19332 15936 19358
rect 14415 19330 14596 19332
rect 14415 19329 14427 19330
rect 14369 19323 14427 19329
rect 15930 19320 15936 19332
rect 15988 19320 15994 19372
rect 16117 19363 16175 19369
rect 16117 19329 16129 19363
rect 16163 19360 16175 19363
rect 16298 19360 16304 19372
rect 16163 19332 16304 19360
rect 16163 19329 16175 19332
rect 16117 19323 16175 19329
rect 16298 19320 16304 19332
rect 16356 19320 16362 19372
rect 16758 19320 16764 19372
rect 16816 19360 16822 19372
rect 16945 19363 17003 19369
rect 16945 19360 16957 19363
rect 16816 19332 16957 19360
rect 16816 19320 16822 19332
rect 16945 19329 16957 19332
rect 16991 19329 17003 19363
rect 16945 19323 17003 19329
rect 19334 19320 19340 19372
rect 19392 19360 19398 19372
rect 19705 19363 19763 19369
rect 19705 19360 19717 19363
rect 19392 19332 19717 19360
rect 19392 19320 19398 19332
rect 19705 19329 19717 19332
rect 19751 19329 19763 19363
rect 21174 19360 21180 19372
rect 21135 19332 21180 19360
rect 19705 19323 19763 19329
rect 21174 19320 21180 19332
rect 21232 19320 21238 19372
rect 1670 19292 1676 19304
rect 1631 19264 1676 19292
rect 1670 19252 1676 19264
rect 1728 19252 1734 19304
rect 1854 19292 1860 19304
rect 1815 19264 1860 19292
rect 1854 19252 1860 19264
rect 1912 19252 1918 19304
rect 2130 19292 2136 19304
rect 2091 19264 2136 19292
rect 2130 19252 2136 19264
rect 2188 19252 2194 19304
rect 12529 19295 12587 19301
rect 12529 19261 12541 19295
rect 12575 19261 12587 19295
rect 12529 19255 12587 19261
rect 12544 19156 12572 19255
rect 14274 19252 14280 19304
rect 14332 19292 14338 19304
rect 15197 19295 15255 19301
rect 15197 19292 15209 19295
rect 14332 19264 15209 19292
rect 14332 19252 14338 19264
rect 15197 19261 15209 19264
rect 15243 19261 15255 19295
rect 15197 19255 15255 19261
rect 15289 19295 15347 19301
rect 15289 19261 15301 19295
rect 15335 19261 15347 19295
rect 15289 19255 15347 19261
rect 19889 19295 19947 19301
rect 19889 19261 19901 19295
rect 19935 19292 19947 19295
rect 20254 19292 20260 19304
rect 19935 19264 20260 19292
rect 19935 19261 19947 19264
rect 19889 19255 19947 19261
rect 13998 19184 14004 19236
rect 14056 19224 14062 19236
rect 14734 19224 14740 19236
rect 14056 19196 14740 19224
rect 14056 19184 14062 19196
rect 14734 19184 14740 19196
rect 14792 19224 14798 19236
rect 15304 19224 15332 19255
rect 20254 19252 20260 19264
rect 20312 19252 20318 19304
rect 14792 19196 15332 19224
rect 14792 19184 14798 19196
rect 13909 19159 13967 19165
rect 13909 19156 13921 19159
rect 12544 19128 13921 19156
rect 13909 19125 13921 19128
rect 13955 19156 13967 19159
rect 14550 19156 14556 19168
rect 13955 19128 14556 19156
rect 13955 19125 13967 19128
rect 13909 19119 13967 19125
rect 14550 19116 14556 19128
rect 14608 19116 14614 19168
rect 17126 19116 17132 19168
rect 17184 19156 17190 19168
rect 18325 19159 18383 19165
rect 18325 19156 18337 19159
rect 17184 19128 18337 19156
rect 17184 19116 17190 19128
rect 18325 19125 18337 19128
rect 18371 19125 18383 19159
rect 18325 19119 18383 19125
rect 20993 19159 21051 19165
rect 20993 19125 21005 19159
rect 21039 19156 21051 19159
rect 21082 19156 21088 19168
rect 21039 19128 21088 19156
rect 21039 19125 21051 19128
rect 20993 19119 21051 19125
rect 21082 19116 21088 19128
rect 21140 19116 21146 19168
rect 27893 19159 27951 19165
rect 27893 19125 27905 19159
rect 27939 19156 27951 19159
rect 28350 19156 28356 19168
rect 27939 19128 28356 19156
rect 27939 19125 27951 19128
rect 27893 19119 27951 19125
rect 28350 19116 28356 19128
rect 28408 19116 28414 19168
rect 1104 19066 28888 19088
rect 1104 19014 4423 19066
rect 4475 19014 4487 19066
rect 4539 19014 4551 19066
rect 4603 19014 4615 19066
rect 4667 19014 4679 19066
rect 4731 19014 11369 19066
rect 11421 19014 11433 19066
rect 11485 19014 11497 19066
rect 11549 19014 11561 19066
rect 11613 19014 11625 19066
rect 11677 19014 18315 19066
rect 18367 19014 18379 19066
rect 18431 19014 18443 19066
rect 18495 19014 18507 19066
rect 18559 19014 18571 19066
rect 18623 19014 25261 19066
rect 25313 19014 25325 19066
rect 25377 19014 25389 19066
rect 25441 19014 25453 19066
rect 25505 19014 25517 19066
rect 25569 19014 28888 19066
rect 1104 18992 28888 19014
rect 1670 18912 1676 18964
rect 1728 18952 1734 18964
rect 1765 18955 1823 18961
rect 1765 18952 1777 18955
rect 1728 18924 1777 18952
rect 1728 18912 1734 18924
rect 1765 18921 1777 18924
rect 1811 18921 1823 18955
rect 1765 18915 1823 18921
rect 1854 18912 1860 18964
rect 1912 18952 1918 18964
rect 2501 18955 2559 18961
rect 2501 18952 2513 18955
rect 1912 18924 2513 18952
rect 1912 18912 1918 18924
rect 2501 18921 2513 18924
rect 2547 18921 2559 18955
rect 2501 18915 2559 18921
rect 12897 18955 12955 18961
rect 12897 18921 12909 18955
rect 12943 18952 12955 18955
rect 12986 18952 12992 18964
rect 12943 18924 12992 18952
rect 12943 18921 12955 18924
rect 12897 18915 12955 18921
rect 12986 18912 12992 18924
rect 13044 18952 13050 18964
rect 13814 18952 13820 18964
rect 13044 18924 13820 18952
rect 13044 18912 13050 18924
rect 13814 18912 13820 18924
rect 13872 18912 13878 18964
rect 16025 18955 16083 18961
rect 16025 18921 16037 18955
rect 16071 18921 16083 18955
rect 16025 18915 16083 18921
rect 16209 18955 16267 18961
rect 16209 18921 16221 18955
rect 16255 18952 16267 18955
rect 16574 18952 16580 18964
rect 16255 18924 16580 18952
rect 16255 18921 16267 18924
rect 16209 18915 16267 18921
rect 16040 18884 16068 18915
rect 16574 18912 16580 18924
rect 16632 18912 16638 18964
rect 17034 18952 17040 18964
rect 16684 18924 17040 18952
rect 16684 18884 16712 18924
rect 17034 18912 17040 18924
rect 17092 18912 17098 18964
rect 24854 18912 24860 18964
rect 24912 18952 24918 18964
rect 25041 18955 25099 18961
rect 25041 18952 25053 18955
rect 24912 18924 25053 18952
rect 24912 18912 24918 18924
rect 25041 18921 25053 18924
rect 25087 18921 25099 18955
rect 25041 18915 25099 18921
rect 16040 18856 16712 18884
rect 23201 18887 23259 18893
rect 23201 18853 23213 18887
rect 23247 18884 23259 18887
rect 24210 18884 24216 18896
rect 23247 18856 24216 18884
rect 23247 18853 23259 18856
rect 23201 18847 23259 18853
rect 24210 18844 24216 18856
rect 24268 18844 24274 18896
rect 14550 18816 14556 18828
rect 12728 18788 14556 18816
rect 2590 18748 2596 18760
rect 2551 18720 2596 18748
rect 2590 18708 2596 18720
rect 2648 18708 2654 18760
rect 12250 18708 12256 18760
rect 12308 18748 12314 18760
rect 12728 18757 12756 18788
rect 14550 18776 14556 18788
rect 14608 18776 14614 18828
rect 18046 18776 18052 18828
rect 18104 18816 18110 18828
rect 20809 18819 20867 18825
rect 20809 18816 20821 18819
rect 18104 18788 20821 18816
rect 18104 18776 18110 18788
rect 20809 18785 20821 18788
rect 20855 18785 20867 18819
rect 24670 18816 24676 18828
rect 24631 18788 24676 18816
rect 20809 18779 20867 18785
rect 24670 18776 24676 18788
rect 24728 18776 24734 18828
rect 26142 18776 26148 18828
rect 26200 18816 26206 18828
rect 26513 18819 26571 18825
rect 26513 18816 26525 18819
rect 26200 18788 26525 18816
rect 26200 18776 26206 18788
rect 26513 18785 26525 18788
rect 26559 18785 26571 18819
rect 28350 18816 28356 18828
rect 28311 18788 28356 18816
rect 26513 18779 26571 18785
rect 28350 18776 28356 18788
rect 28408 18776 28414 18828
rect 12713 18751 12771 18757
rect 12713 18748 12725 18751
rect 12308 18720 12725 18748
rect 12308 18708 12314 18720
rect 12713 18717 12725 18720
rect 12759 18717 12771 18751
rect 12713 18711 12771 18717
rect 12802 18708 12808 18760
rect 12860 18748 12866 18760
rect 12897 18751 12955 18757
rect 12897 18748 12909 18751
rect 12860 18720 12909 18748
rect 12860 18708 12866 18720
rect 12897 18717 12909 18720
rect 12943 18717 12955 18751
rect 12897 18711 12955 18717
rect 13357 18751 13415 18757
rect 13357 18717 13369 18751
rect 13403 18717 13415 18751
rect 13357 18711 13415 18717
rect 13541 18751 13599 18757
rect 13541 18717 13553 18751
rect 13587 18748 13599 18751
rect 13722 18748 13728 18760
rect 13587 18720 13728 18748
rect 13587 18717 13599 18720
rect 13541 18711 13599 18717
rect 13372 18680 13400 18711
rect 13722 18708 13728 18720
rect 13780 18708 13786 18760
rect 15654 18748 15660 18760
rect 15615 18720 15660 18748
rect 15654 18708 15660 18720
rect 15712 18708 15718 18760
rect 16669 18751 16727 18757
rect 16669 18717 16681 18751
rect 16715 18748 16727 18751
rect 16758 18748 16764 18760
rect 16715 18720 16764 18748
rect 16715 18717 16727 18720
rect 16669 18711 16727 18717
rect 16758 18708 16764 18720
rect 16816 18708 16822 18760
rect 16942 18757 16948 18760
rect 16936 18748 16948 18757
rect 16903 18720 16948 18748
rect 16936 18711 16948 18720
rect 16942 18708 16948 18711
rect 17000 18708 17006 18760
rect 18690 18748 18696 18760
rect 18651 18720 18696 18748
rect 18690 18708 18696 18720
rect 18748 18708 18754 18760
rect 19794 18748 19800 18760
rect 19755 18720 19800 18748
rect 19794 18708 19800 18720
rect 19852 18708 19858 18760
rect 21082 18757 21088 18760
rect 21076 18748 21088 18757
rect 21043 18720 21088 18748
rect 21076 18711 21088 18720
rect 21082 18708 21088 18711
rect 21140 18708 21146 18760
rect 22370 18708 22376 18760
rect 22428 18748 22434 18760
rect 22925 18751 22983 18757
rect 22925 18748 22937 18751
rect 22428 18720 22937 18748
rect 22428 18708 22434 18720
rect 22925 18717 22937 18720
rect 22971 18748 22983 18751
rect 23382 18748 23388 18760
rect 22971 18720 23388 18748
rect 22971 18717 22983 18720
rect 22925 18711 22983 18717
rect 23382 18708 23388 18720
rect 23440 18708 23446 18760
rect 23750 18708 23756 18760
rect 23808 18748 23814 18760
rect 24765 18751 24823 18757
rect 24765 18748 24777 18751
rect 23808 18720 24777 18748
rect 23808 18708 23814 18720
rect 24765 18717 24777 18720
rect 24811 18717 24823 18751
rect 24765 18711 24823 18717
rect 24854 18708 24860 18760
rect 24912 18748 24918 18760
rect 25869 18751 25927 18757
rect 25869 18748 25881 18751
rect 24912 18720 25881 18748
rect 24912 18708 24918 18720
rect 25869 18717 25881 18720
rect 25915 18717 25927 18751
rect 25869 18711 25927 18717
rect 13998 18680 14004 18692
rect 13372 18652 14004 18680
rect 13998 18640 14004 18652
rect 14056 18680 14062 18692
rect 14274 18680 14280 18692
rect 14056 18652 14280 18680
rect 14056 18640 14062 18652
rect 14274 18640 14280 18652
rect 14332 18640 14338 18692
rect 14461 18683 14519 18689
rect 14461 18649 14473 18683
rect 14507 18680 14519 18683
rect 14734 18680 14740 18692
rect 14507 18652 14740 18680
rect 14507 18649 14519 18652
rect 14461 18643 14519 18649
rect 14734 18640 14740 18652
rect 14792 18640 14798 18692
rect 15930 18640 15936 18692
rect 15988 18680 15994 18692
rect 19503 18683 19561 18689
rect 19503 18680 19515 18683
rect 15988 18652 19515 18680
rect 15988 18640 15994 18652
rect 19503 18649 19515 18652
rect 19549 18649 19561 18683
rect 19503 18643 19561 18649
rect 20073 18683 20131 18689
rect 20073 18649 20085 18683
rect 20119 18680 20131 18683
rect 20254 18680 20260 18692
rect 20119 18652 20260 18680
rect 20119 18649 20131 18652
rect 20073 18643 20131 18649
rect 20254 18640 20260 18652
rect 20312 18640 20318 18692
rect 20898 18640 20904 18692
rect 20956 18680 20962 18692
rect 23106 18680 23112 18692
rect 20956 18652 23112 18680
rect 20956 18640 20962 18652
rect 23106 18640 23112 18652
rect 23164 18640 23170 18692
rect 23201 18683 23259 18689
rect 23201 18649 23213 18683
rect 23247 18680 23259 18683
rect 23290 18680 23296 18692
rect 23247 18652 23296 18680
rect 23247 18649 23259 18652
rect 23201 18643 23259 18649
rect 23290 18640 23296 18652
rect 23348 18640 23354 18692
rect 27982 18640 27988 18692
rect 28040 18680 28046 18692
rect 28169 18683 28227 18689
rect 28169 18680 28181 18683
rect 28040 18652 28181 18680
rect 28040 18640 28046 18652
rect 28169 18649 28181 18652
rect 28215 18649 28227 18683
rect 28169 18643 28227 18649
rect 13446 18612 13452 18624
rect 13407 18584 13452 18612
rect 13446 18572 13452 18584
rect 13504 18572 13510 18624
rect 14642 18612 14648 18624
rect 14603 18584 14648 18612
rect 14642 18572 14648 18584
rect 14700 18572 14706 18624
rect 16025 18615 16083 18621
rect 16025 18581 16037 18615
rect 16071 18612 16083 18615
rect 17218 18612 17224 18624
rect 16071 18584 17224 18612
rect 16071 18581 16083 18584
rect 16025 18575 16083 18581
rect 17218 18572 17224 18584
rect 17276 18572 17282 18624
rect 17954 18572 17960 18624
rect 18012 18612 18018 18624
rect 18049 18615 18107 18621
rect 18049 18612 18061 18615
rect 18012 18584 18061 18612
rect 18012 18572 18018 18584
rect 18049 18581 18061 18584
rect 18095 18581 18107 18615
rect 18049 18575 18107 18581
rect 18230 18572 18236 18624
rect 18288 18612 18294 18624
rect 18509 18615 18567 18621
rect 18509 18612 18521 18615
rect 18288 18584 18521 18612
rect 18288 18572 18294 18584
rect 18509 18581 18521 18584
rect 18555 18581 18567 18615
rect 18509 18575 18567 18581
rect 19981 18615 20039 18621
rect 19981 18581 19993 18615
rect 20027 18612 20039 18615
rect 20806 18612 20812 18624
rect 20027 18584 20812 18612
rect 20027 18581 20039 18584
rect 19981 18575 20039 18581
rect 20806 18572 20812 18584
rect 20864 18572 20870 18624
rect 22186 18612 22192 18624
rect 22147 18584 22192 18612
rect 22186 18572 22192 18584
rect 22244 18572 22250 18624
rect 23014 18612 23020 18624
rect 22927 18584 23020 18612
rect 23014 18572 23020 18584
rect 23072 18612 23078 18624
rect 23566 18612 23572 18624
rect 23072 18584 23572 18612
rect 23072 18572 23078 18584
rect 23566 18572 23572 18584
rect 23624 18572 23630 18624
rect 25961 18615 26019 18621
rect 25961 18581 25973 18615
rect 26007 18612 26019 18615
rect 26694 18612 26700 18624
rect 26007 18584 26700 18612
rect 26007 18581 26019 18584
rect 25961 18575 26019 18581
rect 26694 18572 26700 18584
rect 26752 18572 26758 18624
rect 1104 18522 29048 18544
rect 1104 18470 7896 18522
rect 7948 18470 7960 18522
rect 8012 18470 8024 18522
rect 8076 18470 8088 18522
rect 8140 18470 8152 18522
rect 8204 18470 14842 18522
rect 14894 18470 14906 18522
rect 14958 18470 14970 18522
rect 15022 18470 15034 18522
rect 15086 18470 15098 18522
rect 15150 18470 21788 18522
rect 21840 18470 21852 18522
rect 21904 18470 21916 18522
rect 21968 18470 21980 18522
rect 22032 18470 22044 18522
rect 22096 18470 28734 18522
rect 28786 18470 28798 18522
rect 28850 18470 28862 18522
rect 28914 18470 28926 18522
rect 28978 18470 28990 18522
rect 29042 18470 29048 18522
rect 1104 18448 29048 18470
rect 16298 18408 16304 18420
rect 16259 18380 16304 18408
rect 16298 18368 16304 18380
rect 16356 18368 16362 18420
rect 17218 18408 17224 18420
rect 17179 18380 17224 18408
rect 17218 18368 17224 18380
rect 17276 18368 17282 18420
rect 21174 18368 21180 18420
rect 21232 18408 21238 18420
rect 21269 18411 21327 18417
rect 21269 18408 21281 18411
rect 21232 18380 21281 18408
rect 21232 18368 21238 18380
rect 21269 18377 21281 18380
rect 21315 18377 21327 18411
rect 21269 18371 21327 18377
rect 22186 18368 22192 18420
rect 22244 18408 22250 18420
rect 22373 18411 22431 18417
rect 22373 18408 22385 18411
rect 22244 18380 22385 18408
rect 22244 18368 22250 18380
rect 22373 18377 22385 18380
rect 22419 18377 22431 18411
rect 22373 18371 22431 18377
rect 22462 18368 22468 18420
rect 22520 18408 22526 18420
rect 22520 18380 22565 18408
rect 22520 18368 22526 18380
rect 23014 18368 23020 18420
rect 23072 18408 23078 18420
rect 23569 18411 23627 18417
rect 23569 18408 23581 18411
rect 23072 18380 23581 18408
rect 23072 18368 23078 18380
rect 23569 18377 23581 18380
rect 23615 18377 23627 18411
rect 23569 18371 23627 18377
rect 24670 18368 24676 18420
rect 24728 18408 24734 18420
rect 27341 18411 27399 18417
rect 27341 18408 27353 18411
rect 24728 18380 27353 18408
rect 24728 18368 24734 18380
rect 27341 18377 27353 18380
rect 27387 18377 27399 18411
rect 27982 18408 27988 18420
rect 27943 18380 27988 18408
rect 27341 18371 27399 18377
rect 27982 18368 27988 18380
rect 28040 18368 28046 18420
rect 13725 18343 13783 18349
rect 13725 18309 13737 18343
rect 13771 18340 13783 18343
rect 14458 18340 14464 18352
rect 13771 18312 14464 18340
rect 13771 18309 13783 18312
rect 13725 18303 13783 18309
rect 14458 18300 14464 18312
rect 14516 18340 14522 18352
rect 16114 18340 16120 18352
rect 14516 18312 14872 18340
rect 16075 18312 16120 18340
rect 14516 18300 14522 18312
rect 1578 18272 1584 18284
rect 1539 18244 1584 18272
rect 1578 18232 1584 18244
rect 1636 18232 1642 18284
rect 12250 18272 12256 18284
rect 12211 18244 12256 18272
rect 12250 18232 12256 18244
rect 12308 18232 12314 18284
rect 12805 18275 12863 18281
rect 12805 18241 12817 18275
rect 12851 18241 12863 18275
rect 12805 18235 12863 18241
rect 11882 18164 11888 18216
rect 11940 18204 11946 18216
rect 12437 18207 12495 18213
rect 12437 18204 12449 18207
rect 11940 18176 12449 18204
rect 11940 18164 11946 18176
rect 12437 18173 12449 18176
rect 12483 18173 12495 18207
rect 12820 18204 12848 18235
rect 12894 18232 12900 18284
rect 12952 18272 12958 18284
rect 13446 18272 13452 18284
rect 12952 18244 12997 18272
rect 13280 18244 13452 18272
rect 12952 18232 12958 18244
rect 13280 18204 13308 18244
rect 13446 18232 13452 18244
rect 13504 18272 13510 18284
rect 13587 18275 13645 18281
rect 13587 18272 13599 18275
rect 13504 18244 13599 18272
rect 13504 18232 13510 18244
rect 13587 18241 13599 18244
rect 13633 18241 13645 18275
rect 13814 18272 13820 18284
rect 13775 18244 13820 18272
rect 13587 18235 13645 18241
rect 13814 18232 13820 18244
rect 13872 18232 13878 18284
rect 13998 18272 14004 18284
rect 13959 18244 14004 18272
rect 13998 18232 14004 18244
rect 14056 18232 14062 18284
rect 14090 18232 14096 18284
rect 14148 18272 14154 18284
rect 14550 18272 14556 18284
rect 14148 18244 14193 18272
rect 14511 18244 14556 18272
rect 14148 18232 14154 18244
rect 14550 18232 14556 18244
rect 14608 18232 14614 18284
rect 14734 18272 14740 18284
rect 14695 18244 14740 18272
rect 14734 18232 14740 18244
rect 14792 18232 14798 18284
rect 14844 18281 14872 18312
rect 16114 18300 16120 18312
rect 16172 18300 16178 18352
rect 16758 18300 16764 18352
rect 16816 18340 16822 18352
rect 18046 18340 18052 18352
rect 16816 18312 18052 18340
rect 16816 18300 16822 18312
rect 18046 18300 18052 18312
rect 18104 18340 18110 18352
rect 18233 18343 18291 18349
rect 18233 18340 18245 18343
rect 18104 18312 18245 18340
rect 18104 18300 18110 18312
rect 18233 18309 18245 18312
rect 18279 18309 18291 18343
rect 18233 18303 18291 18309
rect 19981 18343 20039 18349
rect 19981 18309 19993 18343
rect 20027 18340 20039 18343
rect 22554 18340 22560 18352
rect 20027 18312 22560 18340
rect 20027 18309 20039 18312
rect 19981 18303 20039 18309
rect 22554 18300 22560 18312
rect 22612 18300 22618 18352
rect 23106 18300 23112 18352
rect 23164 18340 23170 18352
rect 24397 18343 24455 18349
rect 24397 18340 24409 18343
rect 23164 18312 24409 18340
rect 23164 18300 23170 18312
rect 24397 18309 24409 18312
rect 24443 18309 24455 18343
rect 24397 18303 24455 18309
rect 25400 18343 25458 18349
rect 25400 18309 25412 18343
rect 25446 18340 25458 18343
rect 25682 18340 25688 18352
rect 25446 18312 25688 18340
rect 25446 18309 25458 18312
rect 25400 18303 25458 18309
rect 25682 18300 25688 18312
rect 25740 18300 25746 18352
rect 14829 18275 14887 18281
rect 14829 18241 14841 18275
rect 14875 18241 14887 18275
rect 15746 18272 15752 18284
rect 15659 18244 15752 18272
rect 14829 18235 14887 18241
rect 15746 18232 15752 18244
rect 15804 18272 15810 18284
rect 16853 18275 16911 18281
rect 16853 18272 16865 18275
rect 15804 18244 16865 18272
rect 15804 18232 15810 18244
rect 16853 18241 16865 18244
rect 16899 18241 16911 18275
rect 17034 18272 17040 18284
rect 16995 18244 17040 18272
rect 16853 18235 16911 18241
rect 17034 18232 17040 18244
rect 17092 18232 17098 18284
rect 21085 18275 21143 18281
rect 21085 18241 21097 18275
rect 21131 18272 21143 18275
rect 23385 18275 23443 18281
rect 23385 18272 23397 18275
rect 21131 18244 22048 18272
rect 21131 18241 21143 18244
rect 21085 18235 21143 18241
rect 20898 18204 20904 18216
rect 12820 18176 13308 18204
rect 20859 18176 20904 18204
rect 12437 18167 12495 18173
rect 20898 18164 20904 18176
rect 20956 18164 20962 18216
rect 1765 18139 1823 18145
rect 1765 18105 1777 18139
rect 1811 18136 1823 18139
rect 15194 18136 15200 18148
rect 1811 18108 15200 18136
rect 1811 18105 1823 18108
rect 1765 18099 1823 18105
rect 15194 18096 15200 18108
rect 15252 18096 15258 18148
rect 22020 18145 22048 18244
rect 23216 18244 23397 18272
rect 22557 18207 22615 18213
rect 22557 18173 22569 18207
rect 22603 18173 22615 18207
rect 22557 18167 22615 18173
rect 22005 18139 22063 18145
rect 22005 18105 22017 18139
rect 22051 18105 22063 18139
rect 22005 18099 22063 18105
rect 13446 18068 13452 18080
rect 13407 18040 13452 18068
rect 13446 18028 13452 18040
rect 13504 18028 13510 18080
rect 14550 18068 14556 18080
rect 14511 18040 14556 18068
rect 14550 18028 14556 18040
rect 14608 18028 14614 18080
rect 16117 18071 16175 18077
rect 16117 18037 16129 18071
rect 16163 18068 16175 18071
rect 16850 18068 16856 18080
rect 16163 18040 16856 18068
rect 16163 18037 16175 18040
rect 16117 18031 16175 18037
rect 16850 18028 16856 18040
rect 16908 18068 16914 18080
rect 17402 18068 17408 18080
rect 16908 18040 17408 18068
rect 16908 18028 16914 18040
rect 17402 18028 17408 18040
rect 17460 18028 17466 18080
rect 19978 18028 19984 18080
rect 20036 18068 20042 18080
rect 22572 18068 22600 18167
rect 23216 18136 23244 18244
rect 23385 18241 23397 18244
rect 23431 18241 23443 18275
rect 23385 18235 23443 18241
rect 23661 18275 23719 18281
rect 23661 18241 23673 18275
rect 23707 18241 23719 18275
rect 23661 18235 23719 18241
rect 24121 18275 24179 18281
rect 24121 18241 24133 18275
rect 24167 18241 24179 18275
rect 24121 18235 24179 18241
rect 23290 18164 23296 18216
rect 23348 18204 23354 18216
rect 23676 18204 23704 18235
rect 23348 18176 23704 18204
rect 24136 18204 24164 18235
rect 24210 18232 24216 18284
rect 24268 18272 24274 18284
rect 24268 18244 24313 18272
rect 24268 18232 24274 18244
rect 25038 18232 25044 18284
rect 25096 18272 25102 18284
rect 25133 18275 25191 18281
rect 25133 18272 25145 18275
rect 25096 18244 25145 18272
rect 25096 18232 25102 18244
rect 25133 18241 25145 18244
rect 25179 18241 25191 18275
rect 27157 18275 27215 18281
rect 27157 18272 27169 18275
rect 25133 18235 25191 18241
rect 26528 18244 27169 18272
rect 24578 18204 24584 18216
rect 24136 18176 24584 18204
rect 23348 18164 23354 18176
rect 24578 18164 24584 18176
rect 24636 18164 24642 18216
rect 23934 18136 23940 18148
rect 23216 18108 23940 18136
rect 23934 18096 23940 18108
rect 23992 18096 23998 18148
rect 26528 18145 26556 18244
rect 27157 18241 27169 18244
rect 27203 18241 27215 18275
rect 27157 18235 27215 18241
rect 27614 18232 27620 18284
rect 27672 18272 27678 18284
rect 27893 18275 27951 18281
rect 27893 18272 27905 18275
rect 27672 18244 27905 18272
rect 27672 18232 27678 18244
rect 27893 18241 27905 18244
rect 27939 18241 27951 18275
rect 27893 18235 27951 18241
rect 26513 18139 26571 18145
rect 26513 18105 26525 18139
rect 26559 18105 26571 18139
rect 26513 18099 26571 18105
rect 23198 18068 23204 18080
rect 20036 18040 22600 18068
rect 23159 18040 23204 18068
rect 20036 18028 20042 18040
rect 23198 18028 23204 18040
rect 23256 18028 23262 18080
rect 24305 18071 24363 18077
rect 24305 18037 24317 18071
rect 24351 18068 24363 18071
rect 24394 18068 24400 18080
rect 24351 18040 24400 18068
rect 24351 18037 24363 18040
rect 24305 18031 24363 18037
rect 24394 18028 24400 18040
rect 24452 18028 24458 18080
rect 1104 17978 28888 18000
rect 1104 17926 4423 17978
rect 4475 17926 4487 17978
rect 4539 17926 4551 17978
rect 4603 17926 4615 17978
rect 4667 17926 4679 17978
rect 4731 17926 11369 17978
rect 11421 17926 11433 17978
rect 11485 17926 11497 17978
rect 11549 17926 11561 17978
rect 11613 17926 11625 17978
rect 11677 17926 18315 17978
rect 18367 17926 18379 17978
rect 18431 17926 18443 17978
rect 18495 17926 18507 17978
rect 18559 17926 18571 17978
rect 18623 17926 25261 17978
rect 25313 17926 25325 17978
rect 25377 17926 25389 17978
rect 25441 17926 25453 17978
rect 25505 17926 25517 17978
rect 25569 17926 28888 17978
rect 1104 17904 28888 17926
rect 13556 17836 14780 17864
rect 2774 17728 2780 17740
rect 2735 17700 2780 17728
rect 2774 17688 2780 17700
rect 2832 17688 2838 17740
rect 1578 17660 1584 17672
rect 1539 17632 1584 17660
rect 1578 17620 1584 17632
rect 1636 17620 1642 17672
rect 13556 17669 13584 17836
rect 14752 17808 14780 17836
rect 16114 17824 16120 17876
rect 16172 17864 16178 17876
rect 16301 17867 16359 17873
rect 16301 17864 16313 17867
rect 16172 17836 16313 17864
rect 16172 17824 16178 17836
rect 16301 17833 16313 17836
rect 16347 17833 16359 17867
rect 16301 17827 16359 17833
rect 18509 17867 18567 17873
rect 18509 17833 18521 17867
rect 18555 17864 18567 17867
rect 18690 17864 18696 17876
rect 18555 17836 18696 17864
rect 18555 17833 18567 17836
rect 18509 17827 18567 17833
rect 18690 17824 18696 17836
rect 18748 17824 18754 17876
rect 21269 17867 21327 17873
rect 21269 17833 21281 17867
rect 21315 17864 21327 17867
rect 21634 17864 21640 17876
rect 21315 17836 21640 17864
rect 21315 17833 21327 17836
rect 21269 17827 21327 17833
rect 21634 17824 21640 17836
rect 21692 17824 21698 17876
rect 23106 17824 23112 17876
rect 23164 17864 23170 17876
rect 23842 17864 23848 17876
rect 23164 17836 23848 17864
rect 23164 17824 23170 17836
rect 23842 17824 23848 17836
rect 23900 17824 23906 17876
rect 24026 17824 24032 17876
rect 24084 17864 24090 17876
rect 24765 17867 24823 17873
rect 24765 17864 24777 17867
rect 24084 17836 24777 17864
rect 24084 17824 24090 17836
rect 24765 17833 24777 17836
rect 24811 17833 24823 17867
rect 24765 17827 24823 17833
rect 14642 17796 14648 17808
rect 14568 17768 14648 17796
rect 14568 17737 14596 17768
rect 14642 17756 14648 17768
rect 14700 17756 14706 17808
rect 14734 17756 14740 17808
rect 14792 17796 14798 17808
rect 19613 17799 19671 17805
rect 19613 17796 19625 17799
rect 14792 17768 19625 17796
rect 14792 17756 14798 17768
rect 19613 17765 19625 17768
rect 19659 17765 19671 17799
rect 19613 17759 19671 17765
rect 19720 17768 23520 17796
rect 13633 17731 13691 17737
rect 13633 17697 13645 17731
rect 13679 17728 13691 17731
rect 14461 17731 14519 17737
rect 14461 17728 14473 17731
rect 13679 17700 14473 17728
rect 13679 17697 13691 17700
rect 13633 17691 13691 17697
rect 14461 17697 14473 17700
rect 14507 17697 14519 17731
rect 14461 17691 14519 17697
rect 14553 17731 14611 17737
rect 14553 17697 14565 17731
rect 14599 17697 14611 17731
rect 14553 17691 14611 17697
rect 16206 17688 16212 17740
rect 16264 17728 16270 17740
rect 19720 17728 19748 17768
rect 16264 17700 19748 17728
rect 20073 17731 20131 17737
rect 16264 17688 16270 17700
rect 20073 17697 20085 17731
rect 20119 17728 20131 17731
rect 20162 17728 20168 17740
rect 20119 17700 20168 17728
rect 20119 17697 20131 17700
rect 20073 17691 20131 17697
rect 20162 17688 20168 17700
rect 20220 17688 20226 17740
rect 23198 17728 23204 17740
rect 23159 17700 23204 17728
rect 23198 17688 23204 17700
rect 23256 17688 23262 17740
rect 23382 17728 23388 17740
rect 23343 17700 23388 17728
rect 23382 17688 23388 17700
rect 23440 17688 23446 17740
rect 13541 17663 13599 17669
rect 13541 17629 13553 17663
rect 13587 17629 13599 17663
rect 13722 17660 13728 17672
rect 13683 17632 13728 17660
rect 13541 17623 13599 17629
rect 13722 17620 13728 17632
rect 13780 17620 13786 17672
rect 13814 17620 13820 17672
rect 13872 17660 13878 17672
rect 14645 17663 14703 17669
rect 14645 17660 14657 17663
rect 13872 17632 14657 17660
rect 13872 17620 13878 17632
rect 14645 17629 14657 17632
rect 14691 17629 14703 17663
rect 14645 17623 14703 17629
rect 14734 17620 14740 17672
rect 14792 17660 14798 17672
rect 14792 17632 14837 17660
rect 14792 17620 14798 17632
rect 15838 17620 15844 17672
rect 15896 17660 15902 17672
rect 15933 17663 15991 17669
rect 15933 17660 15945 17663
rect 15896 17632 15945 17660
rect 15896 17620 15902 17632
rect 15933 17629 15945 17632
rect 15979 17629 15991 17663
rect 15933 17623 15991 17629
rect 18693 17663 18751 17669
rect 18693 17629 18705 17663
rect 18739 17629 18751 17663
rect 18693 17623 18751 17629
rect 1765 17595 1823 17601
rect 1765 17561 1777 17595
rect 1811 17592 1823 17595
rect 2406 17592 2412 17604
rect 1811 17564 2412 17592
rect 1811 17561 1823 17564
rect 1765 17555 1823 17561
rect 2406 17552 2412 17564
rect 2464 17552 2470 17604
rect 16117 17595 16175 17601
rect 12406 17564 14320 17592
rect 7742 17484 7748 17536
rect 7800 17524 7806 17536
rect 12406 17524 12434 17564
rect 14292 17533 14320 17564
rect 16117 17561 16129 17595
rect 16163 17592 16175 17595
rect 16574 17592 16580 17604
rect 16163 17564 16580 17592
rect 16163 17561 16175 17564
rect 16117 17555 16175 17561
rect 16574 17552 16580 17564
rect 16632 17552 16638 17604
rect 18708 17592 18736 17623
rect 18782 17620 18788 17672
rect 18840 17660 18846 17672
rect 19886 17660 19892 17672
rect 18840 17632 19892 17660
rect 18840 17620 18846 17632
rect 19886 17620 19892 17632
rect 19944 17660 19950 17672
rect 20898 17660 20904 17672
rect 19944 17632 20904 17660
rect 19944 17620 19950 17632
rect 20898 17620 20904 17632
rect 20956 17620 20962 17672
rect 22554 17660 22560 17672
rect 22515 17632 22560 17660
rect 22554 17620 22560 17632
rect 22612 17620 22618 17672
rect 23106 17620 23112 17672
rect 23164 17660 23170 17672
rect 23492 17669 23520 17768
rect 23860 17728 23888 17824
rect 27890 17796 27896 17808
rect 26528 17768 27896 17796
rect 26528 17737 26556 17768
rect 27890 17756 27896 17768
rect 27948 17756 27954 17808
rect 26513 17731 26571 17737
rect 23860 17700 24808 17728
rect 23293 17663 23351 17669
rect 23293 17660 23305 17663
rect 23164 17632 23305 17660
rect 23164 17620 23170 17632
rect 23293 17629 23305 17632
rect 23339 17629 23351 17663
rect 23293 17623 23351 17629
rect 23477 17663 23535 17669
rect 23477 17629 23489 17663
rect 23523 17660 23535 17663
rect 23842 17660 23848 17672
rect 23523 17632 23848 17660
rect 23523 17629 23535 17632
rect 23477 17623 23535 17629
rect 23842 17620 23848 17632
rect 23900 17620 23906 17672
rect 19794 17592 19800 17604
rect 18708 17564 19800 17592
rect 19794 17552 19800 17564
rect 19852 17552 19858 17604
rect 20165 17595 20223 17601
rect 20165 17561 20177 17595
rect 20211 17561 20223 17595
rect 20165 17555 20223 17561
rect 7800 17496 12434 17524
rect 14277 17527 14335 17533
rect 7800 17484 7806 17496
rect 14277 17493 14289 17527
rect 14323 17493 14335 17527
rect 20070 17524 20076 17536
rect 20031 17496 20076 17524
rect 14277 17487 14335 17493
rect 20070 17484 20076 17496
rect 20128 17484 20134 17536
rect 20180 17524 20208 17555
rect 23382 17552 23388 17604
rect 23440 17592 23446 17604
rect 24780 17601 24808 17700
rect 26513 17697 26525 17731
rect 26559 17697 26571 17731
rect 26694 17728 26700 17740
rect 26655 17700 26700 17728
rect 26513 17691 26571 17697
rect 26694 17688 26700 17700
rect 26752 17688 26758 17740
rect 28353 17731 28411 17737
rect 28353 17697 28365 17731
rect 28399 17728 28411 17731
rect 28626 17728 28632 17740
rect 28399 17700 28632 17728
rect 28399 17697 28411 17700
rect 28353 17691 28411 17697
rect 28626 17688 28632 17700
rect 28684 17688 28690 17740
rect 24749 17595 24808 17601
rect 23440 17564 24716 17592
rect 23440 17552 23446 17564
rect 20254 17524 20260 17536
rect 20180 17496 20260 17524
rect 20254 17484 20260 17496
rect 20312 17524 20318 17536
rect 22646 17524 22652 17536
rect 20312 17496 22652 17524
rect 20312 17484 20318 17496
rect 22646 17484 22652 17496
rect 22704 17484 22710 17536
rect 23017 17527 23075 17533
rect 23017 17493 23029 17527
rect 23063 17524 23075 17527
rect 23474 17524 23480 17536
rect 23063 17496 23480 17524
rect 23063 17493 23075 17496
rect 23017 17487 23075 17493
rect 23474 17484 23480 17496
rect 23532 17484 23538 17536
rect 24578 17524 24584 17536
rect 24539 17496 24584 17524
rect 24578 17484 24584 17496
rect 24636 17484 24642 17536
rect 24688 17524 24716 17564
rect 24749 17561 24761 17595
rect 24795 17564 24808 17595
rect 24949 17595 25007 17601
rect 24795 17561 24807 17564
rect 24749 17555 24807 17561
rect 24949 17561 24961 17595
rect 24995 17561 25007 17595
rect 24949 17555 25007 17561
rect 24964 17524 24992 17555
rect 25498 17524 25504 17536
rect 24688 17496 25504 17524
rect 25498 17484 25504 17496
rect 25556 17484 25562 17536
rect 1104 17434 29048 17456
rect 1104 17382 7896 17434
rect 7948 17382 7960 17434
rect 8012 17382 8024 17434
rect 8076 17382 8088 17434
rect 8140 17382 8152 17434
rect 8204 17382 14842 17434
rect 14894 17382 14906 17434
rect 14958 17382 14970 17434
rect 15022 17382 15034 17434
rect 15086 17382 15098 17434
rect 15150 17382 21788 17434
rect 21840 17382 21852 17434
rect 21904 17382 21916 17434
rect 21968 17382 21980 17434
rect 22032 17382 22044 17434
rect 22096 17382 28734 17434
rect 28786 17382 28798 17434
rect 28850 17382 28862 17434
rect 28914 17382 28926 17434
rect 28978 17382 28990 17434
rect 29042 17382 29048 17434
rect 1104 17360 29048 17382
rect 2406 17320 2412 17332
rect 2367 17292 2412 17320
rect 2406 17280 2412 17292
rect 2464 17280 2470 17332
rect 15746 17320 15752 17332
rect 15707 17292 15752 17320
rect 15746 17280 15752 17292
rect 15804 17280 15810 17332
rect 19429 17323 19487 17329
rect 19429 17289 19441 17323
rect 19475 17320 19487 17323
rect 20070 17320 20076 17332
rect 19475 17292 20076 17320
rect 19475 17289 19487 17292
rect 19429 17283 19487 17289
rect 20070 17280 20076 17292
rect 20128 17320 20134 17332
rect 20257 17323 20315 17329
rect 20257 17320 20269 17323
rect 20128 17292 20269 17320
rect 20128 17280 20134 17292
rect 20257 17289 20269 17292
rect 20303 17289 20315 17323
rect 20257 17283 20315 17289
rect 20349 17323 20407 17329
rect 20349 17289 20361 17323
rect 20395 17320 20407 17323
rect 23014 17320 23020 17332
rect 20395 17292 23020 17320
rect 20395 17289 20407 17292
rect 20349 17283 20407 17289
rect 23014 17280 23020 17292
rect 23072 17280 23078 17332
rect 24118 17320 24124 17332
rect 23124 17292 24124 17320
rect 13998 17212 14004 17264
rect 14056 17252 14062 17264
rect 18322 17261 18328 17264
rect 14056 17224 18184 17252
rect 14056 17212 14062 17224
rect 1578 17144 1584 17196
rect 1636 17184 1642 17196
rect 1673 17187 1731 17193
rect 1673 17184 1685 17187
rect 1636 17156 1685 17184
rect 1636 17144 1642 17156
rect 1673 17153 1685 17156
rect 1719 17153 1731 17187
rect 2498 17184 2504 17196
rect 2459 17156 2504 17184
rect 1673 17147 1731 17153
rect 2498 17144 2504 17156
rect 2556 17184 2562 17196
rect 4338 17184 4344 17196
rect 2556 17156 4344 17184
rect 2556 17144 2562 17156
rect 4338 17144 4344 17156
rect 4396 17144 4402 17196
rect 14384 17193 14412 17224
rect 14369 17187 14427 17193
rect 14369 17153 14381 17187
rect 14415 17153 14427 17187
rect 14550 17184 14556 17196
rect 14511 17156 14556 17184
rect 14369 17147 14427 17153
rect 14550 17144 14556 17156
rect 14608 17144 14614 17196
rect 15838 17144 15844 17196
rect 15896 17184 15902 17196
rect 15933 17187 15991 17193
rect 15933 17184 15945 17187
rect 15896 17156 15945 17184
rect 15896 17144 15902 17156
rect 15933 17153 15945 17156
rect 15979 17153 15991 17187
rect 18046 17184 18052 17196
rect 18007 17156 18052 17184
rect 15933 17147 15991 17153
rect 18046 17144 18052 17156
rect 18104 17144 18110 17196
rect 18156 17184 18184 17224
rect 18316 17215 18328 17261
rect 18380 17252 18386 17264
rect 22079 17255 22137 17261
rect 22079 17252 22091 17255
rect 18380 17224 18416 17252
rect 18524 17224 22091 17252
rect 18322 17212 18328 17215
rect 18380 17212 18386 17224
rect 18524 17184 18552 17224
rect 22079 17221 22091 17224
rect 22125 17221 22137 17255
rect 22079 17215 22137 17221
rect 22186 17212 22192 17264
rect 22244 17252 22250 17264
rect 22373 17255 22431 17261
rect 22373 17252 22385 17255
rect 22244 17224 22385 17252
rect 22244 17212 22250 17224
rect 22373 17221 22385 17224
rect 22419 17221 22431 17255
rect 22554 17252 22560 17264
rect 22515 17224 22560 17252
rect 22373 17215 22431 17221
rect 22554 17212 22560 17224
rect 22612 17212 22618 17264
rect 22646 17212 22652 17264
rect 22704 17252 22710 17264
rect 23124 17252 23152 17292
rect 24118 17280 24124 17292
rect 24176 17280 24182 17332
rect 25498 17320 25504 17332
rect 25459 17292 25504 17320
rect 25498 17280 25504 17292
rect 25556 17280 25562 17332
rect 25038 17252 25044 17264
rect 22704 17224 23152 17252
rect 24136 17224 25044 17252
rect 22704 17212 22710 17224
rect 18156 17156 18552 17184
rect 21634 17144 21640 17196
rect 21692 17184 21698 17196
rect 24136 17193 24164 17224
rect 25038 17212 25044 17224
rect 25096 17212 25102 17264
rect 24394 17193 24400 17196
rect 24121 17187 24179 17193
rect 24121 17184 24133 17187
rect 21692 17156 24133 17184
rect 21692 17144 21698 17156
rect 24121 17153 24133 17156
rect 24167 17153 24179 17187
rect 24388 17184 24400 17193
rect 24355 17156 24400 17184
rect 24121 17147 24179 17153
rect 24388 17147 24400 17156
rect 24394 17144 24400 17147
rect 24452 17144 24458 17196
rect 26234 17184 26240 17196
rect 26195 17156 26240 17184
rect 26234 17144 26240 17156
rect 26292 17144 26298 17196
rect 27433 17187 27491 17193
rect 27433 17153 27445 17187
rect 27479 17184 27491 17187
rect 28258 17184 28264 17196
rect 27479 17156 28264 17184
rect 27479 17153 27491 17156
rect 27433 17147 27491 17153
rect 16117 17119 16175 17125
rect 16117 17085 16129 17119
rect 16163 17116 16175 17119
rect 16574 17116 16580 17128
rect 16163 17088 16580 17116
rect 16163 17085 16175 17088
rect 16117 17079 16175 17085
rect 16574 17076 16580 17088
rect 16632 17076 16638 17128
rect 19978 17076 19984 17128
rect 20036 17116 20042 17128
rect 20438 17116 20444 17128
rect 20036 17088 20444 17116
rect 20036 17076 20042 17088
rect 20438 17076 20444 17088
rect 20496 17076 20502 17128
rect 14550 17048 14556 17060
rect 14511 17020 14556 17048
rect 14550 17008 14556 17020
rect 14608 17048 14614 17060
rect 14734 17048 14740 17060
rect 14608 17020 14740 17048
rect 14608 17008 14614 17020
rect 14734 17008 14740 17020
rect 14792 17008 14798 17060
rect 19794 17008 19800 17060
rect 19852 17048 19858 17060
rect 19889 17051 19947 17057
rect 19889 17048 19901 17051
rect 19852 17020 19901 17048
rect 19852 17008 19858 17020
rect 19889 17017 19901 17020
rect 19935 17017 19947 17051
rect 27448 17048 27476 17147
rect 28258 17144 28264 17156
rect 28316 17144 28322 17196
rect 19889 17011 19947 17017
rect 25792 17020 27476 17048
rect 20530 16940 20536 16992
rect 20588 16980 20594 16992
rect 25792 16980 25820 17020
rect 20588 16952 25820 16980
rect 20588 16940 20594 16952
rect 25866 16940 25872 16992
rect 25924 16980 25930 16992
rect 26145 16983 26203 16989
rect 26145 16980 26157 16983
rect 25924 16952 26157 16980
rect 25924 16940 25930 16952
rect 26145 16949 26157 16952
rect 26191 16949 26203 16983
rect 26145 16943 26203 16949
rect 26694 16940 26700 16992
rect 26752 16980 26758 16992
rect 27341 16983 27399 16989
rect 27341 16980 27353 16983
rect 26752 16952 27353 16980
rect 26752 16940 26758 16952
rect 27341 16949 27353 16952
rect 27387 16949 27399 16983
rect 27890 16980 27896 16992
rect 27851 16952 27896 16980
rect 27341 16943 27399 16949
rect 27890 16940 27896 16952
rect 27948 16940 27954 16992
rect 1104 16890 28888 16912
rect 1104 16838 4423 16890
rect 4475 16838 4487 16890
rect 4539 16838 4551 16890
rect 4603 16838 4615 16890
rect 4667 16838 4679 16890
rect 4731 16838 11369 16890
rect 11421 16838 11433 16890
rect 11485 16838 11497 16890
rect 11549 16838 11561 16890
rect 11613 16838 11625 16890
rect 11677 16838 18315 16890
rect 18367 16838 18379 16890
rect 18431 16838 18443 16890
rect 18495 16838 18507 16890
rect 18559 16838 18571 16890
rect 18623 16838 25261 16890
rect 25313 16838 25325 16890
rect 25377 16838 25389 16890
rect 25441 16838 25453 16890
rect 25505 16838 25517 16890
rect 25569 16838 28888 16890
rect 1104 16816 28888 16838
rect 15654 16736 15660 16788
rect 15712 16776 15718 16788
rect 15933 16779 15991 16785
rect 15933 16776 15945 16779
rect 15712 16748 15945 16776
rect 15712 16736 15718 16748
rect 15933 16745 15945 16748
rect 15979 16745 15991 16779
rect 15933 16739 15991 16745
rect 16117 16779 16175 16785
rect 16117 16745 16129 16779
rect 16163 16776 16175 16779
rect 16574 16776 16580 16788
rect 16163 16748 16580 16776
rect 16163 16745 16175 16748
rect 16117 16739 16175 16745
rect 16574 16736 16580 16748
rect 16632 16776 16638 16788
rect 17678 16776 17684 16788
rect 16632 16748 17684 16776
rect 16632 16736 16638 16748
rect 17678 16736 17684 16748
rect 17736 16776 17742 16788
rect 17954 16776 17960 16788
rect 17736 16748 17960 16776
rect 17736 16736 17742 16748
rect 17954 16736 17960 16748
rect 18012 16736 18018 16788
rect 24946 16708 24952 16720
rect 22066 16680 24952 16708
rect 1670 16532 1676 16584
rect 1728 16572 1734 16584
rect 1765 16575 1823 16581
rect 1765 16572 1777 16575
rect 1728 16544 1777 16572
rect 1728 16532 1734 16544
rect 1765 16541 1777 16544
rect 1811 16541 1823 16575
rect 1765 16535 1823 16541
rect 19242 16532 19248 16584
rect 19300 16572 19306 16584
rect 20625 16575 20683 16581
rect 20625 16572 20637 16575
rect 19300 16544 20637 16572
rect 19300 16532 19306 16544
rect 20625 16541 20637 16544
rect 20671 16541 20683 16575
rect 20625 16535 20683 16541
rect 21450 16532 21456 16584
rect 21508 16572 21514 16584
rect 22066 16572 22094 16680
rect 24946 16668 24952 16680
rect 25004 16668 25010 16720
rect 27890 16708 27896 16720
rect 26528 16680 27896 16708
rect 23842 16600 23848 16652
rect 23900 16640 23906 16652
rect 26528 16649 26556 16680
rect 27890 16668 27896 16680
rect 27948 16668 27954 16720
rect 25685 16643 25743 16649
rect 25685 16640 25697 16643
rect 23900 16612 25697 16640
rect 23900 16600 23906 16612
rect 25685 16609 25697 16612
rect 25731 16609 25743 16643
rect 25685 16603 25743 16609
rect 26513 16643 26571 16649
rect 26513 16609 26525 16643
rect 26559 16609 26571 16643
rect 26694 16640 26700 16652
rect 26655 16612 26700 16640
rect 26513 16603 26571 16609
rect 26694 16600 26700 16612
rect 26752 16600 26758 16652
rect 23014 16572 23020 16584
rect 21508 16544 22094 16572
rect 22975 16544 23020 16572
rect 21508 16532 21514 16544
rect 23014 16532 23020 16544
rect 23072 16532 23078 16584
rect 23201 16575 23259 16581
rect 23201 16541 23213 16575
rect 23247 16541 23259 16575
rect 23474 16572 23480 16584
rect 23435 16544 23480 16572
rect 23201 16535 23259 16541
rect 15838 16464 15844 16516
rect 15896 16504 15902 16516
rect 16085 16507 16143 16513
rect 16085 16504 16097 16507
rect 15896 16476 16097 16504
rect 15896 16464 15902 16476
rect 16085 16473 16097 16476
rect 16131 16473 16143 16507
rect 16085 16467 16143 16473
rect 16301 16507 16359 16513
rect 16301 16473 16313 16507
rect 16347 16504 16359 16507
rect 17034 16504 17040 16516
rect 16347 16476 17040 16504
rect 16347 16473 16359 16476
rect 16301 16467 16359 16473
rect 17034 16464 17040 16476
rect 17092 16504 17098 16516
rect 18874 16504 18880 16516
rect 17092 16476 18880 16504
rect 17092 16464 17098 16476
rect 18874 16464 18880 16476
rect 18932 16464 18938 16516
rect 20714 16464 20720 16516
rect 20772 16504 20778 16516
rect 20870 16507 20928 16513
rect 20870 16504 20882 16507
rect 20772 16476 20882 16504
rect 20772 16464 20778 16476
rect 20870 16473 20882 16476
rect 20916 16473 20928 16507
rect 23216 16504 23244 16535
rect 23474 16532 23480 16544
rect 23532 16532 23538 16584
rect 24578 16504 24584 16516
rect 23216 16476 24584 16504
rect 20870 16467 20928 16473
rect 24578 16464 24584 16476
rect 24636 16464 24642 16516
rect 24765 16507 24823 16513
rect 24765 16473 24777 16507
rect 24811 16504 24823 16507
rect 25866 16504 25872 16516
rect 24811 16476 25872 16504
rect 24811 16473 24823 16476
rect 24765 16467 24823 16473
rect 25866 16464 25872 16476
rect 25924 16464 25930 16516
rect 25961 16507 26019 16513
rect 25961 16473 25973 16507
rect 26007 16504 26019 16507
rect 26234 16504 26240 16516
rect 26007 16476 26240 16504
rect 26007 16473 26019 16476
rect 25961 16467 26019 16473
rect 26234 16464 26240 16476
rect 26292 16464 26298 16516
rect 28353 16507 28411 16513
rect 28353 16473 28365 16507
rect 28399 16504 28411 16507
rect 28626 16504 28632 16516
rect 28399 16476 28632 16504
rect 28399 16473 28411 16476
rect 28353 16467 28411 16473
rect 28626 16464 28632 16476
rect 28684 16464 28690 16516
rect 22005 16439 22063 16445
rect 22005 16405 22017 16439
rect 22051 16436 22063 16439
rect 22554 16436 22560 16448
rect 22051 16408 22560 16436
rect 22051 16405 22063 16408
rect 22005 16399 22063 16405
rect 22554 16396 22560 16408
rect 22612 16396 22618 16448
rect 23658 16436 23664 16448
rect 23619 16408 23664 16436
rect 23658 16396 23664 16408
rect 23716 16396 23722 16448
rect 1104 16346 29048 16368
rect 1104 16294 7896 16346
rect 7948 16294 7960 16346
rect 8012 16294 8024 16346
rect 8076 16294 8088 16346
rect 8140 16294 8152 16346
rect 8204 16294 14842 16346
rect 14894 16294 14906 16346
rect 14958 16294 14970 16346
rect 15022 16294 15034 16346
rect 15086 16294 15098 16346
rect 15150 16294 21788 16346
rect 21840 16294 21852 16346
rect 21904 16294 21916 16346
rect 21968 16294 21980 16346
rect 22032 16294 22044 16346
rect 22096 16294 28734 16346
rect 28786 16294 28798 16346
rect 28850 16294 28862 16346
rect 28914 16294 28926 16346
rect 28978 16294 28990 16346
rect 29042 16294 29048 16346
rect 1104 16272 29048 16294
rect 11974 16192 11980 16244
rect 12032 16232 12038 16244
rect 20625 16235 20683 16241
rect 12032 16204 18184 16232
rect 12032 16192 12038 16204
rect 18046 16164 18052 16176
rect 16868 16136 18052 16164
rect 1670 16096 1676 16108
rect 1631 16068 1676 16096
rect 1670 16056 1676 16068
rect 1728 16056 1734 16108
rect 16868 16105 16896 16136
rect 18046 16124 18052 16136
rect 18104 16124 18110 16176
rect 18156 16164 18184 16204
rect 20625 16201 20637 16235
rect 20671 16232 20683 16235
rect 20714 16232 20720 16244
rect 20671 16204 20720 16232
rect 20671 16201 20683 16204
rect 20625 16195 20683 16201
rect 20714 16192 20720 16204
rect 20772 16192 20778 16244
rect 26234 16192 26240 16244
rect 26292 16232 26298 16244
rect 28169 16235 28227 16241
rect 28169 16232 28181 16235
rect 26292 16204 28181 16232
rect 26292 16192 26298 16204
rect 28169 16201 28181 16204
rect 28215 16201 28227 16235
rect 28169 16195 28227 16201
rect 24854 16164 24860 16176
rect 18156 16136 24860 16164
rect 24854 16124 24860 16136
rect 24912 16124 24918 16176
rect 17126 16105 17132 16108
rect 16853 16099 16911 16105
rect 16853 16065 16865 16099
rect 16899 16065 16911 16099
rect 16853 16059 16911 16065
rect 17120 16059 17132 16105
rect 17184 16096 17190 16108
rect 20441 16099 20499 16105
rect 17184 16068 17220 16096
rect 17126 16056 17132 16059
rect 17184 16056 17190 16068
rect 20441 16065 20453 16099
rect 20487 16096 20499 16099
rect 21085 16099 21143 16105
rect 21085 16096 21097 16099
rect 20487 16068 21097 16096
rect 20487 16065 20499 16068
rect 20441 16059 20499 16065
rect 21085 16065 21097 16068
rect 21131 16065 21143 16099
rect 21266 16096 21272 16108
rect 21227 16068 21272 16096
rect 21085 16059 21143 16065
rect 21266 16056 21272 16068
rect 21324 16056 21330 16108
rect 21450 16096 21456 16108
rect 21411 16068 21456 16096
rect 21450 16056 21456 16068
rect 21508 16056 21514 16108
rect 26234 16096 26240 16108
rect 26195 16068 26240 16096
rect 26234 16056 26240 16068
rect 26292 16056 26298 16108
rect 26421 16099 26479 16105
rect 26421 16065 26433 16099
rect 26467 16096 26479 16099
rect 27341 16099 27399 16105
rect 27341 16096 27353 16099
rect 26467 16068 27353 16096
rect 26467 16065 26479 16068
rect 26421 16059 26479 16065
rect 27341 16065 27353 16068
rect 27387 16065 27399 16099
rect 27341 16059 27399 16065
rect 28353 16099 28411 16105
rect 28353 16065 28365 16099
rect 28399 16096 28411 16099
rect 29914 16096 29920 16108
rect 28399 16068 29920 16096
rect 28399 16065 28411 16068
rect 28353 16059 28411 16065
rect 29914 16056 29920 16068
rect 29972 16056 29978 16108
rect 1857 16031 1915 16037
rect 1857 15997 1869 16031
rect 1903 16028 1915 16031
rect 2222 16028 2228 16040
rect 1903 16000 2228 16028
rect 1903 15997 1915 16000
rect 1857 15991 1915 15997
rect 2222 15988 2228 16000
rect 2280 15988 2286 16040
rect 2774 16028 2780 16040
rect 2735 16000 2780 16028
rect 2774 15988 2780 16000
rect 2832 15988 2838 16040
rect 25958 15988 25964 16040
rect 26016 16028 26022 16040
rect 26053 16031 26111 16037
rect 26053 16028 26065 16031
rect 26016 16000 26065 16028
rect 26016 15988 26022 16000
rect 26053 15997 26065 16000
rect 26099 15997 26111 16031
rect 26053 15991 26111 15997
rect 17218 15852 17224 15904
rect 17276 15892 17282 15904
rect 18233 15895 18291 15901
rect 18233 15892 18245 15895
rect 17276 15864 18245 15892
rect 17276 15852 17282 15864
rect 18233 15861 18245 15864
rect 18279 15861 18291 15895
rect 27154 15892 27160 15904
rect 27115 15864 27160 15892
rect 18233 15855 18291 15861
rect 27154 15852 27160 15864
rect 27212 15852 27218 15904
rect 1104 15802 28888 15824
rect 1104 15750 4423 15802
rect 4475 15750 4487 15802
rect 4539 15750 4551 15802
rect 4603 15750 4615 15802
rect 4667 15750 4679 15802
rect 4731 15750 11369 15802
rect 11421 15750 11433 15802
rect 11485 15750 11497 15802
rect 11549 15750 11561 15802
rect 11613 15750 11625 15802
rect 11677 15750 18315 15802
rect 18367 15750 18379 15802
rect 18431 15750 18443 15802
rect 18495 15750 18507 15802
rect 18559 15750 18571 15802
rect 18623 15750 25261 15802
rect 25313 15750 25325 15802
rect 25377 15750 25389 15802
rect 25441 15750 25453 15802
rect 25505 15750 25517 15802
rect 25569 15750 28888 15802
rect 1104 15728 28888 15750
rect 2222 15688 2228 15700
rect 2183 15660 2228 15688
rect 2222 15648 2228 15660
rect 2280 15648 2286 15700
rect 20806 15688 20812 15700
rect 20767 15660 20812 15688
rect 20806 15648 20812 15660
rect 20864 15648 20870 15700
rect 10781 15555 10839 15561
rect 10781 15521 10793 15555
rect 10827 15552 10839 15555
rect 12989 15555 13047 15561
rect 12989 15552 13001 15555
rect 10827 15524 13001 15552
rect 10827 15521 10839 15524
rect 10781 15515 10839 15521
rect 12989 15521 13001 15524
rect 13035 15521 13047 15555
rect 12989 15515 13047 15521
rect 13173 15555 13231 15561
rect 13173 15521 13185 15555
rect 13219 15552 13231 15555
rect 13446 15552 13452 15564
rect 13219 15524 13452 15552
rect 13219 15521 13231 15524
rect 13173 15515 13231 15521
rect 13446 15512 13452 15524
rect 13504 15512 13510 15564
rect 21634 15552 21640 15564
rect 21595 15524 21640 15552
rect 21634 15512 21640 15524
rect 21692 15512 21698 15564
rect 25038 15512 25044 15564
rect 25096 15552 25102 15564
rect 26050 15552 26056 15564
rect 25096 15524 26056 15552
rect 25096 15512 25102 15524
rect 26050 15512 26056 15524
rect 26108 15552 26114 15564
rect 26145 15555 26203 15561
rect 26145 15552 26157 15555
rect 26108 15524 26157 15552
rect 26108 15512 26114 15524
rect 26145 15521 26157 15524
rect 26191 15521 26203 15555
rect 26145 15515 26203 15521
rect 2314 15484 2320 15496
rect 2275 15456 2320 15484
rect 2314 15444 2320 15456
rect 2372 15444 2378 15496
rect 10686 15484 10692 15496
rect 10599 15456 10692 15484
rect 10686 15444 10692 15456
rect 10744 15484 10750 15496
rect 17221 15487 17279 15493
rect 10744 15456 11836 15484
rect 10744 15444 10750 15456
rect 11054 15376 11060 15428
rect 11112 15416 11118 15428
rect 11333 15419 11391 15425
rect 11333 15416 11345 15419
rect 11112 15388 11345 15416
rect 11112 15376 11118 15388
rect 11333 15385 11345 15388
rect 11379 15385 11391 15419
rect 11808 15416 11836 15456
rect 17221 15453 17233 15487
rect 17267 15484 17279 15487
rect 18046 15484 18052 15496
rect 17267 15456 18052 15484
rect 17267 15453 17279 15456
rect 17221 15447 17279 15453
rect 18046 15444 18052 15456
rect 18104 15484 18110 15496
rect 19242 15484 19248 15496
rect 18104 15456 19248 15484
rect 18104 15444 18110 15456
rect 19242 15444 19248 15456
rect 19300 15484 19306 15496
rect 19429 15487 19487 15493
rect 19429 15484 19441 15487
rect 19300 15456 19441 15484
rect 19300 15444 19306 15456
rect 19429 15453 19441 15456
rect 19475 15453 19487 15487
rect 25498 15484 25504 15496
rect 25459 15456 25504 15484
rect 19429 15447 19487 15453
rect 25498 15444 25504 15456
rect 25556 15444 25562 15496
rect 26412 15487 26470 15493
rect 26412 15453 26424 15487
rect 26458 15484 26470 15487
rect 27154 15484 27160 15496
rect 26458 15456 27160 15484
rect 26458 15453 26470 15456
rect 26412 15447 26470 15453
rect 27154 15444 27160 15456
rect 27212 15444 27218 15496
rect 27985 15487 28043 15493
rect 27985 15453 27997 15487
rect 28031 15484 28043 15487
rect 28074 15484 28080 15496
rect 28031 15456 28080 15484
rect 28031 15453 28043 15456
rect 27985 15447 28043 15453
rect 28074 15444 28080 15456
rect 28132 15444 28138 15496
rect 11974 15416 11980 15428
rect 11808 15388 11980 15416
rect 11333 15379 11391 15385
rect 11974 15376 11980 15388
rect 12032 15376 12038 15428
rect 17310 15376 17316 15428
rect 17368 15416 17374 15428
rect 19702 15425 19708 15428
rect 17466 15419 17524 15425
rect 17466 15416 17478 15419
rect 17368 15388 17478 15416
rect 17368 15376 17374 15388
rect 17466 15385 17478 15388
rect 17512 15385 17524 15419
rect 17466 15379 17524 15385
rect 19696 15379 19708 15425
rect 19760 15416 19766 15428
rect 19760 15388 19796 15416
rect 19702 15376 19708 15379
rect 19760 15376 19766 15388
rect 21542 15376 21548 15428
rect 21600 15416 21606 15428
rect 21882 15419 21940 15425
rect 21882 15416 21894 15419
rect 21600 15388 21894 15416
rect 21600 15376 21606 15388
rect 21882 15385 21894 15388
rect 21928 15385 21940 15419
rect 21882 15379 21940 15385
rect 18601 15351 18659 15357
rect 18601 15317 18613 15351
rect 18647 15348 18659 15351
rect 18690 15348 18696 15360
rect 18647 15320 18696 15348
rect 18647 15317 18659 15320
rect 18601 15311 18659 15317
rect 18690 15308 18696 15320
rect 18748 15308 18754 15360
rect 23014 15348 23020 15360
rect 22975 15320 23020 15348
rect 23014 15308 23020 15320
rect 23072 15308 23078 15360
rect 25685 15351 25743 15357
rect 25685 15317 25697 15351
rect 25731 15348 25743 15351
rect 27338 15348 27344 15360
rect 25731 15320 27344 15348
rect 25731 15317 25743 15320
rect 25685 15311 25743 15317
rect 27338 15308 27344 15320
rect 27396 15308 27402 15360
rect 27430 15308 27436 15360
rect 27488 15348 27494 15360
rect 27525 15351 27583 15357
rect 27525 15348 27537 15351
rect 27488 15320 27537 15348
rect 27488 15308 27494 15320
rect 27525 15317 27537 15320
rect 27571 15317 27583 15351
rect 27525 15311 27583 15317
rect 28077 15351 28135 15357
rect 28077 15317 28089 15351
rect 28123 15348 28135 15351
rect 28166 15348 28172 15360
rect 28123 15320 28172 15348
rect 28123 15317 28135 15320
rect 28077 15311 28135 15317
rect 28166 15308 28172 15320
rect 28224 15308 28230 15360
rect 1104 15258 29048 15280
rect 1104 15206 7896 15258
rect 7948 15206 7960 15258
rect 8012 15206 8024 15258
rect 8076 15206 8088 15258
rect 8140 15206 8152 15258
rect 8204 15206 14842 15258
rect 14894 15206 14906 15258
rect 14958 15206 14970 15258
rect 15022 15206 15034 15258
rect 15086 15206 15098 15258
rect 15150 15206 21788 15258
rect 21840 15206 21852 15258
rect 21904 15206 21916 15258
rect 21968 15206 21980 15258
rect 22032 15206 22044 15258
rect 22096 15206 28734 15258
rect 28786 15206 28798 15258
rect 28850 15206 28862 15258
rect 28914 15206 28926 15258
rect 28978 15206 28990 15258
rect 29042 15206 29048 15258
rect 1104 15184 29048 15206
rect 20438 15104 20444 15156
rect 20496 15144 20502 15156
rect 20622 15144 20628 15156
rect 20496 15116 20628 15144
rect 20496 15104 20502 15116
rect 20622 15104 20628 15116
rect 20680 15144 20686 15156
rect 20680 15116 21036 15144
rect 20680 15104 20686 15116
rect 19242 15036 19248 15088
rect 19300 15076 19306 15088
rect 21008 15076 21036 15116
rect 21266 15104 21272 15156
rect 21324 15144 21330 15156
rect 22005 15147 22063 15153
rect 22005 15144 22017 15147
rect 21324 15116 22017 15144
rect 21324 15104 21330 15116
rect 22005 15113 22017 15116
rect 22051 15113 22063 15147
rect 22005 15107 22063 15113
rect 22373 15147 22431 15153
rect 22373 15113 22385 15147
rect 22419 15144 22431 15147
rect 22554 15144 22560 15156
rect 22419 15116 22560 15144
rect 22419 15113 22431 15116
rect 22373 15107 22431 15113
rect 22554 15104 22560 15116
rect 22612 15104 22618 15156
rect 23106 15104 23112 15156
rect 23164 15144 23170 15156
rect 23201 15147 23259 15153
rect 23201 15144 23213 15147
rect 23164 15116 23213 15144
rect 23164 15104 23170 15116
rect 23201 15113 23213 15116
rect 23247 15113 23259 15147
rect 23201 15107 23259 15113
rect 26234 15104 26240 15156
rect 26292 15144 26298 15156
rect 27157 15147 27215 15153
rect 27157 15144 27169 15147
rect 26292 15116 27169 15144
rect 26292 15104 26298 15116
rect 27157 15113 27169 15116
rect 27203 15113 27215 15147
rect 27157 15107 27215 15113
rect 27338 15104 27344 15156
rect 27396 15144 27402 15156
rect 27617 15147 27675 15153
rect 27617 15144 27629 15147
rect 27396 15116 27629 15144
rect 27396 15104 27402 15116
rect 27617 15113 27629 15116
rect 27663 15113 27675 15147
rect 27617 15107 27675 15113
rect 19300 15048 20668 15076
rect 21008 15048 22600 15076
rect 19300 15036 19306 15048
rect 17954 15008 17960 15020
rect 18012 15017 18018 15020
rect 17924 14980 17960 15008
rect 17954 14968 17960 14980
rect 18012 14971 18024 15017
rect 18012 14968 18018 14971
rect 18138 14968 18144 15020
rect 18196 15008 18202 15020
rect 18233 15011 18291 15017
rect 18233 15008 18245 15011
rect 18196 14980 18245 15008
rect 18196 14968 18202 14980
rect 18233 14977 18245 14980
rect 18279 14977 18291 15011
rect 20346 15008 20352 15020
rect 20404 15017 20410 15020
rect 20640 15017 20668 15048
rect 20316 14980 20352 15008
rect 18233 14971 18291 14977
rect 20346 14968 20352 14980
rect 20404 14971 20416 15017
rect 20625 15011 20683 15017
rect 20625 14977 20637 15011
rect 20671 14977 20683 15011
rect 20625 14971 20683 14977
rect 20404 14968 20410 14971
rect 22572 14949 22600 15048
rect 23658 15036 23664 15088
rect 23716 15076 23722 15088
rect 24314 15079 24372 15085
rect 24314 15076 24326 15079
rect 23716 15048 24326 15076
rect 23716 15036 23722 15048
rect 24314 15045 24326 15048
rect 24360 15045 24372 15079
rect 24314 15039 24372 15045
rect 26050 15036 26056 15088
rect 26108 15076 26114 15088
rect 26108 15048 26464 15076
rect 26108 15036 26114 15048
rect 24581 15011 24639 15017
rect 24581 14977 24593 15011
rect 24627 15008 24639 15011
rect 25038 15008 25044 15020
rect 24627 14980 25044 15008
rect 24627 14977 24639 14980
rect 24581 14971 24639 14977
rect 25038 14968 25044 14980
rect 25096 14968 25102 15020
rect 25130 14968 25136 15020
rect 25188 15008 25194 15020
rect 26436 15017 26464 15048
rect 26154 15011 26212 15017
rect 26154 15008 26166 15011
rect 25188 14980 26166 15008
rect 25188 14968 25194 14980
rect 26154 14977 26166 14980
rect 26200 14977 26212 15011
rect 26154 14971 26212 14977
rect 26421 15011 26479 15017
rect 26421 14977 26433 15011
rect 26467 14977 26479 15011
rect 26421 14971 26479 14977
rect 27430 14968 27436 15020
rect 27488 15008 27494 15020
rect 27525 15011 27583 15017
rect 27525 15008 27537 15011
rect 27488 14980 27537 15008
rect 27488 14968 27494 14980
rect 27525 14977 27537 14980
rect 27571 14977 27583 15011
rect 27525 14971 27583 14977
rect 22465 14943 22523 14949
rect 22465 14909 22477 14943
rect 22511 14909 22523 14943
rect 22465 14903 22523 14909
rect 22557 14943 22615 14949
rect 22557 14909 22569 14943
rect 22603 14909 22615 14943
rect 22557 14903 22615 14909
rect 19245 14875 19303 14881
rect 19245 14841 19257 14875
rect 19291 14872 19303 14875
rect 19334 14872 19340 14884
rect 19291 14844 19340 14872
rect 19291 14841 19303 14844
rect 19245 14835 19303 14841
rect 19334 14832 19340 14844
rect 19392 14832 19398 14884
rect 22480 14872 22508 14903
rect 27338 14900 27344 14952
rect 27396 14940 27402 14952
rect 27709 14943 27767 14949
rect 27709 14940 27721 14943
rect 27396 14912 27721 14940
rect 27396 14900 27402 14912
rect 27709 14909 27721 14912
rect 27755 14909 27767 14943
rect 27709 14903 27767 14909
rect 22738 14872 22744 14884
rect 22480 14844 22744 14872
rect 22738 14832 22744 14844
rect 22796 14872 22802 14884
rect 23290 14872 23296 14884
rect 22796 14844 23296 14872
rect 22796 14832 22802 14844
rect 23290 14832 23296 14844
rect 23348 14832 23354 14884
rect 16206 14764 16212 14816
rect 16264 14804 16270 14816
rect 16853 14807 16911 14813
rect 16853 14804 16865 14807
rect 16264 14776 16865 14804
rect 16264 14764 16270 14776
rect 16853 14773 16865 14776
rect 16899 14773 16911 14807
rect 19352 14804 19380 14832
rect 21450 14804 21456 14816
rect 19352 14776 21456 14804
rect 16853 14767 16911 14773
rect 21450 14764 21456 14776
rect 21508 14764 21514 14816
rect 24210 14764 24216 14816
rect 24268 14804 24274 14816
rect 25041 14807 25099 14813
rect 25041 14804 25053 14807
rect 24268 14776 25053 14804
rect 24268 14764 24274 14776
rect 25041 14773 25053 14776
rect 25087 14773 25099 14807
rect 25041 14767 25099 14773
rect 1104 14714 28888 14736
rect 1104 14662 4423 14714
rect 4475 14662 4487 14714
rect 4539 14662 4551 14714
rect 4603 14662 4615 14714
rect 4667 14662 4679 14714
rect 4731 14662 11369 14714
rect 11421 14662 11433 14714
rect 11485 14662 11497 14714
rect 11549 14662 11561 14714
rect 11613 14662 11625 14714
rect 11677 14662 18315 14714
rect 18367 14662 18379 14714
rect 18431 14662 18443 14714
rect 18495 14662 18507 14714
rect 18559 14662 18571 14714
rect 18623 14662 25261 14714
rect 25313 14662 25325 14714
rect 25377 14662 25389 14714
rect 25441 14662 25453 14714
rect 25505 14662 25517 14714
rect 25569 14662 28888 14714
rect 1104 14640 28888 14662
rect 16393 14603 16451 14609
rect 16393 14569 16405 14603
rect 16439 14600 16451 14603
rect 17037 14603 17095 14609
rect 17037 14600 17049 14603
rect 16439 14572 17049 14600
rect 16439 14569 16451 14572
rect 16393 14563 16451 14569
rect 17037 14569 17049 14572
rect 17083 14569 17095 14603
rect 17037 14563 17095 14569
rect 17865 14603 17923 14609
rect 17865 14569 17877 14603
rect 17911 14600 17923 14603
rect 17954 14600 17960 14612
rect 17911 14572 17960 14600
rect 17911 14569 17923 14572
rect 17865 14563 17923 14569
rect 17954 14560 17960 14572
rect 18012 14560 18018 14612
rect 19613 14603 19671 14609
rect 19613 14569 19625 14603
rect 19659 14600 19671 14603
rect 19702 14600 19708 14612
rect 19659 14572 19708 14600
rect 19659 14569 19671 14572
rect 19613 14563 19671 14569
rect 19702 14560 19708 14572
rect 19760 14560 19766 14612
rect 17402 14464 17408 14476
rect 17068 14436 17408 14464
rect 3418 14356 3424 14408
rect 3476 14396 3482 14408
rect 3476 14368 3521 14396
rect 3476 14356 3482 14368
rect 15654 14356 15660 14408
rect 15712 14396 15718 14408
rect 16025 14399 16083 14405
rect 16025 14396 16037 14399
rect 15712 14368 16037 14396
rect 15712 14356 15718 14368
rect 16025 14365 16037 14368
rect 16071 14396 16083 14399
rect 16114 14396 16120 14408
rect 16071 14368 16120 14396
rect 16071 14365 16083 14368
rect 16025 14359 16083 14365
rect 16114 14356 16120 14368
rect 16172 14356 16178 14408
rect 1578 14328 1584 14340
rect 1539 14300 1584 14328
rect 1578 14288 1584 14300
rect 1636 14288 1642 14340
rect 2866 14288 2872 14340
rect 2924 14328 2930 14340
rect 3237 14331 3295 14337
rect 3237 14328 3249 14331
rect 2924 14300 3249 14328
rect 2924 14288 2930 14300
rect 3237 14297 3249 14300
rect 3283 14297 3295 14331
rect 16206 14328 16212 14340
rect 16167 14300 16212 14328
rect 3237 14291 3295 14297
rect 16206 14288 16212 14300
rect 16264 14288 16270 14340
rect 16850 14328 16856 14340
rect 16811 14300 16856 14328
rect 16850 14288 16856 14300
rect 16908 14288 16914 14340
rect 16298 14220 16304 14272
rect 16356 14260 16362 14272
rect 17068 14269 17096 14436
rect 17402 14424 17408 14436
rect 17460 14424 17466 14476
rect 26050 14464 26056 14476
rect 26011 14436 26056 14464
rect 26050 14424 26056 14436
rect 26108 14424 26114 14476
rect 27522 14464 27528 14476
rect 27483 14436 27528 14464
rect 27522 14424 27528 14436
rect 27580 14424 27586 14476
rect 28166 14464 28172 14476
rect 28127 14436 28172 14464
rect 28166 14424 28172 14436
rect 28224 14424 28230 14476
rect 17681 14399 17739 14405
rect 17681 14396 17693 14399
rect 17236 14368 17693 14396
rect 17236 14269 17264 14368
rect 17681 14365 17693 14368
rect 17727 14365 17739 14399
rect 19426 14396 19432 14408
rect 19387 14368 19432 14396
rect 17681 14359 17739 14365
rect 19426 14356 19432 14368
rect 19484 14356 19490 14408
rect 28350 14356 28356 14408
rect 28408 14396 28414 14408
rect 28408 14368 28453 14396
rect 28408 14356 28414 14368
rect 25774 14328 25780 14340
rect 25832 14337 25838 14340
rect 25744 14300 25780 14328
rect 25774 14288 25780 14300
rect 25832 14291 25844 14337
rect 25832 14288 25838 14291
rect 17053 14263 17111 14269
rect 17053 14260 17065 14263
rect 16356 14232 17065 14260
rect 16356 14220 16362 14232
rect 17053 14229 17065 14232
rect 17099 14229 17111 14263
rect 17053 14223 17111 14229
rect 17221 14263 17279 14269
rect 17221 14229 17233 14263
rect 17267 14229 17279 14263
rect 17221 14223 17279 14229
rect 24302 14220 24308 14272
rect 24360 14260 24366 14272
rect 24673 14263 24731 14269
rect 24673 14260 24685 14263
rect 24360 14232 24685 14260
rect 24360 14220 24366 14232
rect 24673 14229 24685 14232
rect 24719 14260 24731 14263
rect 26234 14260 26240 14272
rect 24719 14232 26240 14260
rect 24719 14229 24731 14232
rect 24673 14223 24731 14229
rect 26234 14220 26240 14232
rect 26292 14220 26298 14272
rect 1104 14170 29048 14192
rect 1104 14118 7896 14170
rect 7948 14118 7960 14170
rect 8012 14118 8024 14170
rect 8076 14118 8088 14170
rect 8140 14118 8152 14170
rect 8204 14118 14842 14170
rect 14894 14118 14906 14170
rect 14958 14118 14970 14170
rect 15022 14118 15034 14170
rect 15086 14118 15098 14170
rect 15150 14118 21788 14170
rect 21840 14118 21852 14170
rect 21904 14118 21916 14170
rect 21968 14118 21980 14170
rect 22032 14118 22044 14170
rect 22096 14118 28734 14170
rect 28786 14118 28798 14170
rect 28850 14118 28862 14170
rect 28914 14118 28926 14170
rect 28978 14118 28990 14170
rect 29042 14118 29048 14170
rect 1104 14096 29048 14118
rect 2866 14056 2872 14068
rect 2827 14028 2872 14056
rect 2866 14016 2872 14028
rect 2924 14016 2930 14068
rect 16298 14056 16304 14068
rect 16259 14028 16304 14056
rect 16298 14016 16304 14028
rect 16356 14016 16362 14068
rect 17129 14059 17187 14065
rect 17129 14025 17141 14059
rect 17175 14056 17187 14059
rect 17310 14056 17316 14068
rect 17175 14028 17316 14056
rect 17175 14025 17187 14028
rect 17129 14019 17187 14025
rect 17310 14016 17316 14028
rect 17368 14016 17374 14068
rect 19426 14056 19432 14068
rect 19387 14028 19432 14056
rect 19426 14016 19432 14028
rect 19484 14016 19490 14068
rect 20257 14059 20315 14065
rect 20257 14025 20269 14059
rect 20303 14056 20315 14059
rect 20346 14056 20352 14068
rect 20303 14028 20352 14056
rect 20303 14025 20315 14028
rect 20257 14019 20315 14025
rect 20346 14016 20352 14028
rect 20404 14016 20410 14068
rect 22738 14016 22744 14068
rect 22796 14056 22802 14068
rect 23125 14059 23183 14065
rect 23125 14056 23137 14059
rect 22796 14028 23137 14056
rect 22796 14016 22802 14028
rect 23125 14025 23137 14028
rect 23171 14025 23183 14059
rect 23125 14019 23183 14025
rect 23474 14016 23480 14068
rect 23532 14056 23538 14068
rect 23750 14056 23756 14068
rect 23532 14028 23756 14056
rect 23532 14016 23538 14028
rect 23750 14016 23756 14028
rect 23808 14056 23814 14068
rect 23845 14059 23903 14065
rect 23845 14056 23857 14059
rect 23808 14028 23857 14056
rect 23808 14016 23814 14028
rect 23845 14025 23857 14028
rect 23891 14025 23903 14059
rect 23845 14019 23903 14025
rect 23937 14059 23995 14065
rect 23937 14025 23949 14059
rect 23983 14056 23995 14059
rect 24026 14056 24032 14068
rect 23983 14028 24032 14056
rect 23983 14025 23995 14028
rect 23937 14019 23995 14025
rect 24026 14016 24032 14028
rect 24084 14016 24090 14068
rect 24765 14059 24823 14065
rect 24765 14025 24777 14059
rect 24811 14056 24823 14059
rect 25130 14056 25136 14068
rect 24811 14028 25136 14056
rect 24811 14025 24823 14028
rect 24765 14019 24823 14025
rect 25130 14016 25136 14028
rect 25188 14016 25194 14068
rect 25774 14056 25780 14068
rect 25735 14028 25780 14056
rect 25774 14016 25780 14028
rect 25832 14016 25838 14068
rect 3418 13988 3424 14000
rect 2332 13960 3424 13988
rect 2332 13929 2360 13960
rect 3418 13948 3424 13960
rect 3476 13948 3482 14000
rect 22925 13991 22983 13997
rect 22925 13957 22937 13991
rect 22971 13988 22983 13991
rect 23014 13988 23020 14000
rect 22971 13960 23020 13988
rect 22971 13957 22983 13960
rect 22925 13951 22983 13957
rect 23014 13948 23020 13960
rect 23072 13948 23078 14000
rect 2317 13923 2375 13929
rect 2317 13889 2329 13923
rect 2363 13889 2375 13923
rect 2958 13920 2964 13932
rect 2919 13892 2964 13920
rect 2317 13883 2375 13889
rect 2958 13880 2964 13892
rect 3016 13880 3022 13932
rect 16114 13920 16120 13932
rect 16075 13892 16120 13920
rect 16114 13880 16120 13892
rect 16172 13880 16178 13932
rect 16206 13880 16212 13932
rect 16264 13920 16270 13932
rect 16301 13923 16359 13929
rect 16301 13920 16313 13923
rect 16264 13892 16313 13920
rect 16264 13880 16270 13892
rect 16301 13889 16313 13892
rect 16347 13920 16359 13923
rect 16347 13892 16988 13920
rect 16347 13889 16359 13892
rect 16301 13883 16359 13889
rect 16850 13852 16856 13864
rect 16811 13824 16856 13852
rect 16850 13812 16856 13824
rect 16908 13812 16914 13864
rect 16960 13852 16988 13892
rect 17034 13880 17040 13932
rect 17092 13920 17098 13932
rect 17221 13923 17279 13929
rect 17221 13920 17233 13923
rect 17092 13892 17233 13920
rect 17092 13880 17098 13892
rect 17221 13889 17233 13892
rect 17267 13889 17279 13923
rect 17221 13883 17279 13889
rect 17313 13923 17371 13929
rect 17313 13889 17325 13923
rect 17359 13920 17371 13923
rect 17402 13920 17408 13932
rect 17359 13892 17408 13920
rect 17359 13889 17371 13892
rect 17313 13883 17371 13889
rect 17402 13880 17408 13892
rect 17460 13880 17466 13932
rect 17865 13923 17923 13929
rect 17865 13889 17877 13923
rect 17911 13889 17923 13923
rect 17865 13883 17923 13889
rect 18509 13923 18567 13929
rect 18509 13889 18521 13923
rect 18555 13920 18567 13923
rect 18690 13920 18696 13932
rect 18555 13892 18696 13920
rect 18555 13889 18567 13892
rect 18509 13883 18567 13889
rect 17880 13852 17908 13883
rect 18690 13880 18696 13892
rect 18748 13880 18754 13932
rect 19610 13920 19616 13932
rect 19571 13892 19616 13920
rect 19610 13880 19616 13892
rect 19668 13880 19674 13932
rect 19797 13923 19855 13929
rect 19797 13889 19809 13923
rect 19843 13920 19855 13923
rect 19886 13920 19892 13932
rect 19843 13892 19892 13920
rect 19843 13889 19855 13892
rect 19797 13883 19855 13889
rect 19886 13880 19892 13892
rect 19944 13880 19950 13932
rect 20438 13920 20444 13932
rect 20399 13892 20444 13920
rect 20438 13880 20444 13892
rect 20496 13880 20502 13932
rect 23750 13920 23756 13932
rect 23711 13892 23756 13920
rect 23750 13880 23756 13892
rect 23808 13880 23814 13932
rect 24121 13923 24179 13929
rect 24121 13889 24133 13923
rect 24167 13920 24179 13923
rect 24210 13920 24216 13932
rect 24167 13892 24216 13920
rect 24167 13889 24179 13892
rect 24121 13883 24179 13889
rect 16960 13824 17356 13852
rect 17328 13784 17356 13824
rect 17512 13824 17908 13852
rect 17512 13784 17540 13824
rect 21634 13812 21640 13864
rect 21692 13852 21698 13864
rect 22005 13855 22063 13861
rect 22005 13852 22017 13855
rect 21692 13824 22017 13852
rect 21692 13812 21698 13824
rect 22005 13821 22017 13824
rect 22051 13821 22063 13855
rect 22462 13852 22468 13864
rect 22423 13824 22468 13852
rect 22005 13815 22063 13821
rect 22462 13812 22468 13824
rect 22520 13812 22526 13864
rect 23658 13812 23664 13864
rect 23716 13852 23722 13864
rect 24136 13852 24164 13883
rect 24210 13880 24216 13892
rect 24268 13880 24274 13932
rect 24578 13920 24584 13932
rect 24539 13892 24584 13920
rect 24578 13880 24584 13892
rect 24636 13880 24642 13932
rect 25590 13920 25596 13932
rect 25551 13892 25596 13920
rect 25590 13880 25596 13892
rect 25648 13880 25654 13932
rect 28077 13923 28135 13929
rect 28077 13889 28089 13923
rect 28123 13920 28135 13923
rect 28350 13920 28356 13932
rect 28123 13892 28356 13920
rect 28123 13889 28135 13892
rect 28077 13883 28135 13889
rect 28350 13880 28356 13892
rect 28408 13880 28414 13932
rect 23716 13824 24164 13852
rect 23716 13812 23722 13824
rect 17328 13756 17540 13784
rect 18138 13744 18144 13796
rect 18196 13784 18202 13796
rect 18601 13787 18659 13793
rect 18601 13784 18613 13787
rect 18196 13756 18613 13784
rect 18196 13744 18202 13756
rect 18601 13753 18613 13756
rect 18647 13753 18659 13787
rect 18601 13747 18659 13753
rect 22189 13787 22247 13793
rect 22189 13753 22201 13787
rect 22235 13784 22247 13787
rect 22278 13784 22284 13796
rect 22235 13756 22284 13784
rect 22235 13753 22247 13756
rect 22189 13747 22247 13753
rect 22278 13744 22284 13756
rect 22336 13744 22342 13796
rect 24302 13784 24308 13796
rect 23032 13756 24308 13784
rect 3418 13716 3424 13728
rect 3379 13688 3424 13716
rect 3418 13676 3424 13688
rect 3476 13676 3482 13728
rect 17954 13716 17960 13728
rect 17915 13688 17960 13716
rect 17954 13676 17960 13688
rect 18012 13676 18018 13728
rect 18046 13676 18052 13728
rect 18104 13716 18110 13728
rect 23032 13716 23060 13756
rect 24302 13744 24308 13756
rect 24360 13744 24366 13796
rect 18104 13688 23060 13716
rect 18104 13676 18110 13688
rect 23106 13676 23112 13728
rect 23164 13716 23170 13728
rect 23164 13688 23209 13716
rect 23164 13676 23170 13688
rect 23290 13676 23296 13728
rect 23348 13716 23354 13728
rect 24029 13719 24087 13725
rect 23348 13688 23393 13716
rect 23348 13676 23354 13688
rect 24029 13685 24041 13719
rect 24075 13716 24087 13719
rect 24670 13716 24676 13728
rect 24075 13688 24676 13716
rect 24075 13685 24087 13688
rect 24029 13679 24087 13685
rect 24670 13676 24676 13688
rect 24728 13676 24734 13728
rect 1104 13626 28888 13648
rect 1104 13574 4423 13626
rect 4475 13574 4487 13626
rect 4539 13574 4551 13626
rect 4603 13574 4615 13626
rect 4667 13574 4679 13626
rect 4731 13574 11369 13626
rect 11421 13574 11433 13626
rect 11485 13574 11497 13626
rect 11549 13574 11561 13626
rect 11613 13574 11625 13626
rect 11677 13574 18315 13626
rect 18367 13574 18379 13626
rect 18431 13574 18443 13626
rect 18495 13574 18507 13626
rect 18559 13574 18571 13626
rect 18623 13574 25261 13626
rect 25313 13574 25325 13626
rect 25377 13574 25389 13626
rect 25441 13574 25453 13626
rect 25505 13574 25517 13626
rect 25569 13574 28888 13626
rect 1104 13552 28888 13574
rect 18046 13512 18052 13524
rect 18007 13484 18052 13512
rect 18046 13472 18052 13484
rect 18104 13472 18110 13524
rect 19610 13472 19616 13524
rect 19668 13512 19674 13524
rect 19889 13515 19947 13521
rect 19889 13512 19901 13515
rect 19668 13484 19901 13512
rect 19668 13472 19674 13484
rect 19889 13481 19901 13484
rect 19935 13481 19947 13515
rect 22278 13512 22284 13524
rect 22239 13484 22284 13512
rect 19889 13475 19947 13481
rect 22278 13472 22284 13484
rect 22336 13472 22342 13524
rect 23290 13472 23296 13524
rect 23348 13512 23354 13524
rect 24578 13512 24584 13524
rect 23348 13484 23796 13512
rect 24539 13484 24584 13512
rect 23348 13472 23354 13484
rect 23658 13444 23664 13456
rect 20364 13416 23664 13444
rect 1578 13376 1584 13388
rect 1539 13348 1584 13376
rect 1578 13336 1584 13348
rect 1636 13336 1642 13388
rect 3418 13376 3424 13388
rect 3379 13348 3424 13376
rect 3418 13336 3424 13348
rect 3476 13336 3482 13388
rect 20364 13385 20392 13416
rect 20349 13379 20407 13385
rect 20349 13345 20361 13379
rect 20395 13345 20407 13379
rect 20349 13339 20407 13345
rect 20533 13379 20591 13385
rect 20533 13345 20545 13379
rect 20579 13376 20591 13379
rect 20622 13376 20628 13388
rect 20579 13348 20628 13376
rect 20579 13345 20591 13348
rect 20533 13339 20591 13345
rect 20622 13336 20628 13348
rect 20680 13376 20686 13388
rect 21637 13379 21695 13385
rect 21637 13376 21649 13379
rect 20680 13348 21649 13376
rect 20680 13336 20686 13348
rect 21637 13345 21649 13348
rect 21683 13345 21695 13379
rect 22465 13379 22523 13385
rect 22465 13376 22477 13379
rect 21637 13339 21695 13345
rect 22066 13348 22477 13376
rect 17034 13268 17040 13320
rect 17092 13308 17098 13320
rect 17957 13311 18015 13317
rect 17957 13308 17969 13311
rect 17092 13280 17969 13308
rect 17092 13268 17098 13280
rect 17957 13277 17969 13280
rect 18003 13308 18015 13311
rect 18138 13308 18144 13320
rect 18003 13280 18144 13308
rect 18003 13277 18015 13280
rect 17957 13271 18015 13277
rect 18138 13268 18144 13280
rect 18196 13268 18202 13320
rect 18233 13311 18291 13317
rect 18233 13277 18245 13311
rect 18279 13277 18291 13311
rect 18233 13271 18291 13277
rect 1946 13200 1952 13252
rect 2004 13240 2010 13252
rect 3237 13243 3295 13249
rect 3237 13240 3249 13243
rect 2004 13212 3249 13240
rect 2004 13200 2010 13212
rect 3237 13209 3249 13212
rect 3283 13209 3295 13243
rect 18248 13240 18276 13271
rect 18322 13268 18328 13320
rect 18380 13308 18386 13320
rect 18966 13308 18972 13320
rect 18380 13280 18972 13308
rect 18380 13268 18386 13280
rect 18966 13268 18972 13280
rect 19024 13268 19030 13320
rect 20257 13311 20315 13317
rect 20257 13277 20269 13311
rect 20303 13308 20315 13311
rect 20806 13308 20812 13320
rect 20303 13280 20812 13308
rect 20303 13277 20315 13280
rect 20257 13271 20315 13277
rect 20806 13268 20812 13280
rect 20864 13268 20870 13320
rect 21450 13308 21456 13320
rect 21411 13280 21456 13308
rect 21450 13268 21456 13280
rect 21508 13268 21514 13320
rect 21545 13311 21603 13317
rect 21545 13277 21557 13311
rect 21591 13308 21603 13311
rect 22066 13308 22094 13348
rect 22465 13345 22477 13348
rect 22511 13376 22523 13379
rect 23014 13376 23020 13388
rect 22511 13348 23020 13376
rect 22511 13345 22523 13348
rect 22465 13339 22523 13345
rect 23014 13336 23020 13348
rect 23072 13336 23078 13388
rect 23492 13385 23520 13416
rect 23658 13404 23664 13416
rect 23716 13404 23722 13456
rect 23768 13385 23796 13484
rect 24578 13472 24584 13484
rect 24636 13472 24642 13524
rect 24670 13472 24676 13524
rect 24728 13512 24734 13524
rect 24765 13515 24823 13521
rect 24765 13512 24777 13515
rect 24728 13484 24777 13512
rect 24728 13472 24734 13484
rect 24765 13481 24777 13484
rect 24811 13481 24823 13515
rect 25590 13512 25596 13524
rect 25551 13484 25596 13512
rect 24765 13475 24823 13481
rect 25590 13472 25596 13484
rect 25648 13472 25654 13524
rect 23483 13379 23541 13385
rect 23483 13345 23495 13379
rect 23529 13345 23541 13379
rect 23483 13339 23541 13345
rect 23753 13379 23811 13385
rect 23753 13345 23765 13379
rect 23799 13345 23811 13379
rect 23753 13339 23811 13345
rect 21591 13280 22094 13308
rect 22557 13311 22615 13317
rect 21591 13277 21603 13280
rect 21545 13271 21603 13277
rect 22557 13277 22569 13311
rect 22603 13277 22615 13311
rect 22557 13271 22615 13277
rect 22925 13311 22983 13317
rect 22925 13277 22937 13311
rect 22971 13308 22983 13311
rect 23566 13308 23572 13320
rect 22971 13280 23428 13308
rect 23527 13280 23572 13308
rect 22971 13277 22983 13280
rect 22925 13271 22983 13277
rect 3237 13203 3295 13209
rect 17972 13212 18276 13240
rect 22572 13240 22600 13271
rect 23106 13240 23112 13252
rect 22572 13212 23112 13240
rect 17972 13184 18000 13212
rect 23106 13200 23112 13212
rect 23164 13200 23170 13252
rect 23400 13240 23428 13280
rect 23566 13268 23572 13280
rect 23624 13268 23630 13320
rect 23661 13311 23719 13317
rect 23661 13277 23673 13311
rect 23707 13308 23719 13311
rect 24026 13308 24032 13320
rect 23707 13280 24032 13308
rect 23707 13277 23719 13280
rect 23661 13271 23719 13277
rect 23474 13240 23480 13252
rect 23400 13212 23480 13240
rect 23474 13200 23480 13212
rect 23532 13200 23538 13252
rect 17954 13132 17960 13184
rect 18012 13132 18018 13184
rect 18509 13175 18567 13181
rect 18509 13141 18521 13175
rect 18555 13172 18567 13175
rect 18782 13172 18788 13184
rect 18555 13144 18788 13172
rect 18555 13141 18567 13144
rect 18509 13135 18567 13141
rect 18782 13132 18788 13144
rect 18840 13132 18846 13184
rect 21082 13172 21088 13184
rect 21043 13144 21088 13172
rect 21082 13132 21088 13144
rect 21140 13132 21146 13184
rect 22738 13172 22744 13184
rect 22699 13144 22744 13172
rect 22738 13132 22744 13144
rect 22796 13132 22802 13184
rect 22830 13132 22836 13184
rect 22888 13172 22894 13184
rect 23676 13172 23704 13271
rect 24026 13268 24032 13280
rect 24084 13268 24090 13320
rect 25777 13311 25835 13317
rect 25777 13277 25789 13311
rect 25823 13308 25835 13311
rect 25866 13308 25872 13320
rect 25823 13280 25872 13308
rect 25823 13277 25835 13280
rect 25777 13271 25835 13277
rect 25866 13268 25872 13280
rect 25924 13268 25930 13320
rect 25958 13268 25964 13320
rect 26016 13308 26022 13320
rect 26016 13280 26109 13308
rect 26016 13268 26022 13280
rect 24946 13240 24952 13252
rect 24907 13212 24952 13240
rect 24946 13200 24952 13212
rect 25004 13240 25010 13252
rect 25976 13240 26004 13268
rect 25004 13212 26004 13240
rect 25004 13200 25010 13212
rect 22888 13144 23704 13172
rect 23937 13175 23995 13181
rect 22888 13132 22894 13144
rect 23937 13141 23949 13175
rect 23983 13172 23995 13175
rect 24739 13175 24797 13181
rect 24739 13172 24751 13175
rect 23983 13144 24751 13172
rect 23983 13141 23995 13144
rect 23937 13135 23995 13141
rect 24739 13141 24751 13144
rect 24785 13141 24797 13175
rect 24739 13135 24797 13141
rect 1104 13082 29048 13104
rect 1104 13030 7896 13082
rect 7948 13030 7960 13082
rect 8012 13030 8024 13082
rect 8076 13030 8088 13082
rect 8140 13030 8152 13082
rect 8204 13030 14842 13082
rect 14894 13030 14906 13082
rect 14958 13030 14970 13082
rect 15022 13030 15034 13082
rect 15086 13030 15098 13082
rect 15150 13030 21788 13082
rect 21840 13030 21852 13082
rect 21904 13030 21916 13082
rect 21968 13030 21980 13082
rect 22032 13030 22044 13082
rect 22096 13030 28734 13082
rect 28786 13030 28798 13082
rect 28850 13030 28862 13082
rect 28914 13030 28926 13082
rect 28978 13030 28990 13082
rect 29042 13030 29048 13082
rect 1104 13008 29048 13030
rect 1946 12968 1952 12980
rect 1907 12940 1952 12968
rect 1946 12928 1952 12940
rect 2004 12928 2010 12980
rect 20438 12928 20444 12980
rect 20496 12968 20502 12980
rect 20533 12971 20591 12977
rect 20533 12968 20545 12971
rect 20496 12940 20545 12968
rect 20496 12928 20502 12940
rect 20533 12937 20545 12940
rect 20579 12937 20591 12971
rect 20533 12931 20591 12937
rect 22373 12971 22431 12977
rect 22373 12937 22385 12971
rect 22419 12968 22431 12971
rect 22462 12968 22468 12980
rect 22419 12940 22468 12968
rect 22419 12937 22431 12940
rect 22373 12931 22431 12937
rect 22462 12928 22468 12940
rect 22520 12928 22526 12980
rect 23750 12968 23756 12980
rect 22572 12940 23756 12968
rect 2038 12832 2044 12844
rect 1951 12804 2044 12832
rect 2038 12792 2044 12804
rect 2096 12832 2102 12844
rect 4982 12832 4988 12844
rect 2096 12804 4988 12832
rect 2096 12792 2102 12804
rect 4982 12792 4988 12804
rect 5040 12792 5046 12844
rect 16666 12792 16672 12844
rect 16724 12832 16730 12844
rect 16853 12835 16911 12841
rect 16853 12832 16865 12835
rect 16724 12804 16865 12832
rect 16724 12792 16730 12804
rect 16853 12801 16865 12804
rect 16899 12801 16911 12835
rect 16853 12795 16911 12801
rect 18046 12792 18052 12844
rect 18104 12832 18110 12844
rect 18693 12835 18751 12841
rect 18693 12832 18705 12835
rect 18104 12804 18705 12832
rect 18104 12792 18110 12804
rect 18693 12801 18705 12804
rect 18739 12801 18751 12835
rect 18693 12795 18751 12801
rect 18874 12792 18880 12844
rect 18932 12832 18938 12844
rect 19153 12835 19211 12841
rect 19153 12832 19165 12835
rect 18932 12804 19165 12832
rect 18932 12792 18938 12804
rect 19153 12801 19165 12804
rect 19199 12801 19211 12835
rect 19153 12795 19211 12801
rect 19886 12792 19892 12844
rect 19944 12832 19950 12844
rect 20162 12832 20168 12844
rect 19944 12804 20168 12832
rect 19944 12792 19950 12804
rect 20162 12792 20168 12804
rect 20220 12792 20226 12844
rect 20349 12835 20407 12841
rect 20349 12801 20361 12835
rect 20395 12832 20407 12835
rect 21082 12832 21088 12844
rect 20395 12804 21088 12832
rect 20395 12801 20407 12804
rect 20349 12795 20407 12801
rect 21082 12792 21088 12804
rect 21140 12792 21146 12844
rect 22572 12841 22600 12940
rect 23750 12928 23756 12940
rect 23808 12928 23814 12980
rect 25866 12968 25872 12980
rect 25827 12940 25872 12968
rect 25866 12928 25872 12940
rect 25924 12928 25930 12980
rect 26234 12968 26240 12980
rect 26195 12940 26240 12968
rect 26234 12928 26240 12940
rect 26292 12928 26298 12980
rect 23290 12860 23296 12912
rect 23348 12900 23354 12912
rect 23385 12903 23443 12909
rect 23385 12900 23397 12903
rect 23348 12872 23397 12900
rect 23348 12860 23354 12872
rect 23385 12869 23397 12872
rect 23431 12869 23443 12903
rect 23385 12863 23443 12869
rect 23569 12903 23627 12909
rect 23569 12869 23581 12903
rect 23615 12900 23627 12903
rect 23934 12900 23940 12912
rect 23615 12872 23940 12900
rect 23615 12869 23627 12872
rect 23569 12863 23627 12869
rect 23934 12860 23940 12872
rect 23992 12860 23998 12912
rect 22557 12835 22615 12841
rect 22557 12801 22569 12835
rect 22603 12801 22615 12835
rect 22557 12795 22615 12801
rect 22649 12835 22707 12841
rect 22649 12801 22661 12835
rect 22695 12832 22707 12835
rect 23474 12832 23480 12844
rect 22695 12804 23480 12832
rect 22695 12801 22707 12804
rect 22649 12795 22707 12801
rect 23474 12792 23480 12804
rect 23532 12792 23538 12844
rect 26329 12835 26387 12841
rect 26329 12801 26341 12835
rect 26375 12832 26387 12835
rect 26970 12832 26976 12844
rect 26375 12804 26976 12832
rect 26375 12801 26387 12804
rect 26329 12795 26387 12801
rect 26970 12792 26976 12804
rect 27028 12792 27034 12844
rect 27433 12835 27491 12841
rect 27433 12801 27445 12835
rect 27479 12832 27491 12835
rect 27614 12832 27620 12844
rect 27479 12804 27620 12832
rect 27479 12801 27491 12804
rect 27433 12795 27491 12801
rect 27614 12792 27620 12804
rect 27672 12792 27678 12844
rect 16942 12724 16948 12776
rect 17000 12764 17006 12776
rect 17129 12767 17187 12773
rect 17129 12764 17141 12767
rect 17000 12736 17141 12764
rect 17000 12724 17006 12736
rect 17129 12733 17141 12736
rect 17175 12733 17187 12767
rect 22738 12764 22744 12776
rect 22699 12736 22744 12764
rect 17129 12727 17187 12733
rect 17144 12696 17172 12727
rect 22738 12724 22744 12736
rect 22796 12724 22802 12776
rect 22833 12767 22891 12773
rect 22833 12733 22845 12767
rect 22879 12764 22891 12767
rect 23842 12764 23848 12776
rect 22879 12736 23848 12764
rect 22879 12733 22891 12736
rect 22833 12727 22891 12733
rect 23842 12724 23848 12736
rect 23900 12724 23906 12776
rect 26421 12767 26479 12773
rect 26421 12733 26433 12767
rect 26467 12764 26479 12767
rect 27338 12764 27344 12776
rect 26467 12736 27344 12764
rect 26467 12733 26479 12736
rect 26421 12727 26479 12733
rect 17494 12696 17500 12708
rect 17144 12668 17500 12696
rect 17494 12656 17500 12668
rect 17552 12696 17558 12708
rect 26436 12696 26464 12727
rect 27338 12724 27344 12736
rect 27396 12724 27402 12776
rect 17552 12668 26464 12696
rect 17552 12656 17558 12668
rect 26510 12656 26516 12708
rect 26568 12696 26574 12708
rect 27893 12699 27951 12705
rect 27893 12696 27905 12699
rect 26568 12668 27905 12696
rect 26568 12656 26574 12668
rect 27893 12665 27905 12668
rect 27939 12665 27951 12699
rect 27893 12659 27951 12665
rect 18230 12628 18236 12640
rect 18191 12600 18236 12628
rect 18230 12588 18236 12600
rect 18288 12588 18294 12640
rect 18601 12631 18659 12637
rect 18601 12597 18613 12631
rect 18647 12628 18659 12631
rect 18690 12628 18696 12640
rect 18647 12600 18696 12628
rect 18647 12597 18659 12600
rect 18601 12591 18659 12597
rect 18690 12588 18696 12600
rect 18748 12588 18754 12640
rect 19245 12631 19303 12637
rect 19245 12597 19257 12631
rect 19291 12628 19303 12631
rect 20254 12628 20260 12640
rect 19291 12600 20260 12628
rect 19291 12597 19303 12600
rect 19245 12591 19303 12597
rect 20254 12588 20260 12600
rect 20312 12588 20318 12640
rect 26694 12588 26700 12640
rect 26752 12628 26758 12640
rect 27341 12631 27399 12637
rect 27341 12628 27353 12631
rect 26752 12600 27353 12628
rect 26752 12588 26758 12600
rect 27341 12597 27353 12600
rect 27387 12597 27399 12631
rect 27341 12591 27399 12597
rect 1104 12538 28888 12560
rect 1104 12486 4423 12538
rect 4475 12486 4487 12538
rect 4539 12486 4551 12538
rect 4603 12486 4615 12538
rect 4667 12486 4679 12538
rect 4731 12486 11369 12538
rect 11421 12486 11433 12538
rect 11485 12486 11497 12538
rect 11549 12486 11561 12538
rect 11613 12486 11625 12538
rect 11677 12486 18315 12538
rect 18367 12486 18379 12538
rect 18431 12486 18443 12538
rect 18495 12486 18507 12538
rect 18559 12486 18571 12538
rect 18623 12486 25261 12538
rect 25313 12486 25325 12538
rect 25377 12486 25389 12538
rect 25441 12486 25453 12538
rect 25505 12486 25517 12538
rect 25569 12486 28888 12538
rect 1104 12464 28888 12486
rect 3510 12384 3516 12436
rect 3568 12424 3574 12436
rect 11054 12424 11060 12436
rect 3568 12396 11060 12424
rect 3568 12384 3574 12396
rect 11054 12384 11060 12396
rect 11112 12384 11118 12436
rect 17126 12384 17132 12436
rect 17184 12424 17190 12436
rect 17313 12427 17371 12433
rect 17313 12424 17325 12427
rect 17184 12396 17325 12424
rect 17184 12384 17190 12396
rect 17313 12393 17325 12396
rect 17359 12393 17371 12427
rect 17313 12387 17371 12393
rect 21542 12384 21548 12436
rect 21600 12424 21606 12436
rect 21821 12427 21879 12433
rect 21821 12424 21833 12427
rect 21600 12396 21833 12424
rect 21600 12384 21606 12396
rect 21821 12393 21833 12396
rect 21867 12393 21879 12427
rect 21821 12387 21879 12393
rect 21085 12359 21143 12365
rect 21085 12325 21097 12359
rect 21131 12325 21143 12359
rect 21085 12319 21143 12325
rect 16485 12291 16543 12297
rect 16485 12257 16497 12291
rect 16531 12288 16543 12291
rect 20162 12288 20168 12300
rect 16531 12260 20168 12288
rect 16531 12257 16543 12260
rect 16485 12251 16543 12257
rect 20162 12248 20168 12260
rect 20220 12288 20226 12300
rect 21100 12288 21128 12319
rect 24946 12288 24952 12300
rect 20220 12260 21128 12288
rect 21284 12260 24952 12288
rect 20220 12248 20226 12260
rect 1670 12220 1676 12232
rect 1631 12192 1676 12220
rect 1670 12180 1676 12192
rect 1728 12180 1734 12232
rect 16666 12220 16672 12232
rect 16627 12192 16672 12220
rect 16666 12180 16672 12192
rect 16724 12180 16730 12232
rect 21284 12229 21312 12260
rect 24946 12248 24952 12260
rect 25004 12248 25010 12300
rect 26510 12288 26516 12300
rect 26471 12260 26516 12288
rect 26510 12248 26516 12260
rect 26568 12248 26574 12300
rect 26694 12288 26700 12300
rect 26655 12260 26700 12288
rect 26694 12248 26700 12260
rect 26752 12248 26758 12300
rect 28350 12288 28356 12300
rect 28311 12260 28356 12288
rect 28350 12248 28356 12260
rect 28408 12248 28414 12300
rect 16853 12223 16911 12229
rect 16853 12189 16865 12223
rect 16899 12220 16911 12223
rect 17497 12223 17555 12229
rect 17497 12220 17509 12223
rect 16899 12192 17509 12220
rect 16899 12189 16911 12192
rect 16853 12183 16911 12189
rect 17497 12189 17509 12192
rect 17543 12189 17555 12223
rect 17497 12183 17555 12189
rect 21269 12223 21327 12229
rect 21269 12189 21281 12223
rect 21315 12189 21327 12223
rect 21269 12183 21327 12189
rect 21634 12180 21640 12232
rect 21692 12220 21698 12232
rect 22005 12223 22063 12229
rect 22005 12220 22017 12223
rect 21692 12192 22017 12220
rect 21692 12180 21698 12192
rect 22005 12189 22017 12192
rect 22051 12189 22063 12223
rect 22005 12183 22063 12189
rect 1104 11994 29048 12016
rect 1104 11942 7896 11994
rect 7948 11942 7960 11994
rect 8012 11942 8024 11994
rect 8076 11942 8088 11994
rect 8140 11942 8152 11994
rect 8204 11942 14842 11994
rect 14894 11942 14906 11994
rect 14958 11942 14970 11994
rect 15022 11942 15034 11994
rect 15086 11942 15098 11994
rect 15150 11942 21788 11994
rect 21840 11942 21852 11994
rect 21904 11942 21916 11994
rect 21968 11942 21980 11994
rect 22032 11942 22044 11994
rect 22096 11942 28734 11994
rect 28786 11942 28798 11994
rect 28850 11942 28862 11994
rect 28914 11942 28926 11994
rect 28978 11942 28990 11994
rect 29042 11942 29048 11994
rect 1104 11920 29048 11942
rect 16666 11840 16672 11892
rect 16724 11880 16730 11892
rect 16853 11883 16911 11889
rect 16853 11880 16865 11883
rect 16724 11852 16865 11880
rect 16724 11840 16730 11852
rect 16853 11849 16865 11852
rect 16899 11849 16911 11883
rect 16853 11843 16911 11849
rect 18785 11883 18843 11889
rect 18785 11849 18797 11883
rect 18831 11880 18843 11883
rect 18874 11880 18880 11892
rect 18831 11852 18880 11880
rect 18831 11849 18843 11852
rect 18785 11843 18843 11849
rect 18874 11840 18880 11852
rect 18932 11840 18938 11892
rect 18230 11812 18236 11824
rect 18191 11784 18236 11812
rect 18230 11772 18236 11784
rect 18288 11772 18294 11824
rect 1670 11744 1676 11756
rect 1631 11716 1676 11744
rect 1670 11704 1676 11716
rect 1728 11704 1734 11756
rect 17218 11744 17224 11756
rect 17179 11716 17224 11744
rect 17218 11704 17224 11716
rect 17276 11704 17282 11756
rect 17313 11747 17371 11753
rect 17313 11713 17325 11747
rect 17359 11744 17371 11747
rect 18046 11744 18052 11756
rect 17359 11716 18052 11744
rect 17359 11713 17371 11716
rect 17313 11707 17371 11713
rect 18046 11704 18052 11716
rect 18104 11704 18110 11756
rect 18782 11744 18788 11756
rect 18743 11716 18788 11744
rect 18782 11704 18788 11716
rect 18840 11704 18846 11756
rect 27062 11704 27068 11756
rect 27120 11744 27126 11756
rect 27157 11747 27215 11753
rect 27157 11744 27169 11747
rect 27120 11716 27169 11744
rect 27120 11704 27126 11716
rect 27157 11713 27169 11716
rect 27203 11713 27215 11747
rect 27157 11707 27215 11713
rect 1854 11676 1860 11688
rect 1815 11648 1860 11676
rect 1854 11636 1860 11648
rect 1912 11636 1918 11688
rect 2774 11676 2780 11688
rect 2735 11648 2780 11676
rect 2774 11636 2780 11648
rect 2832 11636 2838 11688
rect 17494 11676 17500 11688
rect 17455 11648 17500 11676
rect 17494 11636 17500 11648
rect 17552 11636 17558 11688
rect 18874 11676 18880 11688
rect 18835 11648 18880 11676
rect 18874 11636 18880 11648
rect 18932 11636 18938 11688
rect 26694 11500 26700 11552
rect 26752 11540 26758 11552
rect 27249 11543 27307 11549
rect 27249 11540 27261 11543
rect 26752 11512 27261 11540
rect 26752 11500 26758 11512
rect 27249 11509 27261 11512
rect 27295 11509 27307 11543
rect 27249 11503 27307 11509
rect 1104 11450 28888 11472
rect 1104 11398 4423 11450
rect 4475 11398 4487 11450
rect 4539 11398 4551 11450
rect 4603 11398 4615 11450
rect 4667 11398 4679 11450
rect 4731 11398 11369 11450
rect 11421 11398 11433 11450
rect 11485 11398 11497 11450
rect 11549 11398 11561 11450
rect 11613 11398 11625 11450
rect 11677 11398 18315 11450
rect 18367 11398 18379 11450
rect 18431 11398 18443 11450
rect 18495 11398 18507 11450
rect 18559 11398 18571 11450
rect 18623 11398 25261 11450
rect 25313 11398 25325 11450
rect 25377 11398 25389 11450
rect 25441 11398 25453 11450
rect 25505 11398 25517 11450
rect 25569 11398 28888 11450
rect 1104 11376 28888 11398
rect 1854 11336 1860 11348
rect 1815 11308 1860 11336
rect 1854 11296 1860 11308
rect 1912 11296 1918 11348
rect 18693 11339 18751 11345
rect 18693 11305 18705 11339
rect 18739 11336 18751 11339
rect 18782 11336 18788 11348
rect 18739 11308 18788 11336
rect 18739 11305 18751 11308
rect 18693 11299 18751 11305
rect 18782 11296 18788 11308
rect 18840 11296 18846 11348
rect 18877 11339 18935 11345
rect 18877 11305 18889 11339
rect 18923 11336 18935 11339
rect 19150 11336 19156 11348
rect 18923 11308 19156 11336
rect 18923 11305 18935 11308
rect 18877 11299 18935 11305
rect 19150 11296 19156 11308
rect 19208 11296 19214 11348
rect 4338 11200 4344 11212
rect 4299 11172 4344 11200
rect 4338 11160 4344 11172
rect 4396 11160 4402 11212
rect 26694 11200 26700 11212
rect 26655 11172 26700 11200
rect 26694 11160 26700 11172
rect 26752 11160 26758 11212
rect 1486 11092 1492 11144
rect 1544 11132 1550 11144
rect 1765 11135 1823 11141
rect 1765 11132 1777 11135
rect 1544 11104 1777 11132
rect 1544 11092 1550 11104
rect 1765 11101 1777 11104
rect 1811 11101 1823 11135
rect 1765 11095 1823 11101
rect 2958 11092 2964 11144
rect 3016 11132 3022 11144
rect 3973 11135 4031 11141
rect 3973 11132 3985 11135
rect 3016 11104 3985 11132
rect 3016 11092 3022 11104
rect 3973 11101 3985 11104
rect 4019 11101 4031 11135
rect 17678 11132 17684 11144
rect 17639 11104 17684 11132
rect 3973 11095 4031 11101
rect 17678 11092 17684 11104
rect 17736 11092 17742 11144
rect 26510 11132 26516 11144
rect 26471 11104 26516 11132
rect 26510 11092 26516 11104
rect 26568 11092 26574 11144
rect 18322 11024 18328 11076
rect 18380 11064 18386 11076
rect 18509 11067 18567 11073
rect 18509 11064 18521 11067
rect 18380 11036 18521 11064
rect 18380 11024 18386 11036
rect 18509 11033 18521 11036
rect 18555 11033 18567 11067
rect 18509 11027 18567 11033
rect 28353 11067 28411 11073
rect 28353 11033 28365 11067
rect 28399 11064 28411 11067
rect 29914 11064 29920 11076
rect 28399 11036 29920 11064
rect 28399 11033 28411 11036
rect 28353 11027 28411 11033
rect 29914 11024 29920 11036
rect 29972 11024 29978 11076
rect 17770 10996 17776 11008
rect 17731 10968 17776 10996
rect 17770 10956 17776 10968
rect 17828 10956 17834 11008
rect 18719 10999 18777 11005
rect 18719 10965 18731 10999
rect 18765 10996 18777 10999
rect 19242 10996 19248 11008
rect 18765 10968 19248 10996
rect 18765 10965 18777 10968
rect 18719 10959 18777 10965
rect 19242 10956 19248 10968
rect 19300 10956 19306 11008
rect 1104 10906 29048 10928
rect 1104 10854 7896 10906
rect 7948 10854 7960 10906
rect 8012 10854 8024 10906
rect 8076 10854 8088 10906
rect 8140 10854 8152 10906
rect 8204 10854 14842 10906
rect 14894 10854 14906 10906
rect 14958 10854 14970 10906
rect 15022 10854 15034 10906
rect 15086 10854 15098 10906
rect 15150 10854 21788 10906
rect 21840 10854 21852 10906
rect 21904 10854 21916 10906
rect 21968 10854 21980 10906
rect 22032 10854 22044 10906
rect 22096 10854 28734 10906
rect 28786 10854 28798 10906
rect 28850 10854 28862 10906
rect 28914 10854 28926 10906
rect 28978 10854 28990 10906
rect 29042 10854 29048 10906
rect 1104 10832 29048 10854
rect 18230 10792 18236 10804
rect 18191 10764 18236 10792
rect 18230 10752 18236 10764
rect 18288 10752 18294 10804
rect 18693 10795 18751 10801
rect 18693 10761 18705 10795
rect 18739 10792 18751 10795
rect 18874 10792 18880 10804
rect 18739 10764 18880 10792
rect 18739 10761 18751 10764
rect 18693 10755 18751 10761
rect 18874 10752 18880 10764
rect 18932 10752 18938 10804
rect 17770 10684 17776 10736
rect 17828 10724 17834 10736
rect 17828 10696 20024 10724
rect 17828 10684 17834 10696
rect 17880 10665 17908 10696
rect 17865 10659 17923 10665
rect 17865 10625 17877 10659
rect 17911 10625 17923 10659
rect 18874 10656 18880 10668
rect 18835 10628 18880 10656
rect 17865 10619 17923 10625
rect 18874 10616 18880 10628
rect 18932 10616 18938 10668
rect 18969 10659 19027 10665
rect 18969 10625 18981 10659
rect 19015 10625 19027 10659
rect 19150 10656 19156 10668
rect 19111 10628 19156 10656
rect 18969 10619 19027 10625
rect 17218 10548 17224 10600
rect 17276 10588 17282 10600
rect 17773 10591 17831 10597
rect 17773 10588 17785 10591
rect 17276 10560 17785 10588
rect 17276 10548 17282 10560
rect 17773 10557 17785 10560
rect 17819 10557 17831 10591
rect 17773 10551 17831 10557
rect 17788 10520 17816 10551
rect 17954 10548 17960 10600
rect 18012 10588 18018 10600
rect 18984 10588 19012 10619
rect 19150 10616 19156 10628
rect 19208 10616 19214 10668
rect 19242 10616 19248 10668
rect 19300 10656 19306 10668
rect 19996 10665 20024 10696
rect 19705 10659 19763 10665
rect 19705 10656 19717 10659
rect 19300 10628 19717 10656
rect 19300 10616 19306 10628
rect 19705 10625 19717 10628
rect 19751 10625 19763 10659
rect 19705 10619 19763 10625
rect 19889 10659 19947 10665
rect 19889 10625 19901 10659
rect 19935 10625 19947 10659
rect 19889 10619 19947 10625
rect 19981 10659 20039 10665
rect 19981 10625 19993 10659
rect 20027 10625 20039 10659
rect 20254 10656 20260 10668
rect 20215 10628 20260 10656
rect 19981 10619 20039 10625
rect 18012 10560 19012 10588
rect 18012 10548 18018 10560
rect 19904 10520 19932 10619
rect 20254 10616 20260 10628
rect 20312 10616 20318 10668
rect 26510 10616 26516 10668
rect 26568 10656 26574 10668
rect 27157 10659 27215 10665
rect 27157 10656 27169 10659
rect 26568 10628 27169 10656
rect 26568 10616 26574 10628
rect 27157 10625 27169 10628
rect 27203 10625 27215 10659
rect 27157 10619 27215 10625
rect 20162 10588 20168 10600
rect 20075 10560 20168 10588
rect 20162 10548 20168 10560
rect 20220 10588 20226 10600
rect 27430 10588 27436 10600
rect 20220 10560 27436 10588
rect 20220 10548 20226 10560
rect 27430 10548 27436 10560
rect 27488 10548 27494 10600
rect 17788 10492 19932 10520
rect 17589 10455 17647 10461
rect 17589 10421 17601 10455
rect 17635 10452 17647 10455
rect 18138 10452 18144 10464
rect 17635 10424 18144 10452
rect 17635 10421 17647 10424
rect 17589 10415 17647 10421
rect 18138 10412 18144 10424
rect 18196 10412 18202 10464
rect 27985 10455 28043 10461
rect 27985 10421 27997 10455
rect 28031 10452 28043 10455
rect 28350 10452 28356 10464
rect 28031 10424 28356 10452
rect 28031 10421 28043 10424
rect 27985 10415 28043 10421
rect 28350 10412 28356 10424
rect 28408 10412 28414 10464
rect 1104 10362 28888 10384
rect 1104 10310 4423 10362
rect 4475 10310 4487 10362
rect 4539 10310 4551 10362
rect 4603 10310 4615 10362
rect 4667 10310 4679 10362
rect 4731 10310 11369 10362
rect 11421 10310 11433 10362
rect 11485 10310 11497 10362
rect 11549 10310 11561 10362
rect 11613 10310 11625 10362
rect 11677 10310 18315 10362
rect 18367 10310 18379 10362
rect 18431 10310 18443 10362
rect 18495 10310 18507 10362
rect 18559 10310 18571 10362
rect 18623 10310 25261 10362
rect 25313 10310 25325 10362
rect 25377 10310 25389 10362
rect 25441 10310 25453 10362
rect 25505 10310 25517 10362
rect 25569 10310 28888 10362
rect 1104 10288 28888 10310
rect 18230 10248 18236 10260
rect 18191 10220 18236 10248
rect 18230 10208 18236 10220
rect 18288 10208 18294 10260
rect 18049 10183 18107 10189
rect 18049 10149 18061 10183
rect 18095 10180 18107 10183
rect 19150 10180 19156 10192
rect 18095 10152 19156 10180
rect 18095 10149 18107 10152
rect 18049 10143 18107 10149
rect 19150 10140 19156 10152
rect 19208 10180 19214 10192
rect 19429 10183 19487 10189
rect 19429 10180 19441 10183
rect 19208 10152 19441 10180
rect 19208 10140 19214 10152
rect 19429 10149 19441 10152
rect 19475 10149 19487 10183
rect 19429 10143 19487 10149
rect 18138 10112 18144 10124
rect 18099 10084 18144 10112
rect 18138 10072 18144 10084
rect 18196 10072 18202 10124
rect 19797 10115 19855 10121
rect 19797 10081 19809 10115
rect 19843 10112 19855 10115
rect 20254 10112 20260 10124
rect 19843 10084 20260 10112
rect 19843 10081 19855 10084
rect 19797 10075 19855 10081
rect 20254 10072 20260 10084
rect 20312 10072 20318 10124
rect 27522 10112 27528 10124
rect 27483 10084 27528 10112
rect 27522 10072 27528 10084
rect 27580 10072 27586 10124
rect 28350 10112 28356 10124
rect 28311 10084 28356 10112
rect 28350 10072 28356 10084
rect 28408 10072 28414 10124
rect 1670 10044 1676 10056
rect 1631 10016 1676 10044
rect 1670 10004 1676 10016
rect 1728 10004 1734 10056
rect 2958 10004 2964 10056
rect 3016 10044 3022 10056
rect 3053 10047 3111 10053
rect 3053 10044 3065 10047
rect 3016 10016 3065 10044
rect 3016 10004 3022 10016
rect 3053 10013 3065 10016
rect 3099 10013 3111 10047
rect 17954 10044 17960 10056
rect 17915 10016 17960 10044
rect 3053 10007 3111 10013
rect 17954 10004 17960 10016
rect 18012 10004 18018 10056
rect 19613 10047 19671 10053
rect 19613 10013 19625 10047
rect 19659 10044 19671 10047
rect 20162 10044 20168 10056
rect 19659 10016 20168 10044
rect 19659 10013 19671 10016
rect 19613 10007 19671 10013
rect 20162 10004 20168 10016
rect 20220 10004 20226 10056
rect 17773 9979 17831 9985
rect 17773 9945 17785 9979
rect 17819 9976 17831 9979
rect 18874 9976 18880 9988
rect 17819 9948 18880 9976
rect 17819 9945 17831 9948
rect 17773 9939 17831 9945
rect 18874 9936 18880 9948
rect 18932 9936 18938 9988
rect 28166 9976 28172 9988
rect 28127 9948 28172 9976
rect 28166 9936 28172 9948
rect 28224 9936 28230 9988
rect 2961 9911 3019 9917
rect 2961 9877 2973 9911
rect 3007 9908 3019 9911
rect 4062 9908 4068 9920
rect 3007 9880 4068 9908
rect 3007 9877 3019 9880
rect 2961 9871 3019 9877
rect 4062 9868 4068 9880
rect 4120 9868 4126 9920
rect 1104 9818 29048 9840
rect 1104 9766 7896 9818
rect 7948 9766 7960 9818
rect 8012 9766 8024 9818
rect 8076 9766 8088 9818
rect 8140 9766 8152 9818
rect 8204 9766 14842 9818
rect 14894 9766 14906 9818
rect 14958 9766 14970 9818
rect 15022 9766 15034 9818
rect 15086 9766 15098 9818
rect 15150 9766 21788 9818
rect 21840 9766 21852 9818
rect 21904 9766 21916 9818
rect 21968 9766 21980 9818
rect 22032 9766 22044 9818
rect 22096 9766 28734 9818
rect 28786 9766 28798 9818
rect 28850 9766 28862 9818
rect 28914 9766 28926 9818
rect 28978 9766 28990 9818
rect 29042 9766 29048 9818
rect 1104 9744 29048 9766
rect 27801 9707 27859 9713
rect 27801 9673 27813 9707
rect 27847 9704 27859 9707
rect 28166 9704 28172 9716
rect 27847 9676 28172 9704
rect 27847 9673 27859 9676
rect 27801 9667 27859 9673
rect 28166 9664 28172 9676
rect 28224 9664 28230 9716
rect 1670 9568 1676 9580
rect 1631 9540 1676 9568
rect 1670 9528 1676 9540
rect 1728 9528 1734 9580
rect 20441 9571 20499 9577
rect 20441 9537 20453 9571
rect 20487 9568 20499 9571
rect 20530 9568 20536 9580
rect 20487 9540 20536 9568
rect 20487 9537 20499 9540
rect 20441 9531 20499 9537
rect 20530 9528 20536 9540
rect 20588 9528 20594 9580
rect 27338 9528 27344 9580
rect 27396 9568 27402 9580
rect 27614 9568 27620 9580
rect 27396 9540 27620 9568
rect 27396 9528 27402 9540
rect 27614 9528 27620 9540
rect 27672 9568 27678 9580
rect 27709 9571 27767 9577
rect 27709 9568 27721 9571
rect 27672 9540 27721 9568
rect 27672 9528 27678 9540
rect 27709 9537 27721 9540
rect 27755 9537 27767 9571
rect 27709 9531 27767 9537
rect 1854 9500 1860 9512
rect 1815 9472 1860 9500
rect 1854 9460 1860 9472
rect 1912 9460 1918 9512
rect 2774 9500 2780 9512
rect 2735 9472 2780 9500
rect 2774 9460 2780 9472
rect 2832 9460 2838 9512
rect 4157 9367 4215 9373
rect 4157 9333 4169 9367
rect 4203 9364 4215 9367
rect 4246 9364 4252 9376
rect 4203 9336 4252 9364
rect 4203 9333 4215 9336
rect 4157 9327 4215 9333
rect 4246 9324 4252 9336
rect 4304 9324 4310 9376
rect 20533 9367 20591 9373
rect 20533 9333 20545 9367
rect 20579 9364 20591 9367
rect 20622 9364 20628 9376
rect 20579 9336 20628 9364
rect 20579 9333 20591 9336
rect 20533 9327 20591 9333
rect 20622 9324 20628 9336
rect 20680 9324 20686 9376
rect 1104 9274 28888 9296
rect 1104 9222 4423 9274
rect 4475 9222 4487 9274
rect 4539 9222 4551 9274
rect 4603 9222 4615 9274
rect 4667 9222 4679 9274
rect 4731 9222 11369 9274
rect 11421 9222 11433 9274
rect 11485 9222 11497 9274
rect 11549 9222 11561 9274
rect 11613 9222 11625 9274
rect 11677 9222 18315 9274
rect 18367 9222 18379 9274
rect 18431 9222 18443 9274
rect 18495 9222 18507 9274
rect 18559 9222 18571 9274
rect 18623 9222 25261 9274
rect 25313 9222 25325 9274
rect 25377 9222 25389 9274
rect 25441 9222 25453 9274
rect 25505 9222 25517 9274
rect 25569 9222 28888 9274
rect 1104 9200 28888 9222
rect 2958 9024 2964 9036
rect 2919 8996 2964 9024
rect 2958 8984 2964 8996
rect 3016 8984 3022 9036
rect 1578 8956 1584 8968
rect 1539 8928 1584 8956
rect 1578 8916 1584 8928
rect 1636 8916 1642 8968
rect 26510 8956 26516 8968
rect 26471 8928 26516 8956
rect 26510 8916 26516 8928
rect 26568 8916 26574 8968
rect 28350 8956 28356 8968
rect 28311 8928 28356 8956
rect 28350 8916 28356 8928
rect 28408 8916 28414 8968
rect 1762 8888 1768 8900
rect 1723 8860 1768 8888
rect 1762 8848 1768 8860
rect 1820 8848 1826 8900
rect 26697 8891 26755 8897
rect 26697 8857 26709 8891
rect 26743 8888 26755 8891
rect 27246 8888 27252 8900
rect 26743 8860 27252 8888
rect 26743 8857 26755 8860
rect 26697 8851 26755 8857
rect 27246 8848 27252 8860
rect 27304 8848 27310 8900
rect 1104 8730 29048 8752
rect 1104 8678 7896 8730
rect 7948 8678 7960 8730
rect 8012 8678 8024 8730
rect 8076 8678 8088 8730
rect 8140 8678 8152 8730
rect 8204 8678 14842 8730
rect 14894 8678 14906 8730
rect 14958 8678 14970 8730
rect 15022 8678 15034 8730
rect 15086 8678 15098 8730
rect 15150 8678 21788 8730
rect 21840 8678 21852 8730
rect 21904 8678 21916 8730
rect 21968 8678 21980 8730
rect 22032 8678 22044 8730
rect 22096 8678 28734 8730
rect 28786 8678 28798 8730
rect 28850 8678 28862 8730
rect 28914 8678 28926 8730
rect 28978 8678 28990 8730
rect 29042 8678 29048 8730
rect 1104 8656 29048 8678
rect 1854 8616 1860 8628
rect 1815 8588 1860 8616
rect 1854 8576 1860 8588
rect 1912 8576 1918 8628
rect 4338 8616 4344 8628
rect 2792 8588 4344 8616
rect 1949 8483 2007 8489
rect 1949 8449 1961 8483
rect 1995 8480 2007 8483
rect 2792 8480 2820 8588
rect 4338 8576 4344 8588
rect 4396 8616 4402 8628
rect 27246 8616 27252 8628
rect 4396 8588 6914 8616
rect 27207 8588 27252 8616
rect 4396 8576 4402 8588
rect 4062 8548 4068 8560
rect 4023 8520 4068 8548
rect 4062 8508 4068 8520
rect 4120 8508 4126 8560
rect 1995 8452 2820 8480
rect 1995 8449 2007 8452
rect 1949 8443 2007 8449
rect 4246 8440 4252 8492
rect 4304 8480 4310 8492
rect 6886 8480 6914 8588
rect 27246 8576 27252 8588
rect 27304 8576 27310 8628
rect 26510 8508 26516 8560
rect 26568 8548 26574 8560
rect 26568 8520 27844 8548
rect 26568 8508 26574 8520
rect 27816 8489 27844 8520
rect 27341 8483 27399 8489
rect 27341 8480 27353 8483
rect 4304 8452 4349 8480
rect 6886 8452 27353 8480
rect 4304 8440 4310 8452
rect 27341 8449 27353 8452
rect 27387 8449 27399 8483
rect 27341 8443 27399 8449
rect 27801 8483 27859 8489
rect 27801 8449 27813 8483
rect 27847 8449 27859 8483
rect 27801 8443 27859 8449
rect 3326 8412 3332 8424
rect 3287 8384 3332 8412
rect 3326 8372 3332 8384
rect 3384 8372 3390 8424
rect 27356 8412 27384 8443
rect 27356 8384 27844 8412
rect 27816 8356 27844 8384
rect 27798 8304 27804 8356
rect 27856 8304 27862 8356
rect 26602 8276 26608 8288
rect 26563 8248 26608 8276
rect 26602 8236 26608 8248
rect 26660 8236 26666 8288
rect 1104 8186 28888 8208
rect 1104 8134 4423 8186
rect 4475 8134 4487 8186
rect 4539 8134 4551 8186
rect 4603 8134 4615 8186
rect 4667 8134 4679 8186
rect 4731 8134 11369 8186
rect 11421 8134 11433 8186
rect 11485 8134 11497 8186
rect 11549 8134 11561 8186
rect 11613 8134 11625 8186
rect 11677 8134 18315 8186
rect 18367 8134 18379 8186
rect 18431 8134 18443 8186
rect 18495 8134 18507 8186
rect 18559 8134 18571 8186
rect 18623 8134 25261 8186
rect 25313 8134 25325 8186
rect 25377 8134 25389 8186
rect 25441 8134 25453 8186
rect 25505 8134 25517 8186
rect 25569 8134 28888 8186
rect 1104 8112 28888 8134
rect 1578 8032 1584 8084
rect 1636 8072 1642 8084
rect 1673 8075 1731 8081
rect 1673 8072 1685 8075
rect 1636 8044 1685 8072
rect 1636 8032 1642 8044
rect 1673 8041 1685 8044
rect 1719 8041 1731 8075
rect 1673 8035 1731 8041
rect 1762 8032 1768 8084
rect 1820 8072 1826 8084
rect 2409 8075 2467 8081
rect 2409 8072 2421 8075
rect 1820 8044 2421 8072
rect 1820 8032 1826 8044
rect 2409 8041 2421 8044
rect 2455 8041 2467 8075
rect 2409 8035 2467 8041
rect 27706 7936 27712 7948
rect 26206 7908 27712 7936
rect 1486 7828 1492 7880
rect 1544 7868 1550 7880
rect 2498 7868 2504 7880
rect 1544 7840 2504 7868
rect 1544 7828 1550 7840
rect 2498 7828 2504 7840
rect 2556 7828 2562 7880
rect 3329 7871 3387 7877
rect 3329 7837 3341 7871
rect 3375 7837 3387 7871
rect 3329 7831 3387 7837
rect 3344 7800 3372 7831
rect 3878 7828 3884 7880
rect 3936 7868 3942 7880
rect 3973 7871 4031 7877
rect 3973 7868 3985 7871
rect 3936 7840 3985 7868
rect 3936 7828 3942 7840
rect 3973 7837 3985 7840
rect 4019 7837 4031 7871
rect 3973 7831 4031 7837
rect 25682 7828 25688 7880
rect 25740 7868 25746 7880
rect 25869 7871 25927 7877
rect 25869 7868 25881 7871
rect 25740 7840 25881 7868
rect 25740 7828 25746 7840
rect 25869 7837 25881 7840
rect 25915 7868 25927 7871
rect 26206 7868 26234 7908
rect 27706 7896 27712 7908
rect 27764 7896 27770 7948
rect 25915 7840 26234 7868
rect 26513 7871 26571 7877
rect 25915 7837 25927 7840
rect 25869 7831 25927 7837
rect 26513 7837 26525 7871
rect 26559 7837 26571 7871
rect 26513 7831 26571 7837
rect 4890 7800 4896 7812
rect 3344 7772 4896 7800
rect 4890 7760 4896 7772
rect 4948 7760 4954 7812
rect 4065 7735 4123 7741
rect 4065 7701 4077 7735
rect 4111 7732 4123 7735
rect 4706 7732 4712 7744
rect 4111 7704 4712 7732
rect 4111 7701 4123 7704
rect 4065 7695 4123 7701
rect 4706 7692 4712 7704
rect 4764 7692 4770 7744
rect 25961 7735 26019 7741
rect 25961 7701 25973 7735
rect 26007 7732 26019 7735
rect 26418 7732 26424 7744
rect 26007 7704 26424 7732
rect 26007 7701 26019 7704
rect 25961 7695 26019 7701
rect 26418 7692 26424 7704
rect 26476 7692 26482 7744
rect 26528 7732 26556 7831
rect 26694 7800 26700 7812
rect 26655 7772 26700 7800
rect 26694 7760 26700 7772
rect 26752 7760 26758 7812
rect 28353 7803 28411 7809
rect 28353 7769 28365 7803
rect 28399 7800 28411 7803
rect 29914 7800 29920 7812
rect 28399 7772 29920 7800
rect 28399 7769 28411 7772
rect 28353 7763 28411 7769
rect 29914 7760 29920 7772
rect 29972 7760 29978 7812
rect 27798 7732 27804 7744
rect 26528 7704 27804 7732
rect 27798 7692 27804 7704
rect 27856 7692 27862 7744
rect 1104 7642 29048 7664
rect 1104 7590 7896 7642
rect 7948 7590 7960 7642
rect 8012 7590 8024 7642
rect 8076 7590 8088 7642
rect 8140 7590 8152 7642
rect 8204 7590 14842 7642
rect 14894 7590 14906 7642
rect 14958 7590 14970 7642
rect 15022 7590 15034 7642
rect 15086 7590 15098 7642
rect 15150 7590 21788 7642
rect 21840 7590 21852 7642
rect 21904 7590 21916 7642
rect 21968 7590 21980 7642
rect 22032 7590 22044 7642
rect 22096 7590 28734 7642
rect 28786 7590 28798 7642
rect 28850 7590 28862 7642
rect 28914 7590 28926 7642
rect 28978 7590 28990 7642
rect 29042 7590 29048 7642
rect 1104 7568 29048 7590
rect 3050 7460 3056 7472
rect 3011 7432 3056 7460
rect 3050 7420 3056 7432
rect 3108 7420 3114 7472
rect 4706 7460 4712 7472
rect 4667 7432 4712 7460
rect 4706 7420 4712 7432
rect 4764 7420 4770 7472
rect 26418 7460 26424 7472
rect 26379 7432 26424 7460
rect 26418 7420 26424 7432
rect 26476 7420 26482 7472
rect 4890 7352 4896 7404
rect 4948 7392 4954 7404
rect 4948 7364 4993 7392
rect 4948 7352 4954 7364
rect 26602 7352 26608 7404
rect 26660 7392 26666 7404
rect 27798 7392 27804 7404
rect 26660 7364 26705 7392
rect 27759 7364 27804 7392
rect 26660 7352 26666 7364
rect 27798 7352 27804 7364
rect 27856 7352 27862 7404
rect 26142 7324 26148 7336
rect 26103 7296 26148 7324
rect 26142 7284 26148 7296
rect 26200 7284 26206 7336
rect 1670 7148 1676 7200
rect 1728 7188 1734 7200
rect 1765 7191 1823 7197
rect 1765 7188 1777 7191
rect 1728 7160 1777 7188
rect 1728 7148 1734 7160
rect 1765 7157 1777 7160
rect 1811 7157 1823 7191
rect 27154 7188 27160 7200
rect 27115 7160 27160 7188
rect 1765 7151 1823 7157
rect 27154 7148 27160 7160
rect 27212 7148 27218 7200
rect 1104 7098 28888 7120
rect 1104 7046 4423 7098
rect 4475 7046 4487 7098
rect 4539 7046 4551 7098
rect 4603 7046 4615 7098
rect 4667 7046 4679 7098
rect 4731 7046 11369 7098
rect 11421 7046 11433 7098
rect 11485 7046 11497 7098
rect 11549 7046 11561 7098
rect 11613 7046 11625 7098
rect 11677 7046 18315 7098
rect 18367 7046 18379 7098
rect 18431 7046 18443 7098
rect 18495 7046 18507 7098
rect 18559 7046 18571 7098
rect 18623 7046 25261 7098
rect 25313 7046 25325 7098
rect 25377 7046 25389 7098
rect 25441 7046 25453 7098
rect 25505 7046 25517 7098
rect 25569 7046 28888 7098
rect 1104 7024 28888 7046
rect 3970 6944 3976 6996
rect 4028 6984 4034 6996
rect 5350 6984 5356 6996
rect 4028 6956 5356 6984
rect 4028 6944 4034 6956
rect 5350 6944 5356 6956
rect 5408 6944 5414 6996
rect 7742 6876 7748 6928
rect 7800 6876 7806 6928
rect 3970 6848 3976 6860
rect 2424 6820 3976 6848
rect 1578 6780 1584 6792
rect 1539 6752 1584 6780
rect 1578 6740 1584 6752
rect 1636 6740 1642 6792
rect 2424 6789 2452 6820
rect 3970 6808 3976 6820
rect 4028 6808 4034 6860
rect 4062 6808 4068 6860
rect 4120 6848 4126 6860
rect 5445 6851 5503 6857
rect 4120 6820 4476 6848
rect 4120 6808 4126 6820
rect 2409 6783 2467 6789
rect 2409 6749 2421 6783
rect 2455 6749 2467 6783
rect 2866 6780 2872 6792
rect 2827 6752 2872 6780
rect 2409 6743 2467 6749
rect 2866 6740 2872 6752
rect 2924 6740 2930 6792
rect 4341 6783 4399 6789
rect 4341 6749 4353 6783
rect 4387 6749 4399 6783
rect 4341 6743 4399 6749
rect 2590 6672 2596 6724
rect 2648 6712 2654 6724
rect 4356 6712 4384 6743
rect 2648 6684 4384 6712
rect 4448 6712 4476 6820
rect 5445 6817 5457 6851
rect 5491 6848 5503 6851
rect 7653 6851 7711 6857
rect 7653 6848 7665 6851
rect 5491 6820 7665 6848
rect 5491 6817 5503 6820
rect 5445 6811 5503 6817
rect 7653 6817 7665 6820
rect 7699 6817 7711 6851
rect 7760 6848 7788 6876
rect 7837 6851 7895 6857
rect 7837 6848 7849 6851
rect 7760 6820 7849 6848
rect 7653 6811 7711 6817
rect 7837 6817 7849 6820
rect 7883 6817 7895 6851
rect 26418 6848 26424 6860
rect 7837 6811 7895 6817
rect 12406 6820 26424 6848
rect 5350 6780 5356 6792
rect 5263 6752 5356 6780
rect 5350 6740 5356 6752
rect 5408 6780 5414 6792
rect 5534 6780 5540 6792
rect 5408 6752 5540 6780
rect 5408 6740 5414 6752
rect 5534 6740 5540 6752
rect 5592 6740 5598 6792
rect 5997 6715 6055 6721
rect 5997 6712 6009 6715
rect 4448 6684 6009 6712
rect 2648 6672 2654 6684
rect 2317 6647 2375 6653
rect 2317 6613 2329 6647
rect 2363 6644 2375 6647
rect 3050 6644 3056 6656
rect 2363 6616 3056 6644
rect 2363 6613 2375 6616
rect 2317 6607 2375 6613
rect 3050 6604 3056 6616
rect 3108 6604 3114 6656
rect 4154 6604 4160 6656
rect 4212 6644 4218 6656
rect 4249 6647 4307 6653
rect 4249 6644 4261 6647
rect 4212 6616 4261 6644
rect 4212 6604 4218 6616
rect 4249 6613 4261 6616
rect 4295 6613 4307 6647
rect 4356 6644 4384 6684
rect 5997 6681 6009 6684
rect 6043 6681 6055 6715
rect 5997 6675 6055 6681
rect 12406 6644 12434 6820
rect 26418 6808 26424 6820
rect 26476 6808 26482 6860
rect 26513 6851 26571 6857
rect 26513 6817 26525 6851
rect 26559 6848 26571 6851
rect 27154 6848 27160 6860
rect 26559 6820 27160 6848
rect 26559 6817 26571 6820
rect 26513 6811 26571 6817
rect 27154 6808 27160 6820
rect 27212 6808 27218 6860
rect 28350 6848 28356 6860
rect 28311 6820 28356 6848
rect 28350 6808 28356 6820
rect 28408 6808 28414 6860
rect 25774 6740 25780 6792
rect 25832 6780 25838 6792
rect 25869 6783 25927 6789
rect 25869 6780 25881 6783
rect 25832 6752 25881 6780
rect 25832 6740 25838 6752
rect 25869 6749 25881 6752
rect 25915 6749 25927 6783
rect 25869 6743 25927 6749
rect 25961 6715 26019 6721
rect 25961 6681 25973 6715
rect 26007 6712 26019 6715
rect 26697 6715 26755 6721
rect 26697 6712 26709 6715
rect 26007 6684 26709 6712
rect 26007 6681 26019 6684
rect 25961 6675 26019 6681
rect 26697 6681 26709 6684
rect 26743 6681 26755 6715
rect 26697 6675 26755 6681
rect 4356 6616 12434 6644
rect 4249 6607 4307 6613
rect 1104 6554 29048 6576
rect 1104 6502 7896 6554
rect 7948 6502 7960 6554
rect 8012 6502 8024 6554
rect 8076 6502 8088 6554
rect 8140 6502 8152 6554
rect 8204 6502 14842 6554
rect 14894 6502 14906 6554
rect 14958 6502 14970 6554
rect 15022 6502 15034 6554
rect 15086 6502 15098 6554
rect 15150 6502 21788 6554
rect 21840 6502 21852 6554
rect 21904 6502 21916 6554
rect 21968 6502 21980 6554
rect 22032 6502 22044 6554
rect 22096 6502 28734 6554
rect 28786 6502 28798 6554
rect 28850 6502 28862 6554
rect 28914 6502 28926 6554
rect 28978 6502 28990 6554
rect 29042 6502 29048 6554
rect 1104 6480 29048 6502
rect 26694 6400 26700 6452
rect 26752 6440 26758 6452
rect 27249 6443 27307 6449
rect 27249 6440 27261 6443
rect 26752 6412 27261 6440
rect 26752 6400 26758 6412
rect 27249 6409 27261 6412
rect 27295 6409 27307 6443
rect 27249 6403 27307 6409
rect 4154 6372 4160 6384
rect 4115 6344 4160 6372
rect 4154 6332 4160 6344
rect 4212 6332 4218 6384
rect 1670 6304 1676 6316
rect 1631 6276 1676 6304
rect 1670 6264 1676 6276
rect 1728 6264 1734 6316
rect 26418 6264 26424 6316
rect 26476 6304 26482 6316
rect 27341 6307 27399 6313
rect 27341 6304 27353 6307
rect 26476 6276 27353 6304
rect 26476 6264 26482 6276
rect 27341 6273 27353 6276
rect 27387 6304 27399 6307
rect 27982 6304 27988 6316
rect 27387 6276 27988 6304
rect 27387 6273 27399 6276
rect 27341 6267 27399 6273
rect 27982 6264 27988 6276
rect 28040 6264 28046 6316
rect 1854 6236 1860 6248
rect 1815 6208 1860 6236
rect 1854 6196 1860 6208
rect 1912 6196 1918 6248
rect 3142 6236 3148 6248
rect 3103 6208 3148 6236
rect 3142 6196 3148 6208
rect 3200 6196 3206 6248
rect 3970 6236 3976 6248
rect 3931 6208 3976 6236
rect 3970 6196 3976 6208
rect 4028 6196 4034 6248
rect 4338 6196 4344 6248
rect 4396 6236 4402 6248
rect 4433 6239 4491 6245
rect 4433 6236 4445 6239
rect 4396 6208 4445 6236
rect 4396 6196 4402 6208
rect 4433 6205 4445 6208
rect 4479 6205 4491 6239
rect 4433 6199 4491 6205
rect 27893 6103 27951 6109
rect 27893 6069 27905 6103
rect 27939 6100 27951 6103
rect 28166 6100 28172 6112
rect 27939 6072 28172 6100
rect 27939 6069 27951 6072
rect 27893 6063 27951 6069
rect 28166 6060 28172 6072
rect 28224 6060 28230 6112
rect 1104 6010 28888 6032
rect 1104 5958 4423 6010
rect 4475 5958 4487 6010
rect 4539 5958 4551 6010
rect 4603 5958 4615 6010
rect 4667 5958 4679 6010
rect 4731 5958 11369 6010
rect 11421 5958 11433 6010
rect 11485 5958 11497 6010
rect 11549 5958 11561 6010
rect 11613 5958 11625 6010
rect 11677 5958 18315 6010
rect 18367 5958 18379 6010
rect 18431 5958 18443 6010
rect 18495 5958 18507 6010
rect 18559 5958 18571 6010
rect 18623 5958 25261 6010
rect 25313 5958 25325 6010
rect 25377 5958 25389 6010
rect 25441 5958 25453 6010
rect 25505 5958 25517 6010
rect 25569 5958 28888 6010
rect 1104 5936 28888 5958
rect 3970 5856 3976 5908
rect 4028 5896 4034 5908
rect 4065 5899 4123 5905
rect 4065 5896 4077 5899
rect 4028 5868 4077 5896
rect 4028 5856 4034 5868
rect 4065 5865 4077 5868
rect 4111 5865 4123 5899
rect 4065 5859 4123 5865
rect 1578 5760 1584 5772
rect 1539 5732 1584 5760
rect 1578 5720 1584 5732
rect 1636 5720 1642 5772
rect 2774 5760 2780 5772
rect 2735 5732 2780 5760
rect 2774 5720 2780 5732
rect 2832 5720 2838 5772
rect 27522 5760 27528 5772
rect 27483 5732 27528 5760
rect 27522 5720 27528 5732
rect 27580 5720 27586 5772
rect 28166 5760 28172 5772
rect 28127 5732 28172 5760
rect 28166 5720 28172 5732
rect 28224 5720 28230 5772
rect 28350 5652 28356 5704
rect 28408 5692 28414 5704
rect 28408 5664 28453 5692
rect 28408 5652 28414 5664
rect 1762 5624 1768 5636
rect 1723 5596 1768 5624
rect 1762 5584 1768 5596
rect 1820 5584 1826 5636
rect 1104 5466 29048 5488
rect 1104 5414 7896 5466
rect 7948 5414 7960 5466
rect 8012 5414 8024 5466
rect 8076 5414 8088 5466
rect 8140 5414 8152 5466
rect 8204 5414 14842 5466
rect 14894 5414 14906 5466
rect 14958 5414 14970 5466
rect 15022 5414 15034 5466
rect 15086 5414 15098 5466
rect 15150 5414 21788 5466
rect 21840 5414 21852 5466
rect 21904 5414 21916 5466
rect 21968 5414 21980 5466
rect 22032 5414 22044 5466
rect 22096 5414 28734 5466
rect 28786 5414 28798 5466
rect 28850 5414 28862 5466
rect 28914 5414 28926 5466
rect 28978 5414 28990 5466
rect 29042 5414 29048 5466
rect 1104 5392 29048 5414
rect 1762 5312 1768 5364
rect 1820 5352 1826 5364
rect 1949 5355 2007 5361
rect 1949 5352 1961 5355
rect 1820 5324 1961 5352
rect 1820 5312 1826 5324
rect 1949 5321 1961 5324
rect 1995 5321 2007 5355
rect 2498 5352 2504 5364
rect 1949 5315 2007 5321
rect 2056 5324 2504 5352
rect 2056 5228 2084 5324
rect 2498 5312 2504 5324
rect 2556 5352 2562 5364
rect 2556 5324 6914 5352
rect 2556 5312 2562 5324
rect 3050 5284 3056 5296
rect 3011 5256 3056 5284
rect 3050 5244 3056 5256
rect 3108 5244 3114 5296
rect 2038 5216 2044 5228
rect 1951 5188 2044 5216
rect 2038 5176 2044 5188
rect 2096 5176 2102 5228
rect 2866 5216 2872 5228
rect 2827 5188 2872 5216
rect 2866 5176 2872 5188
rect 2924 5176 2930 5228
rect 6886 5216 6914 5324
rect 12805 5219 12863 5225
rect 12805 5216 12817 5219
rect 6886 5188 12817 5216
rect 12805 5185 12817 5188
rect 12851 5185 12863 5219
rect 12805 5179 12863 5185
rect 28077 5219 28135 5225
rect 28077 5185 28089 5219
rect 28123 5216 28135 5219
rect 28350 5216 28356 5228
rect 28123 5188 28356 5216
rect 28123 5185 28135 5188
rect 28077 5179 28135 5185
rect 28350 5176 28356 5188
rect 28408 5176 28414 5228
rect 4709 5151 4767 5157
rect 4709 5117 4721 5151
rect 4755 5148 4767 5151
rect 4798 5148 4804 5160
rect 4755 5120 4804 5148
rect 4755 5117 4767 5120
rect 4709 5111 4767 5117
rect 4798 5108 4804 5120
rect 4856 5108 4862 5160
rect 4246 4972 4252 5024
rect 4304 5012 4310 5024
rect 5169 5015 5227 5021
rect 5169 5012 5181 5015
rect 4304 4984 5181 5012
rect 4304 4972 4310 4984
rect 5169 4981 5181 4984
rect 5215 4981 5227 5015
rect 5169 4975 5227 4981
rect 12897 5015 12955 5021
rect 12897 4981 12909 5015
rect 12943 5012 12955 5015
rect 12986 5012 12992 5024
rect 12943 4984 12992 5012
rect 12943 4981 12955 4984
rect 12897 4975 12955 4981
rect 12986 4972 12992 4984
rect 13044 4972 13050 5024
rect 1104 4922 28888 4944
rect 1104 4870 4423 4922
rect 4475 4870 4487 4922
rect 4539 4870 4551 4922
rect 4603 4870 4615 4922
rect 4667 4870 4679 4922
rect 4731 4870 11369 4922
rect 11421 4870 11433 4922
rect 11485 4870 11497 4922
rect 11549 4870 11561 4922
rect 11613 4870 11625 4922
rect 11677 4870 18315 4922
rect 18367 4870 18379 4922
rect 18431 4870 18443 4922
rect 18495 4870 18507 4922
rect 18559 4870 18571 4922
rect 18623 4870 25261 4922
rect 25313 4870 25325 4922
rect 25377 4870 25389 4922
rect 25441 4870 25453 4922
rect 25505 4870 25517 4922
rect 25569 4870 28888 4922
rect 1104 4848 28888 4870
rect 1854 4768 1860 4820
rect 1912 4808 1918 4820
rect 1949 4811 2007 4817
rect 1949 4808 1961 4811
rect 1912 4780 1961 4808
rect 1912 4768 1918 4780
rect 1949 4777 1961 4780
rect 1995 4777 2007 4811
rect 1949 4771 2007 4777
rect 4982 4672 4988 4684
rect 4816 4644 4988 4672
rect 2038 4604 2044 4616
rect 1999 4576 2044 4604
rect 2038 4564 2044 4576
rect 2096 4564 2102 4616
rect 3142 4604 3148 4616
rect 3103 4576 3148 4604
rect 3142 4564 3148 4576
rect 3200 4564 3206 4616
rect 3970 4604 3976 4616
rect 3931 4576 3976 4604
rect 3970 4564 3976 4576
rect 4028 4564 4034 4616
rect 4816 4613 4844 4644
rect 4982 4632 4988 4644
rect 5040 4672 5046 4684
rect 5718 4672 5724 4684
rect 5040 4644 5724 4672
rect 5040 4632 5046 4644
rect 5718 4632 5724 4644
rect 5776 4632 5782 4684
rect 20622 4672 20628 4684
rect 20583 4644 20628 4672
rect 20622 4632 20628 4644
rect 20680 4632 20686 4684
rect 21266 4672 21272 4684
rect 21227 4644 21272 4672
rect 21266 4632 21272 4644
rect 21324 4632 21330 4684
rect 27522 4672 27528 4684
rect 27483 4644 27528 4672
rect 27522 4632 27528 4644
rect 27580 4632 27586 4684
rect 4801 4607 4859 4613
rect 4801 4573 4813 4607
rect 4847 4573 4859 4607
rect 4801 4567 4859 4573
rect 4890 4564 4896 4616
rect 4948 4604 4954 4616
rect 5261 4607 5319 4613
rect 5261 4604 5273 4607
rect 4948 4576 5273 4604
rect 4948 4564 4954 4576
rect 5261 4573 5273 4576
rect 5307 4573 5319 4607
rect 5261 4567 5319 4573
rect 5534 4564 5540 4616
rect 5592 4604 5598 4616
rect 5997 4607 6055 4613
rect 5997 4604 6009 4607
rect 5592 4576 6009 4604
rect 5592 4564 5598 4576
rect 5997 4573 6009 4576
rect 6043 4604 6055 4607
rect 6043 4576 6914 4604
rect 6043 4573 6055 4576
rect 5997 4567 6055 4573
rect 6886 4536 6914 4576
rect 12802 4564 12808 4616
rect 12860 4604 12866 4616
rect 12897 4607 12955 4613
rect 12897 4604 12909 4607
rect 12860 4576 12909 4604
rect 12860 4564 12866 4576
rect 12897 4573 12909 4576
rect 12943 4573 12955 4607
rect 20438 4604 20444 4616
rect 20399 4576 20444 4604
rect 12897 4567 12955 4573
rect 20438 4564 20444 4576
rect 20496 4564 20502 4616
rect 25774 4604 25780 4616
rect 25735 4576 25780 4604
rect 25774 4564 25780 4576
rect 25832 4564 25838 4616
rect 26510 4604 26516 4616
rect 26471 4576 26516 4604
rect 26510 4564 26516 4576
rect 26568 4564 26574 4616
rect 16758 4536 16764 4548
rect 6886 4508 16764 4536
rect 16758 4496 16764 4508
rect 16816 4496 16822 4548
rect 26694 4536 26700 4548
rect 26655 4508 26700 4536
rect 26694 4496 26700 4508
rect 26752 4496 26758 4548
rect 4154 4428 4160 4480
rect 4212 4468 4218 4480
rect 4709 4471 4767 4477
rect 4709 4468 4721 4471
rect 4212 4440 4721 4468
rect 4212 4428 4218 4440
rect 4709 4437 4721 4440
rect 4755 4437 4767 4471
rect 4709 4431 4767 4437
rect 6089 4471 6147 4477
rect 6089 4437 6101 4471
rect 6135 4468 6147 4471
rect 6730 4468 6736 4480
rect 6135 4440 6736 4468
rect 6135 4437 6147 4440
rect 6089 4431 6147 4437
rect 6730 4428 6736 4440
rect 6788 4428 6794 4480
rect 25866 4468 25872 4480
rect 25827 4440 25872 4468
rect 25866 4428 25872 4440
rect 25924 4428 25930 4480
rect 1104 4378 29048 4400
rect 1104 4326 7896 4378
rect 7948 4326 7960 4378
rect 8012 4326 8024 4378
rect 8076 4326 8088 4378
rect 8140 4326 8152 4378
rect 8204 4326 14842 4378
rect 14894 4326 14906 4378
rect 14958 4326 14970 4378
rect 15022 4326 15034 4378
rect 15086 4326 15098 4378
rect 15150 4326 21788 4378
rect 21840 4326 21852 4378
rect 21904 4326 21916 4378
rect 21968 4326 21980 4378
rect 22032 4326 22044 4378
rect 22096 4326 28734 4378
rect 28786 4326 28798 4378
rect 28850 4326 28862 4378
rect 28914 4326 28926 4378
rect 28978 4326 28990 4378
rect 29042 4326 29048 4378
rect 1104 4304 29048 4326
rect 26694 4224 26700 4276
rect 26752 4264 26758 4276
rect 27249 4267 27307 4273
rect 27249 4264 27261 4267
rect 26752 4236 27261 4264
rect 26752 4224 26758 4236
rect 27249 4233 27261 4236
rect 27295 4233 27307 4267
rect 27249 4227 27307 4233
rect 4154 4196 4160 4208
rect 4115 4168 4160 4196
rect 4154 4156 4160 4168
rect 4212 4156 4218 4208
rect 12986 4196 12992 4208
rect 12947 4168 12992 4196
rect 12986 4156 12992 4168
rect 13044 4156 13050 4208
rect 3970 4128 3976 4140
rect 3931 4100 3976 4128
rect 3970 4088 3976 4100
rect 4028 4088 4034 4140
rect 11974 4128 11980 4140
rect 11935 4100 11980 4128
rect 11974 4088 11980 4100
rect 12032 4088 12038 4140
rect 12802 4128 12808 4140
rect 12763 4100 12808 4128
rect 12802 4088 12808 4100
rect 12860 4088 12866 4140
rect 17126 4128 17132 4140
rect 17087 4100 17132 4128
rect 17126 4088 17132 4100
rect 17184 4088 17190 4140
rect 20438 4088 20444 4140
rect 20496 4128 20502 4140
rect 20533 4131 20591 4137
rect 20533 4128 20545 4131
rect 20496 4100 20545 4128
rect 20496 4088 20502 4100
rect 20533 4097 20545 4100
rect 20579 4097 20591 4131
rect 20533 4091 20591 4097
rect 27341 4131 27399 4137
rect 27341 4097 27353 4131
rect 27387 4128 27399 4131
rect 27614 4128 27620 4140
rect 27387 4100 27620 4128
rect 27387 4097 27399 4100
rect 27341 4091 27399 4097
rect 27614 4088 27620 4100
rect 27672 4088 27678 4140
rect 658 4020 664 4072
rect 716 4060 722 4072
rect 1673 4063 1731 4069
rect 1673 4060 1685 4063
rect 716 4032 1685 4060
rect 716 4020 722 4032
rect 1673 4029 1685 4032
rect 1719 4029 1731 4063
rect 1673 4023 1731 4029
rect 1854 4020 1860 4072
rect 1912 4060 1918 4072
rect 3329 4063 3387 4069
rect 3329 4060 3341 4063
rect 1912 4032 3341 4060
rect 1912 4020 1918 4032
rect 3329 4029 3341 4032
rect 3375 4029 3387 4063
rect 3329 4023 3387 4029
rect 3513 4063 3571 4069
rect 3513 4029 3525 4063
rect 3559 4060 3571 4063
rect 4890 4060 4896 4072
rect 3559 4032 4896 4060
rect 3559 4029 3571 4032
rect 3513 4023 3571 4029
rect 4890 4020 4896 4032
rect 4948 4020 4954 4072
rect 4985 4063 5043 4069
rect 4985 4029 4997 4063
rect 5031 4029 5043 4063
rect 7742 4060 7748 4072
rect 7703 4032 7748 4060
rect 4985 4023 5043 4029
rect 3234 3952 3240 4004
rect 3292 3992 3298 4004
rect 5000 3992 5028 4023
rect 7742 4020 7748 4032
rect 7800 4020 7806 4072
rect 7929 4063 7987 4069
rect 7929 4029 7941 4063
rect 7975 4029 7987 4063
rect 8386 4060 8392 4072
rect 8347 4032 8392 4060
rect 7929 4023 7987 4029
rect 3292 3964 5028 3992
rect 3292 3952 3298 3964
rect 7650 3952 7656 4004
rect 7708 3992 7714 4004
rect 7944 3992 7972 4023
rect 8386 4020 8392 4032
rect 8444 4020 8450 4072
rect 7708 3964 7972 3992
rect 11992 3992 12020 4088
rect 13538 4060 13544 4072
rect 13499 4032 13544 4060
rect 13538 4020 13544 4032
rect 13596 4020 13602 4072
rect 16758 4020 16764 4072
rect 16816 4060 16822 4072
rect 25774 4060 25780 4072
rect 16816 4032 25780 4060
rect 16816 4020 16822 4032
rect 25774 4020 25780 4032
rect 25832 4020 25838 4072
rect 26142 4060 26148 4072
rect 26103 4032 26148 4060
rect 26142 4020 26148 4032
rect 26200 4020 26206 4072
rect 26418 4060 26424 4072
rect 26379 4032 26424 4060
rect 26418 4020 26424 4032
rect 26476 4020 26482 4072
rect 26605 4063 26663 4069
rect 26605 4029 26617 4063
rect 26651 4060 26663 4063
rect 27893 4063 27951 4069
rect 27893 4060 27905 4063
rect 26651 4032 27905 4060
rect 26651 4029 26663 4032
rect 26605 4023 26663 4029
rect 27893 4029 27905 4032
rect 27939 4029 27951 4063
rect 27893 4023 27951 4029
rect 14182 3992 14188 4004
rect 11992 3964 14188 3992
rect 7708 3952 7714 3964
rect 14182 3952 14188 3964
rect 14240 3952 14246 4004
rect 14550 3952 14556 4004
rect 14608 3992 14614 4004
rect 18690 3992 18696 4004
rect 14608 3964 18696 3992
rect 14608 3952 14614 3964
rect 18690 3952 18696 3964
rect 18748 3952 18754 4004
rect 6546 3924 6552 3936
rect 6507 3896 6552 3924
rect 6546 3884 6552 3896
rect 6604 3884 6610 3936
rect 12066 3924 12072 3936
rect 12027 3896 12072 3924
rect 12066 3884 12072 3896
rect 12124 3884 12130 3936
rect 17218 3924 17224 3936
rect 17179 3896 17224 3924
rect 17218 3884 17224 3896
rect 17276 3884 17282 3936
rect 1104 3834 28888 3856
rect 1104 3782 4423 3834
rect 4475 3782 4487 3834
rect 4539 3782 4551 3834
rect 4603 3782 4615 3834
rect 4667 3782 4679 3834
rect 4731 3782 11369 3834
rect 11421 3782 11433 3834
rect 11485 3782 11497 3834
rect 11549 3782 11561 3834
rect 11613 3782 11625 3834
rect 11677 3782 18315 3834
rect 18367 3782 18379 3834
rect 18431 3782 18443 3834
rect 18495 3782 18507 3834
rect 18559 3782 18571 3834
rect 18623 3782 25261 3834
rect 25313 3782 25325 3834
rect 25377 3782 25389 3834
rect 25441 3782 25453 3834
rect 25505 3782 25517 3834
rect 25569 3782 28888 3834
rect 1104 3760 28888 3782
rect 7742 3680 7748 3732
rect 7800 3720 7806 3732
rect 7837 3723 7895 3729
rect 7837 3720 7849 3723
rect 7800 3692 7849 3720
rect 7800 3680 7806 3692
rect 7837 3689 7849 3692
rect 7883 3689 7895 3723
rect 18046 3720 18052 3732
rect 18007 3692 18052 3720
rect 7837 3683 7895 3689
rect 18046 3680 18052 3692
rect 18104 3680 18110 3732
rect 25682 3720 25688 3732
rect 18248 3692 25688 3720
rect 3142 3544 3148 3596
rect 3200 3584 3206 3596
rect 3421 3587 3479 3593
rect 3421 3584 3433 3587
rect 3200 3556 3433 3584
rect 3200 3544 3206 3556
rect 3421 3553 3433 3556
rect 3467 3553 3479 3587
rect 5810 3584 5816 3596
rect 5771 3556 5816 3584
rect 3421 3547 3479 3553
rect 5810 3544 5816 3556
rect 5868 3544 5874 3596
rect 11882 3584 11888 3596
rect 11843 3556 11888 3584
rect 11882 3544 11888 3556
rect 11940 3544 11946 3596
rect 12066 3584 12072 3596
rect 12027 3556 12072 3584
rect 12066 3544 12072 3556
rect 12124 3544 12130 3596
rect 12434 3544 12440 3596
rect 12492 3584 12498 3596
rect 18248 3584 18276 3692
rect 25682 3680 25688 3692
rect 25740 3680 25746 3732
rect 26418 3680 26424 3732
rect 26476 3720 26482 3732
rect 28077 3723 28135 3729
rect 28077 3720 28089 3723
rect 26476 3692 28089 3720
rect 26476 3680 26482 3692
rect 28077 3689 28089 3692
rect 28123 3689 28135 3723
rect 28077 3683 28135 3689
rect 18690 3612 18696 3664
rect 18748 3652 18754 3664
rect 18748 3624 25728 3652
rect 18748 3612 18754 3624
rect 25700 3593 25728 3624
rect 25685 3587 25743 3593
rect 12492 3556 12537 3584
rect 17236 3556 18276 3584
rect 18432 3556 22048 3584
rect 12492 3544 12498 3556
rect 4617 3519 4675 3525
rect 4617 3485 4629 3519
rect 4663 3516 4675 3519
rect 5077 3519 5135 3525
rect 5077 3516 5089 3519
rect 4663 3488 5089 3516
rect 4663 3485 4675 3488
rect 4617 3479 4675 3485
rect 5077 3485 5089 3488
rect 5123 3485 5135 3519
rect 5077 3479 5135 3485
rect 8938 3476 8944 3528
rect 8996 3516 9002 3528
rect 9125 3519 9183 3525
rect 9125 3516 9137 3519
rect 8996 3488 9137 3516
rect 8996 3476 9002 3488
rect 9125 3485 9137 3488
rect 9171 3485 9183 3519
rect 9950 3516 9956 3528
rect 9911 3488 9956 3516
rect 9125 3479 9183 3485
rect 9950 3476 9956 3488
rect 10008 3476 10014 3528
rect 10594 3516 10600 3528
rect 10507 3488 10600 3516
rect 10594 3476 10600 3488
rect 10652 3516 10658 3528
rect 11425 3519 11483 3525
rect 10652 3488 11376 3516
rect 10652 3476 10658 3488
rect 1578 3448 1584 3460
rect 1539 3420 1584 3448
rect 1578 3408 1584 3420
rect 1636 3408 1642 3460
rect 2498 3408 2504 3460
rect 2556 3448 2562 3460
rect 3237 3451 3295 3457
rect 3237 3448 3249 3451
rect 2556 3420 3249 3448
rect 2556 3408 2562 3420
rect 3237 3417 3249 3420
rect 3283 3417 3295 3451
rect 5258 3448 5264 3460
rect 5219 3420 5264 3448
rect 3237 3411 3295 3417
rect 5258 3408 5264 3420
rect 5316 3408 5322 3460
rect 11348 3448 11376 3488
rect 11425 3485 11437 3519
rect 11471 3516 11483 3519
rect 11698 3516 11704 3528
rect 11471 3488 11704 3516
rect 11471 3485 11483 3488
rect 11425 3479 11483 3485
rect 11698 3476 11704 3488
rect 11756 3476 11762 3528
rect 14274 3476 14280 3528
rect 14332 3516 14338 3528
rect 14369 3519 14427 3525
rect 14369 3516 14381 3519
rect 14332 3488 14381 3516
rect 14332 3476 14338 3488
rect 14369 3485 14381 3488
rect 14415 3485 14427 3519
rect 16298 3516 16304 3528
rect 16259 3488 16304 3516
rect 14369 3479 14427 3485
rect 16298 3476 16304 3488
rect 16356 3476 16362 3528
rect 16758 3516 16764 3528
rect 16719 3488 16764 3516
rect 16758 3476 16764 3488
rect 16816 3476 16822 3528
rect 17236 3448 17264 3556
rect 17402 3516 17408 3528
rect 17363 3488 17408 3516
rect 17402 3476 17408 3488
rect 17460 3476 17466 3528
rect 17494 3476 17500 3528
rect 17552 3516 17558 3528
rect 18233 3519 18291 3525
rect 18233 3516 18245 3519
rect 17552 3488 18245 3516
rect 17552 3476 17558 3488
rect 18233 3485 18245 3488
rect 18279 3485 18291 3519
rect 18233 3479 18291 3485
rect 11348 3420 17264 3448
rect 9122 3340 9128 3392
rect 9180 3380 9186 3392
rect 9861 3383 9919 3389
rect 9861 3380 9873 3383
rect 9180 3352 9873 3380
rect 9180 3340 9186 3352
rect 9861 3349 9873 3352
rect 9907 3349 9919 3383
rect 9861 3343 9919 3349
rect 10689 3383 10747 3389
rect 10689 3349 10701 3383
rect 10735 3380 10747 3383
rect 11882 3380 11888 3392
rect 10735 3352 11888 3380
rect 10735 3349 10747 3352
rect 10689 3343 10747 3349
rect 11882 3340 11888 3352
rect 11940 3340 11946 3392
rect 16853 3383 16911 3389
rect 16853 3349 16865 3383
rect 16899 3380 16911 3383
rect 17034 3380 17040 3392
rect 16899 3352 17040 3380
rect 16899 3349 16911 3352
rect 16853 3343 16911 3349
rect 17034 3340 17040 3352
rect 17092 3340 17098 3392
rect 17126 3340 17132 3392
rect 17184 3380 17190 3392
rect 18432 3380 18460 3556
rect 19242 3476 19248 3528
rect 19300 3516 19306 3528
rect 19429 3519 19487 3525
rect 19429 3516 19441 3519
rect 19300 3488 19441 3516
rect 19300 3476 19306 3488
rect 19429 3485 19441 3488
rect 19475 3485 19487 3519
rect 19429 3479 19487 3485
rect 20257 3519 20315 3525
rect 20257 3485 20269 3519
rect 20303 3485 20315 3519
rect 21542 3516 21548 3528
rect 21503 3488 21548 3516
rect 20257 3479 20315 3485
rect 20272 3448 20300 3479
rect 21542 3476 21548 3488
rect 21600 3476 21606 3528
rect 22020 3525 22048 3556
rect 25685 3553 25697 3587
rect 25731 3553 25743 3587
rect 25866 3584 25872 3596
rect 25827 3556 25872 3584
rect 25685 3547 25743 3553
rect 25866 3544 25872 3556
rect 25924 3544 25930 3596
rect 22005 3519 22063 3525
rect 22005 3485 22017 3519
rect 22051 3485 22063 3519
rect 23842 3516 23848 3528
rect 23803 3488 23848 3516
rect 22005 3479 22063 3485
rect 23842 3476 23848 3488
rect 23900 3476 23906 3528
rect 24302 3476 24308 3528
rect 24360 3516 24366 3528
rect 24581 3519 24639 3525
rect 24581 3516 24593 3519
rect 24360 3488 24593 3516
rect 24360 3476 24366 3488
rect 24581 3485 24593 3488
rect 24627 3485 24639 3519
rect 27614 3516 27620 3528
rect 24581 3479 24639 3485
rect 27080 3488 27620 3516
rect 27080 3448 27108 3488
rect 27614 3476 27620 3488
rect 27672 3476 27678 3528
rect 27890 3476 27896 3528
rect 27948 3516 27954 3528
rect 27985 3519 28043 3525
rect 27985 3516 27997 3519
rect 27948 3488 27997 3516
rect 27948 3476 27954 3488
rect 27985 3485 27997 3488
rect 28031 3485 28043 3519
rect 27985 3479 28043 3485
rect 20272 3420 27108 3448
rect 27430 3408 27436 3460
rect 27488 3448 27494 3460
rect 27525 3451 27583 3457
rect 27525 3448 27537 3451
rect 27488 3420 27537 3448
rect 27488 3408 27494 3420
rect 27525 3417 27537 3420
rect 27571 3417 27583 3451
rect 27525 3411 27583 3417
rect 17184 3352 18460 3380
rect 17184 3340 17190 3352
rect 19426 3340 19432 3392
rect 19484 3380 19490 3392
rect 20165 3383 20223 3389
rect 20165 3380 20177 3383
rect 19484 3352 20177 3380
rect 19484 3340 19490 3352
rect 20165 3349 20177 3352
rect 20211 3349 20223 3383
rect 20165 3343 20223 3349
rect 22097 3383 22155 3389
rect 22097 3349 22109 3383
rect 22143 3380 22155 3383
rect 22186 3380 22192 3392
rect 22143 3352 22192 3380
rect 22143 3349 22155 3352
rect 22097 3343 22155 3349
rect 22186 3340 22192 3352
rect 22244 3340 22250 3392
rect 23937 3383 23995 3389
rect 23937 3349 23949 3383
rect 23983 3380 23995 3383
rect 24486 3380 24492 3392
rect 23983 3352 24492 3380
rect 23983 3349 23995 3352
rect 23937 3343 23995 3349
rect 24486 3340 24492 3352
rect 24544 3340 24550 3392
rect 1104 3290 29048 3312
rect 1104 3238 7896 3290
rect 7948 3238 7960 3290
rect 8012 3238 8024 3290
rect 8076 3238 8088 3290
rect 8140 3238 8152 3290
rect 8204 3238 14842 3290
rect 14894 3238 14906 3290
rect 14958 3238 14970 3290
rect 15022 3238 15034 3290
rect 15086 3238 15098 3290
rect 15150 3238 21788 3290
rect 21840 3238 21852 3290
rect 21904 3238 21916 3290
rect 21968 3238 21980 3290
rect 22032 3238 22044 3290
rect 22096 3238 28734 3290
rect 28786 3238 28798 3290
rect 28850 3238 28862 3290
rect 28914 3238 28926 3290
rect 28978 3238 28990 3290
rect 29042 3238 29048 3290
rect 1104 3216 29048 3238
rect 1854 3176 1860 3188
rect 1815 3148 1860 3176
rect 1854 3136 1860 3148
rect 1912 3136 1918 3188
rect 2498 3176 2504 3188
rect 2459 3148 2504 3176
rect 2498 3136 2504 3148
rect 2556 3136 2562 3188
rect 9950 3176 9956 3188
rect 6886 3148 9956 3176
rect 6886 3108 6914 3148
rect 9950 3136 9956 3148
rect 10008 3136 10014 3188
rect 14182 3136 14188 3188
rect 14240 3176 14246 3188
rect 17126 3176 17132 3188
rect 14240 3148 17132 3176
rect 14240 3136 14246 3148
rect 17126 3136 17132 3148
rect 17184 3136 17190 3188
rect 9122 3108 9128 3120
rect 2608 3080 6914 3108
rect 9083 3080 9128 3108
rect 2608 3049 2636 3080
rect 9122 3068 9128 3080
rect 9180 3068 9186 3120
rect 11882 3108 11888 3120
rect 11843 3080 11888 3108
rect 11882 3068 11888 3080
rect 11940 3068 11946 3120
rect 17034 3108 17040 3120
rect 16995 3080 17040 3108
rect 17034 3068 17040 3080
rect 17092 3068 17098 3120
rect 19426 3108 19432 3120
rect 19387 3080 19432 3108
rect 19426 3068 19432 3080
rect 19484 3068 19490 3120
rect 22186 3108 22192 3120
rect 22147 3080 22192 3108
rect 22186 3068 22192 3080
rect 22244 3068 22250 3120
rect 24486 3108 24492 3120
rect 24447 3080 24492 3108
rect 24486 3068 24492 3080
rect 24544 3068 24550 3120
rect 1949 3043 2007 3049
rect 1949 3009 1961 3043
rect 1995 3040 2007 3043
rect 2593 3043 2651 3049
rect 2593 3040 2605 3043
rect 1995 3012 2605 3040
rect 1995 3009 2007 3012
rect 1949 3003 2007 3009
rect 2593 3009 2605 3012
rect 2639 3009 2651 3043
rect 6546 3040 6552 3052
rect 6507 3012 6552 3040
rect 2593 3003 2651 3009
rect 6546 3000 6552 3012
rect 6604 3000 6610 3052
rect 8938 3040 8944 3052
rect 8899 3012 8944 3040
rect 8938 3000 8944 3012
rect 8996 3000 9002 3052
rect 11698 3040 11704 3052
rect 11659 3012 11704 3040
rect 11698 3000 11704 3012
rect 11756 3000 11762 3052
rect 14274 3040 14280 3052
rect 14235 3012 14280 3040
rect 14274 3000 14280 3012
rect 14332 3000 14338 3052
rect 16298 3000 16304 3052
rect 16356 3040 16362 3052
rect 16853 3043 16911 3049
rect 16853 3040 16865 3043
rect 16356 3012 16865 3040
rect 16356 3000 16362 3012
rect 16853 3009 16865 3012
rect 16899 3009 16911 3043
rect 19242 3040 19248 3052
rect 19203 3012 19248 3040
rect 16853 3003 16911 3009
rect 19242 3000 19248 3012
rect 19300 3000 19306 3052
rect 21542 3000 21548 3052
rect 21600 3040 21606 3052
rect 22005 3043 22063 3049
rect 22005 3040 22017 3043
rect 21600 3012 22017 3040
rect 21600 3000 21606 3012
rect 22005 3009 22017 3012
rect 22051 3009 22063 3043
rect 24302 3040 24308 3052
rect 24263 3012 24308 3040
rect 22005 3003 22063 3009
rect 24302 3000 24308 3012
rect 24360 3000 24366 3052
rect 26510 3000 26516 3052
rect 26568 3040 26574 3052
rect 27157 3043 27215 3049
rect 27157 3040 27169 3043
rect 26568 3012 27169 3040
rect 26568 3000 26574 3012
rect 27157 3009 27169 3012
rect 27203 3009 27215 3043
rect 27157 3003 27215 3009
rect 27890 3000 27896 3052
rect 27948 3040 27954 3052
rect 27985 3043 28043 3049
rect 27985 3040 27997 3043
rect 27948 3012 27997 3040
rect 27948 3000 27954 3012
rect 27985 3009 27997 3012
rect 28031 3009 28043 3043
rect 27985 3003 28043 3009
rect 3237 2975 3295 2981
rect 3237 2941 3249 2975
rect 3283 2972 3295 2975
rect 3697 2975 3755 2981
rect 3697 2972 3709 2975
rect 3283 2944 3709 2972
rect 3283 2941 3295 2944
rect 3237 2935 3295 2941
rect 3697 2941 3709 2944
rect 3743 2941 3755 2975
rect 3878 2972 3884 2984
rect 3839 2944 3884 2972
rect 3697 2935 3755 2941
rect 3878 2932 3884 2944
rect 3936 2932 3942 2984
rect 3970 2932 3976 2984
rect 4028 2972 4034 2984
rect 4157 2975 4215 2981
rect 4157 2972 4169 2975
rect 4028 2944 4169 2972
rect 4028 2932 4034 2944
rect 4157 2941 4169 2944
rect 4203 2941 4215 2975
rect 6730 2972 6736 2984
rect 6691 2944 6736 2972
rect 4157 2935 4215 2941
rect 6730 2932 6736 2944
rect 6788 2932 6794 2984
rect 7009 2975 7067 2981
rect 7009 2972 7021 2975
rect 6886 2944 7021 2972
rect 6454 2864 6460 2916
rect 6512 2904 6518 2916
rect 6886 2904 6914 2944
rect 7009 2941 7021 2944
rect 7055 2941 7067 2975
rect 9674 2972 9680 2984
rect 9635 2944 9680 2972
rect 7009 2935 7067 2941
rect 9674 2932 9680 2944
rect 9732 2932 9738 2984
rect 10962 2932 10968 2984
rect 11020 2972 11026 2984
rect 12161 2975 12219 2981
rect 12161 2972 12173 2975
rect 11020 2944 12173 2972
rect 11020 2932 11026 2944
rect 12161 2941 12173 2944
rect 12207 2941 12219 2975
rect 14458 2972 14464 2984
rect 14419 2944 14464 2972
rect 12161 2935 12219 2941
rect 14458 2932 14464 2944
rect 14516 2932 14522 2984
rect 14734 2972 14740 2984
rect 14695 2944 14740 2972
rect 14734 2932 14740 2944
rect 14792 2932 14798 2984
rect 16758 2932 16764 2984
rect 16816 2972 16822 2984
rect 17313 2975 17371 2981
rect 17313 2972 17325 2975
rect 16816 2944 17325 2972
rect 16816 2932 16822 2944
rect 17313 2941 17325 2944
rect 17359 2941 17371 2975
rect 19978 2972 19984 2984
rect 19939 2944 19984 2972
rect 17313 2935 17371 2941
rect 19978 2932 19984 2944
rect 20036 2932 20042 2984
rect 22465 2975 22523 2981
rect 22465 2972 22477 2975
rect 22066 2944 22477 2972
rect 6512 2876 6914 2904
rect 6512 2864 6518 2876
rect 21634 2864 21640 2916
rect 21692 2904 21698 2916
rect 22066 2904 22094 2944
rect 22465 2941 22477 2944
rect 22511 2941 22523 2975
rect 25130 2972 25136 2984
rect 25091 2944 25136 2972
rect 22465 2935 22523 2941
rect 25130 2932 25136 2944
rect 25188 2932 25194 2984
rect 21692 2876 22094 2904
rect 21692 2864 21698 2876
rect 2590 2796 2596 2848
rect 2648 2836 2654 2848
rect 4798 2836 4804 2848
rect 2648 2808 4804 2836
rect 2648 2796 2654 2808
rect 4798 2796 4804 2808
rect 4856 2796 4862 2848
rect 26418 2796 26424 2848
rect 26476 2836 26482 2848
rect 27893 2839 27951 2845
rect 27893 2836 27905 2839
rect 26476 2808 27905 2836
rect 26476 2796 26482 2808
rect 27893 2805 27905 2808
rect 27939 2805 27951 2839
rect 27893 2799 27951 2805
rect 1104 2746 28888 2768
rect 1104 2694 4423 2746
rect 4475 2694 4487 2746
rect 4539 2694 4551 2746
rect 4603 2694 4615 2746
rect 4667 2694 4679 2746
rect 4731 2694 11369 2746
rect 11421 2694 11433 2746
rect 11485 2694 11497 2746
rect 11549 2694 11561 2746
rect 11613 2694 11625 2746
rect 11677 2694 18315 2746
rect 18367 2694 18379 2746
rect 18431 2694 18443 2746
rect 18495 2694 18507 2746
rect 18559 2694 18571 2746
rect 18623 2694 25261 2746
rect 25313 2694 25325 2746
rect 25377 2694 25389 2746
rect 25441 2694 25453 2746
rect 25505 2694 25517 2746
rect 25569 2694 28888 2746
rect 1104 2672 28888 2694
rect 3878 2592 3884 2644
rect 3936 2632 3942 2644
rect 4065 2635 4123 2641
rect 4065 2632 4077 2635
rect 3936 2604 4077 2632
rect 3936 2592 3942 2604
rect 4065 2601 4077 2604
rect 4111 2601 4123 2635
rect 5258 2632 5264 2644
rect 5219 2604 5264 2632
rect 4065 2595 4123 2601
rect 5258 2592 5264 2604
rect 5316 2592 5322 2644
rect 7650 2592 7656 2644
rect 7708 2632 7714 2644
rect 8021 2635 8079 2641
rect 8021 2632 8033 2635
rect 7708 2604 8033 2632
rect 7708 2592 7714 2604
rect 8021 2601 8033 2604
rect 8067 2601 8079 2635
rect 8021 2595 8079 2601
rect 14369 2635 14427 2641
rect 14369 2601 14381 2635
rect 14415 2632 14427 2635
rect 14458 2632 14464 2644
rect 14415 2604 14464 2632
rect 14415 2601 14427 2604
rect 14369 2595 14427 2601
rect 14458 2592 14464 2604
rect 14516 2592 14522 2644
rect 16209 2635 16267 2641
rect 16209 2601 16221 2635
rect 16255 2632 16267 2635
rect 16850 2632 16856 2644
rect 16255 2604 16856 2632
rect 16255 2601 16267 2604
rect 16209 2595 16267 2601
rect 16850 2592 16856 2604
rect 16908 2592 16914 2644
rect 23842 2632 23848 2644
rect 16960 2604 23848 2632
rect 2314 2524 2320 2576
rect 2372 2564 2378 2576
rect 16960 2564 16988 2604
rect 23842 2592 23848 2604
rect 23900 2592 23906 2644
rect 27062 2592 27068 2644
rect 27120 2632 27126 2644
rect 27157 2635 27215 2641
rect 27157 2632 27169 2635
rect 27120 2604 27169 2632
rect 27120 2592 27126 2604
rect 27157 2601 27169 2604
rect 27203 2601 27215 2635
rect 27157 2595 27215 2601
rect 17402 2564 17408 2576
rect 2372 2536 16988 2564
rect 17052 2536 17408 2564
rect 2372 2524 2378 2536
rect 2774 2456 2780 2508
rect 2832 2496 2838 2508
rect 3421 2499 3479 2505
rect 2832 2468 2877 2496
rect 2832 2456 2838 2468
rect 3421 2465 3433 2499
rect 3467 2496 3479 2499
rect 3786 2496 3792 2508
rect 3467 2468 3792 2496
rect 3467 2465 3479 2468
rect 3421 2459 3479 2465
rect 3786 2456 3792 2468
rect 3844 2456 3850 2508
rect 4154 2428 4160 2440
rect 4115 2400 4160 2428
rect 4154 2388 4160 2400
rect 4212 2388 4218 2440
rect 5169 2431 5227 2437
rect 5169 2397 5181 2431
rect 5215 2430 5227 2431
rect 5276 2430 5304 2536
rect 9398 2496 9404 2508
rect 9359 2468 9404 2496
rect 9398 2456 9404 2468
rect 9456 2456 9462 2508
rect 17052 2505 17080 2536
rect 17402 2524 17408 2536
rect 17460 2524 17466 2576
rect 17037 2499 17095 2505
rect 17037 2465 17049 2499
rect 17083 2465 17095 2499
rect 17218 2496 17224 2508
rect 17179 2468 17224 2496
rect 17037 2459 17095 2465
rect 17218 2456 17224 2468
rect 17276 2456 17282 2508
rect 18046 2496 18052 2508
rect 18007 2468 18052 2496
rect 18046 2456 18052 2468
rect 18104 2456 18110 2508
rect 26142 2496 26148 2508
rect 26103 2468 26148 2496
rect 26142 2456 26148 2468
rect 26200 2456 26206 2508
rect 26418 2496 26424 2508
rect 26379 2468 26424 2496
rect 26418 2456 26424 2468
rect 26476 2456 26482 2508
rect 26605 2499 26663 2505
rect 26605 2465 26617 2499
rect 26651 2496 26663 2499
rect 27801 2499 27859 2505
rect 27801 2496 27813 2499
rect 26651 2468 27813 2496
rect 26651 2465 26663 2468
rect 26605 2459 26663 2465
rect 27801 2465 27813 2468
rect 27847 2465 27859 2499
rect 27801 2459 27859 2465
rect 5215 2402 5304 2430
rect 5215 2397 5227 2402
rect 5169 2391 5227 2397
rect 5718 2388 5724 2440
rect 5776 2428 5782 2440
rect 5997 2431 6055 2437
rect 5997 2428 6009 2431
rect 5776 2400 6009 2428
rect 5776 2388 5782 2400
rect 5997 2397 6009 2400
rect 6043 2428 6055 2431
rect 8113 2431 8171 2437
rect 8113 2428 8125 2431
rect 6043 2400 8125 2428
rect 6043 2397 6055 2400
rect 5997 2391 6055 2397
rect 8113 2397 8125 2400
rect 8159 2397 8171 2431
rect 8113 2391 8171 2397
rect 9030 2388 9036 2440
rect 9088 2428 9094 2440
rect 9125 2431 9183 2437
rect 9125 2428 9137 2431
rect 9088 2400 9137 2428
rect 9088 2388 9094 2400
rect 9125 2397 9137 2400
rect 9171 2397 9183 2431
rect 9125 2391 9183 2397
rect 14182 2388 14188 2440
rect 14240 2428 14246 2440
rect 14277 2431 14335 2437
rect 14277 2428 14289 2431
rect 14240 2400 14289 2428
rect 14240 2388 14246 2400
rect 14277 2397 14289 2400
rect 14323 2397 14335 2431
rect 14277 2391 14335 2397
rect 27062 2388 27068 2440
rect 27120 2428 27126 2440
rect 27341 2431 27399 2437
rect 27341 2428 27353 2431
rect 27120 2400 27353 2428
rect 27120 2388 27126 2400
rect 27341 2397 27353 2400
rect 27387 2397 27399 2431
rect 27341 2391 27399 2397
rect 3237 2363 3295 2369
rect 3237 2329 3249 2363
rect 3283 2360 3295 2363
rect 5905 2363 5963 2369
rect 5905 2360 5917 2363
rect 3283 2332 5917 2360
rect 3283 2329 3295 2332
rect 3237 2323 3295 2329
rect 5905 2329 5917 2332
rect 5951 2329 5963 2363
rect 16114 2360 16120 2372
rect 16075 2332 16120 2360
rect 5905 2323 5963 2329
rect 16114 2320 16120 2332
rect 16172 2320 16178 2372
rect 4062 2252 4068 2304
rect 4120 2292 4126 2304
rect 12434 2292 12440 2304
rect 4120 2264 12440 2292
rect 4120 2252 4126 2264
rect 12434 2252 12440 2264
rect 12492 2252 12498 2304
rect 1104 2202 29048 2224
rect 1104 2150 7896 2202
rect 7948 2150 7960 2202
rect 8012 2150 8024 2202
rect 8076 2150 8088 2202
rect 8140 2150 8152 2202
rect 8204 2150 14842 2202
rect 14894 2150 14906 2202
rect 14958 2150 14970 2202
rect 15022 2150 15034 2202
rect 15086 2150 15098 2202
rect 15150 2150 21788 2202
rect 21840 2150 21852 2202
rect 21904 2150 21916 2202
rect 21968 2150 21980 2202
rect 22032 2150 22044 2202
rect 22096 2150 28734 2202
rect 28786 2150 28798 2202
rect 28850 2150 28862 2202
rect 28914 2150 28926 2202
rect 28978 2150 28990 2202
rect 29042 2150 29048 2202
rect 1104 2128 29048 2150
rect 4154 2048 4160 2100
rect 4212 2088 4218 2100
rect 10594 2088 10600 2100
rect 4212 2060 10600 2088
rect 4212 2048 4218 2060
rect 10594 2048 10600 2060
rect 10652 2048 10658 2100
<< via1 >>
rect 20 47404 72 47456
rect 940 47404 992 47456
rect 4423 47302 4475 47354
rect 4487 47302 4539 47354
rect 4551 47302 4603 47354
rect 4615 47302 4667 47354
rect 4679 47302 4731 47354
rect 11369 47302 11421 47354
rect 11433 47302 11485 47354
rect 11497 47302 11549 47354
rect 11561 47302 11613 47354
rect 11625 47302 11677 47354
rect 18315 47302 18367 47354
rect 18379 47302 18431 47354
rect 18443 47302 18495 47354
rect 18507 47302 18559 47354
rect 18571 47302 18623 47354
rect 25261 47302 25313 47354
rect 25325 47302 25377 47354
rect 25389 47302 25441 47354
rect 25453 47302 25505 47354
rect 25517 47302 25569 47354
rect 22192 47132 22244 47184
rect 1952 47107 2004 47116
rect 1952 47073 1961 47107
rect 1961 47073 1995 47107
rect 1995 47073 2004 47107
rect 1952 47064 2004 47073
rect 10324 47107 10376 47116
rect 10324 47073 10333 47107
rect 10333 47073 10367 47107
rect 10367 47073 10376 47107
rect 10324 47064 10376 47073
rect 3516 46996 3568 47048
rect 5816 47039 5868 47048
rect 5816 47005 5825 47039
rect 5825 47005 5859 47039
rect 5859 47005 5868 47039
rect 5816 46996 5868 47005
rect 6460 46996 6512 47048
rect 7012 46996 7064 47048
rect 9312 47039 9364 47048
rect 9312 47005 9321 47039
rect 9321 47005 9355 47039
rect 9355 47005 9364 47039
rect 9312 46996 9364 47005
rect 11704 47039 11756 47048
rect 11704 47005 11713 47039
rect 11713 47005 11747 47039
rect 11747 47005 11756 47039
rect 11704 46996 11756 47005
rect 13912 46996 13964 47048
rect 14372 46996 14424 47048
rect 16856 47039 16908 47048
rect 16856 47005 16865 47039
rect 16865 47005 16899 47039
rect 16899 47005 16908 47039
rect 16856 46996 16908 47005
rect 18512 47039 18564 47048
rect 18512 47005 18521 47039
rect 18521 47005 18555 47039
rect 18555 47005 18564 47039
rect 18512 46996 18564 47005
rect 20812 47039 20864 47048
rect 20812 47005 20821 47039
rect 20821 47005 20855 47039
rect 20855 47005 20864 47039
rect 20812 46996 20864 47005
rect 22468 47064 22520 47116
rect 23204 47107 23256 47116
rect 23204 47073 23213 47107
rect 23213 47073 23247 47107
rect 23247 47073 23256 47107
rect 23204 47064 23256 47073
rect 26608 47107 26660 47116
rect 26608 47073 26617 47107
rect 26617 47073 26651 47107
rect 26651 47073 26660 47107
rect 26608 47064 26660 47073
rect 24768 47039 24820 47048
rect 24768 47005 24777 47039
rect 24777 47005 24811 47039
rect 24811 47005 24820 47039
rect 24768 46996 24820 47005
rect 27436 46996 27488 47048
rect 27804 47039 27856 47048
rect 27804 47005 27813 47039
rect 27813 47005 27847 47039
rect 27847 47005 27856 47039
rect 27804 46996 27856 47005
rect 3240 46971 3292 46980
rect 3240 46937 3249 46971
rect 3249 46937 3283 46971
rect 3283 46937 3292 46971
rect 3240 46928 3292 46937
rect 9864 46928 9916 46980
rect 23020 46928 23072 46980
rect 24952 46971 25004 46980
rect 24952 46937 24961 46971
rect 24961 46937 24995 46971
rect 24995 46937 25004 46971
rect 24952 46928 25004 46937
rect 26700 46928 26752 46980
rect 6000 46903 6052 46912
rect 6000 46869 6009 46903
rect 6009 46869 6043 46903
rect 6043 46869 6052 46903
rect 6000 46860 6052 46869
rect 6736 46903 6788 46912
rect 6736 46869 6745 46903
rect 6745 46869 6779 46903
rect 6779 46869 6788 46903
rect 6736 46860 6788 46869
rect 7896 46758 7948 46810
rect 7960 46758 8012 46810
rect 8024 46758 8076 46810
rect 8088 46758 8140 46810
rect 8152 46758 8204 46810
rect 14842 46758 14894 46810
rect 14906 46758 14958 46810
rect 14970 46758 15022 46810
rect 15034 46758 15086 46810
rect 15098 46758 15150 46810
rect 21788 46758 21840 46810
rect 21852 46758 21904 46810
rect 21916 46758 21968 46810
rect 21980 46758 22032 46810
rect 22044 46758 22096 46810
rect 28734 46758 28786 46810
rect 28798 46758 28850 46810
rect 28862 46758 28914 46810
rect 28926 46758 28978 46810
rect 28990 46758 29042 46810
rect 26700 46588 26752 46640
rect 7012 46563 7064 46572
rect 7012 46529 7021 46563
rect 7021 46529 7055 46563
rect 7055 46529 7064 46563
rect 7012 46520 7064 46529
rect 13912 46563 13964 46572
rect 13912 46529 13921 46563
rect 13921 46529 13955 46563
rect 13955 46529 13964 46563
rect 14372 46563 14424 46572
rect 13912 46520 13964 46529
rect 14372 46529 14381 46563
rect 14381 46529 14415 46563
rect 14415 46529 14424 46563
rect 14372 46520 14424 46529
rect 16856 46563 16908 46572
rect 16856 46529 16865 46563
rect 16865 46529 16899 46563
rect 16899 46529 16908 46563
rect 16856 46520 16908 46529
rect 18512 46520 18564 46572
rect 20812 46520 20864 46572
rect 27620 46588 27672 46640
rect 27160 46563 27212 46572
rect 4068 46452 4120 46504
rect 2596 46384 2648 46436
rect 7840 46452 7892 46504
rect 8392 46495 8444 46504
rect 8392 46461 8401 46495
rect 8401 46461 8435 46495
rect 8435 46461 8444 46495
rect 8392 46452 8444 46461
rect 10508 46452 10560 46504
rect 10968 46495 11020 46504
rect 10968 46461 10977 46495
rect 10977 46461 11011 46495
rect 11011 46461 11020 46495
rect 10968 46452 11020 46461
rect 13452 46495 13504 46504
rect 13452 46461 13461 46495
rect 13461 46461 13495 46495
rect 13495 46461 13504 46495
rect 13452 46452 13504 46461
rect 13544 46452 13596 46504
rect 14556 46495 14608 46504
rect 14556 46461 14565 46495
rect 14565 46461 14599 46495
rect 14599 46461 14608 46495
rect 14556 46452 14608 46461
rect 14740 46452 14792 46504
rect 16396 46452 16448 46504
rect 19340 46495 19392 46504
rect 10324 46384 10376 46436
rect 16764 46384 16816 46436
rect 19340 46461 19349 46495
rect 19349 46461 19383 46495
rect 19383 46461 19392 46495
rect 19340 46452 19392 46461
rect 18696 46384 18748 46436
rect 22376 46452 22428 46504
rect 21272 46384 21324 46436
rect 24308 46452 24360 46504
rect 1584 46316 1636 46368
rect 10600 46316 10652 46368
rect 18144 46316 18196 46368
rect 27160 46529 27169 46563
rect 27169 46529 27203 46563
rect 27203 46529 27212 46563
rect 27160 46520 27212 46529
rect 28356 46452 28408 46504
rect 26700 46384 26752 46436
rect 26424 46316 26476 46368
rect 4423 46214 4475 46266
rect 4487 46214 4539 46266
rect 4551 46214 4603 46266
rect 4615 46214 4667 46266
rect 4679 46214 4731 46266
rect 11369 46214 11421 46266
rect 11433 46214 11485 46266
rect 11497 46214 11549 46266
rect 11561 46214 11613 46266
rect 11625 46214 11677 46266
rect 18315 46214 18367 46266
rect 18379 46214 18431 46266
rect 18443 46214 18495 46266
rect 18507 46214 18559 46266
rect 18571 46214 18623 46266
rect 25261 46214 25313 46266
rect 25325 46214 25377 46266
rect 25389 46214 25441 46266
rect 25453 46214 25505 46266
rect 25517 46214 25569 46266
rect 4068 46155 4120 46164
rect 4068 46121 4077 46155
rect 4077 46121 4111 46155
rect 4111 46121 4120 46155
rect 4068 46112 4120 46121
rect 7840 46155 7892 46164
rect 7840 46121 7849 46155
rect 7849 46121 7883 46155
rect 7883 46121 7892 46155
rect 7840 46112 7892 46121
rect 9864 46155 9916 46164
rect 9864 46121 9873 46155
rect 9873 46121 9907 46155
rect 9907 46121 9916 46155
rect 9864 46112 9916 46121
rect 10508 46155 10560 46164
rect 10508 46121 10517 46155
rect 10517 46121 10551 46155
rect 10551 46121 10560 46155
rect 10508 46112 10560 46121
rect 13544 46155 13596 46164
rect 13544 46121 13553 46155
rect 13553 46121 13587 46155
rect 13587 46121 13596 46155
rect 13544 46112 13596 46121
rect 14556 46155 14608 46164
rect 14556 46121 14565 46155
rect 14565 46121 14599 46155
rect 14599 46121 14608 46155
rect 14556 46112 14608 46121
rect 16396 46155 16448 46164
rect 16396 46121 16405 46155
rect 16405 46121 16439 46155
rect 16439 46121 16448 46155
rect 16396 46112 16448 46121
rect 19340 46112 19392 46164
rect 27344 46112 27396 46164
rect 1584 46019 1636 46028
rect 1584 45985 1593 46019
rect 1593 45985 1627 46019
rect 1627 45985 1636 46019
rect 1584 45976 1636 45985
rect 2964 46019 3016 46028
rect 2964 45985 2973 46019
rect 2973 45985 3007 46019
rect 3007 45985 3016 46019
rect 2964 45976 3016 45985
rect 4804 45908 4856 45960
rect 7748 45908 7800 45960
rect 11704 45976 11756 46028
rect 11796 46019 11848 46028
rect 11796 45985 11805 46019
rect 11805 45985 11839 46019
rect 11839 45985 11848 46019
rect 11796 45976 11848 45985
rect 9956 45951 10008 45960
rect 9956 45917 9965 45951
rect 9965 45917 9999 45951
rect 9999 45917 10008 45951
rect 10600 45951 10652 45960
rect 9956 45908 10008 45917
rect 10600 45917 10609 45951
rect 10609 45917 10643 45951
rect 10643 45917 10652 45951
rect 10600 45908 10652 45917
rect 13636 45951 13688 45960
rect 13636 45917 13645 45951
rect 13645 45917 13679 45951
rect 13679 45917 13688 45951
rect 13636 45908 13688 45917
rect 1952 45840 2004 45892
rect 11796 45840 11848 45892
rect 22192 46044 22244 46096
rect 19984 46019 20036 46028
rect 19984 45985 19993 46019
rect 19993 45985 20027 46019
rect 20027 45985 20036 46019
rect 19984 45976 20036 45985
rect 22560 46019 22612 46028
rect 22560 45985 22569 46019
rect 22569 45985 22603 46019
rect 22603 45985 22612 46019
rect 22560 45976 22612 45985
rect 27068 45976 27120 46028
rect 27436 46019 27488 46028
rect 27436 45985 27445 46019
rect 27445 45985 27479 46019
rect 27479 45985 27488 46019
rect 27436 45976 27488 45985
rect 14464 45951 14516 45960
rect 14464 45917 14473 45951
rect 14473 45917 14507 45951
rect 14507 45917 14516 45951
rect 14464 45908 14516 45917
rect 18144 45908 18196 45960
rect 19432 45951 19484 45960
rect 19432 45917 19441 45951
rect 19441 45917 19475 45951
rect 19475 45917 19484 45951
rect 19432 45908 19484 45917
rect 23848 45908 23900 45960
rect 27528 45908 27580 45960
rect 19616 45883 19668 45892
rect 19616 45849 19625 45883
rect 19625 45849 19659 45883
rect 19659 45849 19668 45883
rect 19616 45840 19668 45849
rect 22284 45883 22336 45892
rect 22284 45849 22293 45883
rect 22293 45849 22327 45883
rect 22327 45849 22336 45883
rect 22284 45840 22336 45849
rect 25136 45840 25188 45892
rect 27252 45883 27304 45892
rect 27252 45849 27261 45883
rect 27261 45849 27295 45883
rect 27295 45849 27304 45883
rect 27252 45840 27304 45849
rect 23572 45772 23624 45824
rect 7896 45670 7948 45722
rect 7960 45670 8012 45722
rect 8024 45670 8076 45722
rect 8088 45670 8140 45722
rect 8152 45670 8204 45722
rect 14842 45670 14894 45722
rect 14906 45670 14958 45722
rect 14970 45670 15022 45722
rect 15034 45670 15086 45722
rect 15098 45670 15150 45722
rect 21788 45670 21840 45722
rect 21852 45670 21904 45722
rect 21916 45670 21968 45722
rect 21980 45670 22032 45722
rect 22044 45670 22096 45722
rect 28734 45670 28786 45722
rect 28798 45670 28850 45722
rect 28862 45670 28914 45722
rect 28926 45670 28978 45722
rect 28990 45670 29042 45722
rect 1952 45611 2004 45620
rect 1952 45577 1961 45611
rect 1961 45577 1995 45611
rect 1995 45577 2004 45611
rect 1952 45568 2004 45577
rect 11796 45611 11848 45620
rect 2412 45500 2464 45552
rect 3240 45500 3292 45552
rect 11796 45577 11805 45611
rect 11805 45577 11839 45611
rect 11839 45577 11848 45611
rect 11796 45568 11848 45577
rect 19616 45568 19668 45620
rect 22284 45568 22336 45620
rect 27252 45611 27304 45620
rect 27252 45577 27261 45611
rect 27261 45577 27295 45611
rect 27295 45577 27304 45611
rect 27252 45568 27304 45577
rect 13636 45500 13688 45552
rect 23020 45543 23072 45552
rect 2320 45364 2372 45416
rect 3516 45432 3568 45484
rect 9312 45432 9364 45484
rect 10324 45475 10376 45484
rect 10324 45441 10333 45475
rect 10333 45441 10367 45475
rect 10367 45441 10376 45475
rect 10324 45432 10376 45441
rect 11888 45475 11940 45484
rect 11888 45441 11897 45475
rect 11897 45441 11931 45475
rect 11931 45441 11940 45475
rect 19340 45475 19392 45484
rect 11888 45432 11940 45441
rect 9956 45364 10008 45416
rect 19340 45441 19349 45475
rect 19349 45441 19383 45475
rect 19383 45441 19392 45475
rect 19340 45432 19392 45441
rect 19432 45432 19484 45484
rect 20628 45475 20680 45484
rect 20628 45441 20637 45475
rect 20637 45441 20671 45475
rect 20671 45441 20680 45475
rect 20628 45432 20680 45441
rect 22376 45432 22428 45484
rect 23020 45509 23029 45543
rect 23029 45509 23063 45543
rect 23063 45509 23072 45543
rect 23020 45500 23072 45509
rect 26240 45500 26292 45552
rect 26424 45543 26476 45552
rect 26424 45509 26433 45543
rect 26433 45509 26467 45543
rect 26467 45509 26476 45543
rect 26424 45500 26476 45509
rect 23112 45475 23164 45484
rect 23112 45441 23121 45475
rect 23121 45441 23155 45475
rect 23155 45441 23164 45475
rect 23112 45432 23164 45441
rect 24308 45475 24360 45484
rect 24308 45441 24317 45475
rect 24317 45441 24351 45475
rect 24351 45441 24360 45475
rect 24308 45432 24360 45441
rect 26700 45432 26752 45484
rect 27344 45475 27396 45484
rect 27344 45441 27353 45475
rect 27353 45441 27387 45475
rect 27387 45441 27396 45475
rect 27344 45432 27396 45441
rect 25780 45364 25832 45416
rect 27712 45568 27764 45620
rect 27896 45475 27948 45484
rect 27896 45441 27905 45475
rect 27905 45441 27939 45475
rect 27939 45441 27948 45475
rect 27896 45432 27948 45441
rect 20628 45296 20680 45348
rect 27160 45296 27212 45348
rect 26424 45228 26476 45280
rect 4423 45126 4475 45178
rect 4487 45126 4539 45178
rect 4551 45126 4603 45178
rect 4615 45126 4667 45178
rect 4679 45126 4731 45178
rect 11369 45126 11421 45178
rect 11433 45126 11485 45178
rect 11497 45126 11549 45178
rect 11561 45126 11613 45178
rect 11625 45126 11677 45178
rect 18315 45126 18367 45178
rect 18379 45126 18431 45178
rect 18443 45126 18495 45178
rect 18507 45126 18559 45178
rect 18571 45126 18623 45178
rect 25261 45126 25313 45178
rect 25325 45126 25377 45178
rect 25389 45126 25441 45178
rect 25453 45126 25505 45178
rect 25517 45126 25569 45178
rect 22468 45067 22520 45076
rect 22468 45033 22477 45067
rect 22477 45033 22511 45067
rect 22511 45033 22520 45067
rect 22468 45024 22520 45033
rect 24768 45067 24820 45076
rect 24768 45033 24777 45067
rect 24777 45033 24811 45067
rect 24811 45033 24820 45067
rect 24768 45024 24820 45033
rect 24952 45024 25004 45076
rect 26240 45024 26292 45076
rect 27896 45024 27948 45076
rect 4804 44956 4856 45008
rect 23112 44956 23164 45008
rect 27804 44956 27856 45008
rect 25136 44888 25188 44940
rect 3056 44820 3108 44872
rect 3148 44820 3200 44872
rect 25964 44888 26016 44940
rect 28356 44931 28408 44940
rect 28356 44897 28365 44931
rect 28365 44897 28399 44931
rect 28399 44897 28408 44931
rect 28356 44888 28408 44897
rect 25872 44863 25924 44872
rect 25872 44829 25881 44863
rect 25881 44829 25915 44863
rect 25915 44829 25924 44863
rect 25872 44820 25924 44829
rect 27252 44752 27304 44804
rect 27804 44684 27856 44736
rect 7896 44582 7948 44634
rect 7960 44582 8012 44634
rect 8024 44582 8076 44634
rect 8088 44582 8140 44634
rect 8152 44582 8204 44634
rect 14842 44582 14894 44634
rect 14906 44582 14958 44634
rect 14970 44582 15022 44634
rect 15034 44582 15086 44634
rect 15098 44582 15150 44634
rect 21788 44582 21840 44634
rect 21852 44582 21904 44634
rect 21916 44582 21968 44634
rect 21980 44582 22032 44634
rect 22044 44582 22096 44634
rect 28734 44582 28786 44634
rect 28798 44582 28850 44634
rect 28862 44582 28914 44634
rect 28926 44582 28978 44634
rect 28990 44582 29042 44634
rect 27252 44523 27304 44532
rect 27252 44489 27261 44523
rect 27261 44489 27295 44523
rect 27295 44489 27304 44523
rect 27252 44480 27304 44489
rect 26424 44455 26476 44464
rect 26424 44421 26433 44455
rect 26433 44421 26467 44455
rect 26467 44421 26476 44455
rect 26424 44412 26476 44421
rect 2412 44344 2464 44396
rect 3148 44387 3200 44396
rect 3148 44353 3157 44387
rect 3157 44353 3191 44387
rect 3191 44353 3200 44387
rect 3148 44344 3200 44353
rect 26884 44344 26936 44396
rect 27344 44387 27396 44396
rect 27344 44353 27353 44387
rect 27353 44353 27387 44387
rect 27387 44353 27396 44387
rect 27344 44344 27396 44353
rect 27804 44387 27856 44396
rect 27804 44353 27813 44387
rect 27813 44353 27847 44387
rect 27847 44353 27856 44387
rect 27804 44344 27856 44353
rect 3332 44319 3384 44328
rect 3332 44285 3341 44319
rect 3341 44285 3375 44319
rect 3375 44285 3384 44319
rect 3332 44276 3384 44285
rect 3608 44319 3660 44328
rect 3608 44285 3617 44319
rect 3617 44285 3651 44319
rect 3651 44285 3660 44319
rect 3608 44276 3660 44285
rect 26056 44319 26108 44328
rect 26056 44285 26065 44319
rect 26065 44285 26099 44319
rect 26099 44285 26108 44319
rect 26056 44276 26108 44285
rect 27528 44276 27580 44328
rect 3608 44140 3660 44192
rect 4423 44038 4475 44090
rect 4487 44038 4539 44090
rect 4551 44038 4603 44090
rect 4615 44038 4667 44090
rect 4679 44038 4731 44090
rect 11369 44038 11421 44090
rect 11433 44038 11485 44090
rect 11497 44038 11549 44090
rect 11561 44038 11613 44090
rect 11625 44038 11677 44090
rect 18315 44038 18367 44090
rect 18379 44038 18431 44090
rect 18443 44038 18495 44090
rect 18507 44038 18559 44090
rect 18571 44038 18623 44090
rect 25261 44038 25313 44090
rect 25325 44038 25377 44090
rect 25389 44038 25441 44090
rect 25453 44038 25505 44090
rect 25517 44038 25569 44090
rect 3332 43936 3384 43988
rect 112 43800 164 43852
rect 3056 43800 3108 43852
rect 11888 43800 11940 43852
rect 25872 43843 25924 43852
rect 25872 43809 25881 43843
rect 25881 43809 25915 43843
rect 25915 43809 25924 43843
rect 25872 43800 25924 43809
rect 26148 43800 26200 43852
rect 4160 43775 4212 43784
rect 4160 43741 4169 43775
rect 4169 43741 4203 43775
rect 4203 43741 4212 43775
rect 4160 43732 4212 43741
rect 4620 43775 4672 43784
rect 4620 43741 4629 43775
rect 4629 43741 4663 43775
rect 4663 43741 4672 43775
rect 4620 43732 4672 43741
rect 27252 43732 27304 43784
rect 3240 43707 3292 43716
rect 3240 43673 3249 43707
rect 3249 43673 3283 43707
rect 3283 43673 3292 43707
rect 3240 43664 3292 43673
rect 26056 43707 26108 43716
rect 26056 43673 26065 43707
rect 26065 43673 26099 43707
rect 26099 43673 26108 43707
rect 26056 43664 26108 43673
rect 7896 43494 7948 43546
rect 7960 43494 8012 43546
rect 8024 43494 8076 43546
rect 8088 43494 8140 43546
rect 8152 43494 8204 43546
rect 14842 43494 14894 43546
rect 14906 43494 14958 43546
rect 14970 43494 15022 43546
rect 15034 43494 15086 43546
rect 15098 43494 15150 43546
rect 21788 43494 21840 43546
rect 21852 43494 21904 43546
rect 21916 43494 21968 43546
rect 21980 43494 22032 43546
rect 22044 43494 22096 43546
rect 28734 43494 28786 43546
rect 28798 43494 28850 43546
rect 28862 43494 28914 43546
rect 28926 43494 28978 43546
rect 28990 43494 29042 43546
rect 26056 43392 26108 43444
rect 20 43324 72 43376
rect 3608 43367 3660 43376
rect 3608 43333 3617 43367
rect 3617 43333 3651 43367
rect 3651 43333 3660 43367
rect 3608 43324 3660 43333
rect 4620 43256 4672 43308
rect 25780 43256 25832 43308
rect 27068 43256 27120 43308
rect 26976 43188 27028 43240
rect 27896 43256 27948 43308
rect 26424 43052 26476 43104
rect 28080 43095 28132 43104
rect 28080 43061 28089 43095
rect 28089 43061 28123 43095
rect 28123 43061 28132 43095
rect 28080 43052 28132 43061
rect 4423 42950 4475 43002
rect 4487 42950 4539 43002
rect 4551 42950 4603 43002
rect 4615 42950 4667 43002
rect 4679 42950 4731 43002
rect 11369 42950 11421 43002
rect 11433 42950 11485 43002
rect 11497 42950 11549 43002
rect 11561 42950 11613 43002
rect 11625 42950 11677 43002
rect 18315 42950 18367 43002
rect 18379 42950 18431 43002
rect 18443 42950 18495 43002
rect 18507 42950 18559 43002
rect 18571 42950 18623 43002
rect 25261 42950 25313 43002
rect 25325 42950 25377 43002
rect 25389 42950 25441 43002
rect 25453 42950 25505 43002
rect 25517 42950 25569 43002
rect 3240 42712 3292 42764
rect 28080 42712 28132 42764
rect 2412 42687 2464 42696
rect 2412 42653 2421 42687
rect 2421 42653 2455 42687
rect 2455 42653 2464 42687
rect 2412 42644 2464 42653
rect 3424 42576 3476 42628
rect 26148 42576 26200 42628
rect 27804 42576 27856 42628
rect 7896 42406 7948 42458
rect 7960 42406 8012 42458
rect 8024 42406 8076 42458
rect 8088 42406 8140 42458
rect 8152 42406 8204 42458
rect 14842 42406 14894 42458
rect 14906 42406 14958 42458
rect 14970 42406 15022 42458
rect 15034 42406 15086 42458
rect 15098 42406 15150 42458
rect 21788 42406 21840 42458
rect 21852 42406 21904 42458
rect 21916 42406 21968 42458
rect 21980 42406 22032 42458
rect 22044 42406 22096 42458
rect 28734 42406 28786 42458
rect 28798 42406 28850 42458
rect 28862 42406 28914 42458
rect 28926 42406 28978 42458
rect 28990 42406 29042 42458
rect 27804 42347 27856 42356
rect 27804 42313 27813 42347
rect 27813 42313 27847 42347
rect 27847 42313 27856 42347
rect 27804 42304 27856 42313
rect 26424 42279 26476 42288
rect 26424 42245 26433 42279
rect 26433 42245 26467 42279
rect 26467 42245 26476 42279
rect 26424 42236 26476 42245
rect 2504 42168 2556 42220
rect 27252 42168 27304 42220
rect 27620 42168 27672 42220
rect 26056 42143 26108 42152
rect 26056 42109 26065 42143
rect 26065 42109 26099 42143
rect 26099 42109 26108 42143
rect 26056 42100 26108 42109
rect 1676 41964 1728 42016
rect 3240 41964 3292 42016
rect 4423 41862 4475 41914
rect 4487 41862 4539 41914
rect 4551 41862 4603 41914
rect 4615 41862 4667 41914
rect 4679 41862 4731 41914
rect 11369 41862 11421 41914
rect 11433 41862 11485 41914
rect 11497 41862 11549 41914
rect 11561 41862 11613 41914
rect 11625 41862 11677 41914
rect 18315 41862 18367 41914
rect 18379 41862 18431 41914
rect 18443 41862 18495 41914
rect 18507 41862 18559 41914
rect 18571 41862 18623 41914
rect 25261 41862 25313 41914
rect 25325 41862 25377 41914
rect 25389 41862 25441 41914
rect 25453 41862 25505 41914
rect 25517 41862 25569 41914
rect 1584 41667 1636 41676
rect 1584 41633 1593 41667
rect 1593 41633 1627 41667
rect 1627 41633 1636 41667
rect 1584 41624 1636 41633
rect 3240 41667 3292 41676
rect 3240 41633 3249 41667
rect 3249 41633 3283 41667
rect 3283 41633 3292 41667
rect 3240 41624 3292 41633
rect 3424 41667 3476 41676
rect 3424 41633 3433 41667
rect 3433 41633 3467 41667
rect 3467 41633 3476 41667
rect 3424 41624 3476 41633
rect 27528 41667 27580 41676
rect 27528 41633 27537 41667
rect 27537 41633 27571 41667
rect 27571 41633 27580 41667
rect 27528 41624 27580 41633
rect 27344 41488 27396 41540
rect 27896 41420 27948 41472
rect 7896 41318 7948 41370
rect 7960 41318 8012 41370
rect 8024 41318 8076 41370
rect 8088 41318 8140 41370
rect 8152 41318 8204 41370
rect 14842 41318 14894 41370
rect 14906 41318 14958 41370
rect 14970 41318 15022 41370
rect 15034 41318 15086 41370
rect 15098 41318 15150 41370
rect 21788 41318 21840 41370
rect 21852 41318 21904 41370
rect 21916 41318 21968 41370
rect 21980 41318 22032 41370
rect 22044 41318 22096 41370
rect 28734 41318 28786 41370
rect 28798 41318 28850 41370
rect 28862 41318 28914 41370
rect 28926 41318 28978 41370
rect 28990 41318 29042 41370
rect 1676 41123 1728 41132
rect 1676 41089 1685 41123
rect 1685 41089 1719 41123
rect 1719 41089 1728 41123
rect 1676 41080 1728 41089
rect 27896 41123 27948 41132
rect 27896 41089 27905 41123
rect 27905 41089 27939 41123
rect 27939 41089 27948 41123
rect 27896 41080 27948 41089
rect 2228 41012 2280 41064
rect 2780 41055 2832 41064
rect 2780 41021 2789 41055
rect 2789 41021 2823 41055
rect 2823 41021 2832 41055
rect 2780 41012 2832 41021
rect 26516 40876 26568 40928
rect 4423 40774 4475 40826
rect 4487 40774 4539 40826
rect 4551 40774 4603 40826
rect 4615 40774 4667 40826
rect 4679 40774 4731 40826
rect 11369 40774 11421 40826
rect 11433 40774 11485 40826
rect 11497 40774 11549 40826
rect 11561 40774 11613 40826
rect 11625 40774 11677 40826
rect 18315 40774 18367 40826
rect 18379 40774 18431 40826
rect 18443 40774 18495 40826
rect 18507 40774 18559 40826
rect 18571 40774 18623 40826
rect 25261 40774 25313 40826
rect 25325 40774 25377 40826
rect 25389 40774 25441 40826
rect 25453 40774 25505 40826
rect 25517 40774 25569 40826
rect 2228 40715 2280 40724
rect 2228 40681 2237 40715
rect 2237 40681 2271 40715
rect 2271 40681 2280 40715
rect 2228 40672 2280 40681
rect 26516 40579 26568 40588
rect 26516 40545 26525 40579
rect 26525 40545 26559 40579
rect 26559 40545 26568 40579
rect 26516 40536 26568 40545
rect 28632 40536 28684 40588
rect 2320 40511 2372 40520
rect 2320 40477 2329 40511
rect 2329 40477 2363 40511
rect 2363 40477 2372 40511
rect 2320 40468 2372 40477
rect 26700 40443 26752 40452
rect 26700 40409 26709 40443
rect 26709 40409 26743 40443
rect 26743 40409 26752 40443
rect 26700 40400 26752 40409
rect 7896 40230 7948 40282
rect 7960 40230 8012 40282
rect 8024 40230 8076 40282
rect 8088 40230 8140 40282
rect 8152 40230 8204 40282
rect 14842 40230 14894 40282
rect 14906 40230 14958 40282
rect 14970 40230 15022 40282
rect 15034 40230 15086 40282
rect 15098 40230 15150 40282
rect 21788 40230 21840 40282
rect 21852 40230 21904 40282
rect 21916 40230 21968 40282
rect 21980 40230 22032 40282
rect 22044 40230 22096 40282
rect 28734 40230 28786 40282
rect 28798 40230 28850 40282
rect 28862 40230 28914 40282
rect 28926 40230 28978 40282
rect 28990 40230 29042 40282
rect 27344 40035 27396 40044
rect 27344 40001 27353 40035
rect 27353 40001 27387 40035
rect 27387 40001 27396 40035
rect 27344 39992 27396 40001
rect 26976 39924 27028 39976
rect 1676 39788 1728 39840
rect 27896 39831 27948 39840
rect 27896 39797 27905 39831
rect 27905 39797 27939 39831
rect 27939 39797 27948 39831
rect 27896 39788 27948 39797
rect 4423 39686 4475 39738
rect 4487 39686 4539 39738
rect 4551 39686 4603 39738
rect 4615 39686 4667 39738
rect 4679 39686 4731 39738
rect 11369 39686 11421 39738
rect 11433 39686 11485 39738
rect 11497 39686 11549 39738
rect 11561 39686 11613 39738
rect 11625 39686 11677 39738
rect 18315 39686 18367 39738
rect 18379 39686 18431 39738
rect 18443 39686 18495 39738
rect 18507 39686 18559 39738
rect 18571 39686 18623 39738
rect 25261 39686 25313 39738
rect 25325 39686 25377 39738
rect 25389 39686 25441 39738
rect 25453 39686 25505 39738
rect 25517 39686 25569 39738
rect 27896 39448 27948 39500
rect 29920 39448 29972 39500
rect 2780 39380 2832 39432
rect 3240 39423 3292 39432
rect 3240 39389 3249 39423
rect 3249 39389 3283 39423
rect 3283 39389 3292 39423
rect 3240 39380 3292 39389
rect 4344 39312 4396 39364
rect 1768 39244 1820 39296
rect 2964 39244 3016 39296
rect 26424 39312 26476 39364
rect 26332 39244 26384 39296
rect 7896 39142 7948 39194
rect 7960 39142 8012 39194
rect 8024 39142 8076 39194
rect 8088 39142 8140 39194
rect 8152 39142 8204 39194
rect 14842 39142 14894 39194
rect 14906 39142 14958 39194
rect 14970 39142 15022 39194
rect 15034 39142 15086 39194
rect 15098 39142 15150 39194
rect 21788 39142 21840 39194
rect 21852 39142 21904 39194
rect 21916 39142 21968 39194
rect 21980 39142 22032 39194
rect 22044 39142 22096 39194
rect 28734 39142 28786 39194
rect 28798 39142 28850 39194
rect 28862 39142 28914 39194
rect 28926 39142 28978 39194
rect 28990 39142 29042 39194
rect 2964 39015 3016 39024
rect 2964 38981 2973 39015
rect 2973 38981 3007 39015
rect 3007 38981 3016 39015
rect 2964 38972 3016 38981
rect 2780 38947 2832 38956
rect 2780 38913 2789 38947
rect 2789 38913 2823 38947
rect 2823 38913 2832 38947
rect 2780 38904 2832 38913
rect 18972 38947 19024 38956
rect 18972 38913 18981 38947
rect 18981 38913 19015 38947
rect 19015 38913 19024 38947
rect 18972 38904 19024 38913
rect 20076 38947 20128 38956
rect 4252 38879 4304 38888
rect 4252 38845 4261 38879
rect 4261 38845 4295 38879
rect 4295 38845 4304 38879
rect 4252 38836 4304 38845
rect 20076 38913 20085 38947
rect 20085 38913 20119 38947
rect 20119 38913 20128 38947
rect 20076 38904 20128 38913
rect 20720 38947 20772 38956
rect 20720 38913 20729 38947
rect 20729 38913 20763 38947
rect 20763 38913 20772 38947
rect 20720 38904 20772 38913
rect 26700 39040 26752 39092
rect 20536 38836 20588 38888
rect 21640 38836 21692 38888
rect 2872 38768 2924 38820
rect 19708 38768 19760 38820
rect 20076 38768 20128 38820
rect 26332 38904 26384 38956
rect 27344 38947 27396 38956
rect 27344 38913 27353 38947
rect 27353 38913 27387 38947
rect 27387 38913 27396 38947
rect 27344 38904 27396 38913
rect 21824 38768 21876 38820
rect 26516 38768 26568 38820
rect 1584 38743 1636 38752
rect 1584 38709 1593 38743
rect 1593 38709 1627 38743
rect 1627 38709 1636 38743
rect 1584 38700 1636 38709
rect 19616 38743 19668 38752
rect 19616 38709 19625 38743
rect 19625 38709 19659 38743
rect 19659 38709 19668 38743
rect 19616 38700 19668 38709
rect 20352 38700 20404 38752
rect 21272 38743 21324 38752
rect 21272 38709 21281 38743
rect 21281 38709 21315 38743
rect 21315 38709 21324 38743
rect 21272 38700 21324 38709
rect 26700 38700 26752 38752
rect 4423 38598 4475 38650
rect 4487 38598 4539 38650
rect 4551 38598 4603 38650
rect 4615 38598 4667 38650
rect 4679 38598 4731 38650
rect 11369 38598 11421 38650
rect 11433 38598 11485 38650
rect 11497 38598 11549 38650
rect 11561 38598 11613 38650
rect 11625 38598 11677 38650
rect 18315 38598 18367 38650
rect 18379 38598 18431 38650
rect 18443 38598 18495 38650
rect 18507 38598 18559 38650
rect 18571 38598 18623 38650
rect 25261 38598 25313 38650
rect 25325 38598 25377 38650
rect 25389 38598 25441 38650
rect 25453 38598 25505 38650
rect 25517 38598 25569 38650
rect 18696 38539 18748 38548
rect 18696 38505 18705 38539
rect 18705 38505 18739 38539
rect 18739 38505 18748 38539
rect 18696 38496 18748 38505
rect 18972 38496 19024 38548
rect 1676 38428 1728 38480
rect 1768 38403 1820 38412
rect 1768 38369 1777 38403
rect 1777 38369 1811 38403
rect 1811 38369 1820 38403
rect 1768 38360 1820 38369
rect 2780 38403 2832 38412
rect 2780 38369 2789 38403
rect 2789 38369 2823 38403
rect 2823 38369 2832 38403
rect 2780 38360 2832 38369
rect 18052 38224 18104 38276
rect 19616 38224 19668 38276
rect 20720 38496 20772 38548
rect 26424 38496 26476 38548
rect 20076 38428 20128 38480
rect 26516 38403 26568 38412
rect 26516 38369 26525 38403
rect 26525 38369 26559 38403
rect 26559 38369 26568 38403
rect 26516 38360 26568 38369
rect 26700 38403 26752 38412
rect 26700 38369 26709 38403
rect 26709 38369 26743 38403
rect 26743 38369 26752 38403
rect 26700 38360 26752 38369
rect 28632 38360 28684 38412
rect 21824 38335 21876 38344
rect 21824 38301 21833 38335
rect 21833 38301 21867 38335
rect 21867 38301 21876 38335
rect 21824 38292 21876 38301
rect 21272 38224 21324 38276
rect 21640 38224 21692 38276
rect 26884 38224 26936 38276
rect 20444 38156 20496 38208
rect 21364 38199 21416 38208
rect 21364 38165 21373 38199
rect 21373 38165 21407 38199
rect 21407 38165 21416 38199
rect 21364 38156 21416 38165
rect 7896 38054 7948 38106
rect 7960 38054 8012 38106
rect 8024 38054 8076 38106
rect 8088 38054 8140 38106
rect 8152 38054 8204 38106
rect 14842 38054 14894 38106
rect 14906 38054 14958 38106
rect 14970 38054 15022 38106
rect 15034 38054 15086 38106
rect 15098 38054 15150 38106
rect 21788 38054 21840 38106
rect 21852 38054 21904 38106
rect 21916 38054 21968 38106
rect 21980 38054 22032 38106
rect 22044 38054 22096 38106
rect 28734 38054 28786 38106
rect 28798 38054 28850 38106
rect 28862 38054 28914 38106
rect 28926 38054 28978 38106
rect 28990 38054 29042 38106
rect 20720 37952 20772 38004
rect 20812 37952 20864 38004
rect 19616 37884 19668 37936
rect 20996 37884 21048 37936
rect 1676 37791 1728 37800
rect 1676 37757 1685 37791
rect 1685 37757 1719 37791
rect 1719 37757 1728 37791
rect 1676 37748 1728 37757
rect 2780 37748 2832 37800
rect 18696 37816 18748 37868
rect 19064 37859 19116 37868
rect 19064 37825 19073 37859
rect 19073 37825 19107 37859
rect 19107 37825 19116 37859
rect 19064 37816 19116 37825
rect 19984 37816 20036 37868
rect 21364 37816 21416 37868
rect 27344 37859 27396 37868
rect 27344 37825 27353 37859
rect 27353 37825 27387 37859
rect 27387 37825 27396 37859
rect 27344 37816 27396 37825
rect 27988 37816 28040 37868
rect 21640 37748 21692 37800
rect 27712 37791 27764 37800
rect 27712 37757 27721 37791
rect 27721 37757 27755 37791
rect 27755 37757 27764 37791
rect 27712 37748 27764 37757
rect 20536 37680 20588 37732
rect 20720 37680 20772 37732
rect 18236 37612 18288 37664
rect 20076 37612 20128 37664
rect 22376 37612 22428 37664
rect 4423 37510 4475 37562
rect 4487 37510 4539 37562
rect 4551 37510 4603 37562
rect 4615 37510 4667 37562
rect 4679 37510 4731 37562
rect 11369 37510 11421 37562
rect 11433 37510 11485 37562
rect 11497 37510 11549 37562
rect 11561 37510 11613 37562
rect 11625 37510 11677 37562
rect 18315 37510 18367 37562
rect 18379 37510 18431 37562
rect 18443 37510 18495 37562
rect 18507 37510 18559 37562
rect 18571 37510 18623 37562
rect 25261 37510 25313 37562
rect 25325 37510 25377 37562
rect 25389 37510 25441 37562
rect 25453 37510 25505 37562
rect 25517 37510 25569 37562
rect 18236 37451 18288 37460
rect 18236 37417 18245 37451
rect 18245 37417 18279 37451
rect 18279 37417 18288 37451
rect 18236 37408 18288 37417
rect 19340 37408 19392 37460
rect 19616 37451 19668 37460
rect 19616 37417 19625 37451
rect 19625 37417 19659 37451
rect 19659 37417 19668 37451
rect 19616 37408 19668 37417
rect 20444 37451 20496 37460
rect 20444 37417 20453 37451
rect 20453 37417 20487 37451
rect 20487 37417 20496 37451
rect 20444 37408 20496 37417
rect 1492 37204 1544 37256
rect 16856 37315 16908 37324
rect 16856 37281 16865 37315
rect 16865 37281 16899 37315
rect 16899 37281 16908 37315
rect 16856 37272 16908 37281
rect 19064 37340 19116 37392
rect 20812 37340 20864 37392
rect 19524 37272 19576 37324
rect 21364 37272 21416 37324
rect 2780 37204 2832 37256
rect 2688 37136 2740 37188
rect 6000 37204 6052 37256
rect 19984 37247 20036 37256
rect 4344 37136 4396 37188
rect 15292 37136 15344 37188
rect 17960 37136 18012 37188
rect 18052 37179 18104 37188
rect 18052 37145 18061 37179
rect 18061 37145 18095 37179
rect 18095 37145 18104 37179
rect 19984 37213 19993 37247
rect 19993 37213 20027 37247
rect 20027 37213 20036 37247
rect 19984 37204 20036 37213
rect 20720 37204 20772 37256
rect 20996 37204 21048 37256
rect 28356 37247 28408 37256
rect 28356 37213 28365 37247
rect 28365 37213 28399 37247
rect 28399 37213 28408 37247
rect 28356 37204 28408 37213
rect 18052 37136 18104 37145
rect 17408 37111 17460 37120
rect 17408 37077 17417 37111
rect 17417 37077 17451 37111
rect 17451 37077 17460 37111
rect 17408 37068 17460 37077
rect 18420 37111 18472 37120
rect 18420 37077 18429 37111
rect 18429 37077 18463 37111
rect 18463 37077 18472 37111
rect 18420 37068 18472 37077
rect 26148 37136 26200 37188
rect 27896 37136 27948 37188
rect 20812 37111 20864 37120
rect 20812 37077 20821 37111
rect 20821 37077 20855 37111
rect 20855 37077 20864 37111
rect 20812 37068 20864 37077
rect 7896 36966 7948 37018
rect 7960 36966 8012 37018
rect 8024 36966 8076 37018
rect 8088 36966 8140 37018
rect 8152 36966 8204 37018
rect 14842 36966 14894 37018
rect 14906 36966 14958 37018
rect 14970 36966 15022 37018
rect 15034 36966 15086 37018
rect 15098 36966 15150 37018
rect 21788 36966 21840 37018
rect 21852 36966 21904 37018
rect 21916 36966 21968 37018
rect 21980 36966 22032 37018
rect 22044 36966 22096 37018
rect 28734 36966 28786 37018
rect 28798 36966 28850 37018
rect 28862 36966 28914 37018
rect 28926 36966 28978 37018
rect 28990 36966 29042 37018
rect 15752 36864 15804 36916
rect 18052 36864 18104 36916
rect 21364 36907 21416 36916
rect 21364 36873 21373 36907
rect 21373 36873 21407 36907
rect 21407 36873 21416 36907
rect 21364 36864 21416 36873
rect 27896 36907 27948 36916
rect 27896 36873 27905 36907
rect 27905 36873 27939 36907
rect 27939 36873 27948 36907
rect 27896 36864 27948 36873
rect 4344 36796 4396 36848
rect 19432 36796 19484 36848
rect 2596 36771 2648 36780
rect 2596 36737 2605 36771
rect 2605 36737 2639 36771
rect 2639 36737 2648 36771
rect 2596 36728 2648 36737
rect 17408 36728 17460 36780
rect 18420 36771 18472 36780
rect 18420 36737 18429 36771
rect 18429 36737 18463 36771
rect 18463 36737 18472 36771
rect 18420 36728 18472 36737
rect 21456 36771 21508 36780
rect 21456 36737 21465 36771
rect 21465 36737 21499 36771
rect 21499 36737 21508 36771
rect 21456 36728 21508 36737
rect 24860 36728 24912 36780
rect 2136 36660 2188 36712
rect 2412 36703 2464 36712
rect 2412 36669 2421 36703
rect 2421 36669 2455 36703
rect 2455 36669 2464 36703
rect 2412 36660 2464 36669
rect 4160 36660 4212 36712
rect 9588 36660 9640 36712
rect 16672 36660 16724 36712
rect 27344 36771 27396 36780
rect 27344 36737 27353 36771
rect 27353 36737 27387 36771
rect 27387 36737 27396 36771
rect 27344 36728 27396 36737
rect 27804 36771 27856 36780
rect 27804 36737 27813 36771
rect 27813 36737 27847 36771
rect 27847 36737 27856 36771
rect 27804 36728 27856 36737
rect 10692 36524 10744 36576
rect 17776 36524 17828 36576
rect 18788 36524 18840 36576
rect 20812 36524 20864 36576
rect 24676 36524 24728 36576
rect 24768 36524 24820 36576
rect 4423 36422 4475 36474
rect 4487 36422 4539 36474
rect 4551 36422 4603 36474
rect 4615 36422 4667 36474
rect 4679 36422 4731 36474
rect 11369 36422 11421 36474
rect 11433 36422 11485 36474
rect 11497 36422 11549 36474
rect 11561 36422 11613 36474
rect 11625 36422 11677 36474
rect 18315 36422 18367 36474
rect 18379 36422 18431 36474
rect 18443 36422 18495 36474
rect 18507 36422 18559 36474
rect 18571 36422 18623 36474
rect 25261 36422 25313 36474
rect 25325 36422 25377 36474
rect 25389 36422 25441 36474
rect 25453 36422 25505 36474
rect 25517 36422 25569 36474
rect 20720 36320 20772 36372
rect 28356 36320 28408 36372
rect 3516 36184 3568 36236
rect 4252 36184 4304 36236
rect 4804 36227 4856 36236
rect 4804 36193 4813 36227
rect 4813 36193 4847 36227
rect 4847 36193 4856 36227
rect 4804 36184 4856 36193
rect 15660 36184 15712 36236
rect 16856 36184 16908 36236
rect 23572 36227 23624 36236
rect 2412 36159 2464 36168
rect 2412 36125 2421 36159
rect 2421 36125 2455 36159
rect 2455 36125 2464 36159
rect 2412 36116 2464 36125
rect 2596 36116 2648 36168
rect 3976 36159 4028 36168
rect 3976 36125 3985 36159
rect 3985 36125 4019 36159
rect 4019 36125 4028 36159
rect 3976 36116 4028 36125
rect 16580 36116 16632 36168
rect 17776 36159 17828 36168
rect 17776 36125 17785 36159
rect 17785 36125 17819 36159
rect 17819 36125 17828 36159
rect 17776 36116 17828 36125
rect 20076 36159 20128 36168
rect 20076 36125 20085 36159
rect 20085 36125 20119 36159
rect 20119 36125 20128 36159
rect 20076 36116 20128 36125
rect 2964 36048 3016 36100
rect 3240 36091 3292 36100
rect 3240 36057 3249 36091
rect 3249 36057 3283 36091
rect 3283 36057 3292 36091
rect 3240 36048 3292 36057
rect 5908 36091 5960 36100
rect 5908 36057 5917 36091
rect 5917 36057 5951 36091
rect 5951 36057 5960 36091
rect 5908 36048 5960 36057
rect 9588 36048 9640 36100
rect 9772 36048 9824 36100
rect 14464 36048 14516 36100
rect 18236 36048 18288 36100
rect 23572 36193 23581 36227
rect 23581 36193 23615 36227
rect 23615 36193 23624 36227
rect 23572 36184 23624 36193
rect 20352 36159 20404 36168
rect 20352 36125 20386 36159
rect 20386 36125 20404 36159
rect 20352 36116 20404 36125
rect 23480 36116 23532 36168
rect 24492 36184 24544 36236
rect 24768 36227 24820 36236
rect 24768 36193 24777 36227
rect 24777 36193 24811 36227
rect 24811 36193 24820 36227
rect 24768 36184 24820 36193
rect 27436 36227 27488 36236
rect 27436 36193 27445 36227
rect 27445 36193 27479 36227
rect 27479 36193 27488 36227
rect 27436 36184 27488 36193
rect 25780 36159 25832 36168
rect 25780 36125 25789 36159
rect 25789 36125 25823 36159
rect 25823 36125 25832 36159
rect 25780 36116 25832 36125
rect 26240 36048 26292 36100
rect 6736 35980 6788 36032
rect 16488 36023 16540 36032
rect 16488 35989 16497 36023
rect 16497 35989 16531 36023
rect 16531 35989 16540 36023
rect 16488 35980 16540 35989
rect 17132 36023 17184 36032
rect 17132 35989 17141 36023
rect 17141 35989 17175 36023
rect 17175 35989 17184 36023
rect 17132 35980 17184 35989
rect 17592 36023 17644 36032
rect 17592 35989 17601 36023
rect 17601 35989 17635 36023
rect 17635 35989 17644 36023
rect 17592 35980 17644 35989
rect 18144 35980 18196 36032
rect 19340 35980 19392 36032
rect 22652 35980 22704 36032
rect 23112 36023 23164 36032
rect 23112 35989 23121 36023
rect 23121 35989 23155 36023
rect 23155 35989 23164 36023
rect 23112 35980 23164 35989
rect 23756 35980 23808 36032
rect 25688 35980 25740 36032
rect 7896 35878 7948 35930
rect 7960 35878 8012 35930
rect 8024 35878 8076 35930
rect 8088 35878 8140 35930
rect 8152 35878 8204 35930
rect 14842 35878 14894 35930
rect 14906 35878 14958 35930
rect 14970 35878 15022 35930
rect 15034 35878 15086 35930
rect 15098 35878 15150 35930
rect 21788 35878 21840 35930
rect 21852 35878 21904 35930
rect 21916 35878 21968 35930
rect 21980 35878 22032 35930
rect 22044 35878 22096 35930
rect 28734 35878 28786 35930
rect 28798 35878 28850 35930
rect 28862 35878 28914 35930
rect 28926 35878 28978 35930
rect 28990 35878 29042 35930
rect 1676 35751 1728 35760
rect 1676 35717 1685 35751
rect 1685 35717 1719 35751
rect 1719 35717 1728 35751
rect 1676 35708 1728 35717
rect 5908 35708 5960 35760
rect 16580 35708 16632 35760
rect 17132 35751 17184 35760
rect 17132 35717 17166 35751
rect 17166 35717 17184 35751
rect 17132 35708 17184 35717
rect 3516 35683 3568 35692
rect 3516 35649 3525 35683
rect 3525 35649 3559 35683
rect 3559 35649 3568 35683
rect 3976 35683 4028 35692
rect 3516 35640 3568 35649
rect 3976 35649 3985 35683
rect 3985 35649 4019 35683
rect 4019 35649 4028 35683
rect 3976 35640 4028 35649
rect 7748 35640 7800 35692
rect 16488 35640 16540 35692
rect 20076 35708 20128 35760
rect 18788 35640 18840 35692
rect 22468 35640 22520 35692
rect 22652 35683 22704 35692
rect 22652 35649 22686 35683
rect 22686 35649 22704 35683
rect 22652 35640 22704 35649
rect 24860 35708 24912 35760
rect 24768 35640 24820 35692
rect 26240 35819 26292 35828
rect 26240 35785 26249 35819
rect 26249 35785 26283 35819
rect 26283 35785 26292 35819
rect 26240 35776 26292 35785
rect 26700 35640 26752 35692
rect 3056 35572 3108 35624
rect 4344 35615 4396 35624
rect 4344 35581 4353 35615
rect 4353 35581 4387 35615
rect 4387 35581 4396 35615
rect 4344 35572 4396 35581
rect 16672 35572 16724 35624
rect 16856 35615 16908 35624
rect 16856 35581 16865 35615
rect 16865 35581 16899 35615
rect 16899 35581 16908 35615
rect 16856 35572 16908 35581
rect 18236 35547 18288 35556
rect 18236 35513 18245 35547
rect 18245 35513 18279 35547
rect 18279 35513 18288 35547
rect 18236 35504 18288 35513
rect 19616 35436 19668 35488
rect 23756 35479 23808 35488
rect 23756 35445 23765 35479
rect 23765 35445 23799 35479
rect 23799 35445 23808 35479
rect 23756 35436 23808 35445
rect 24124 35436 24176 35488
rect 26240 35436 26292 35488
rect 26516 35436 26568 35488
rect 4423 35334 4475 35386
rect 4487 35334 4539 35386
rect 4551 35334 4603 35386
rect 4615 35334 4667 35386
rect 4679 35334 4731 35386
rect 11369 35334 11421 35386
rect 11433 35334 11485 35386
rect 11497 35334 11549 35386
rect 11561 35334 11613 35386
rect 11625 35334 11677 35386
rect 18315 35334 18367 35386
rect 18379 35334 18431 35386
rect 18443 35334 18495 35386
rect 18507 35334 18559 35386
rect 18571 35334 18623 35386
rect 25261 35334 25313 35386
rect 25325 35334 25377 35386
rect 25389 35334 25441 35386
rect 25453 35334 25505 35386
rect 25517 35334 25569 35386
rect 3056 35275 3108 35284
rect 3056 35241 3065 35275
rect 3065 35241 3099 35275
rect 3099 35241 3108 35275
rect 3056 35232 3108 35241
rect 20536 35232 20588 35284
rect 21640 35232 21692 35284
rect 23480 35275 23532 35284
rect 23480 35241 23489 35275
rect 23489 35241 23523 35275
rect 23523 35241 23532 35275
rect 23480 35232 23532 35241
rect 24768 35275 24820 35284
rect 24768 35241 24777 35275
rect 24777 35241 24811 35275
rect 24811 35241 24820 35275
rect 24768 35232 24820 35241
rect 25780 35232 25832 35284
rect 2412 35139 2464 35148
rect 2412 35105 2421 35139
rect 2421 35105 2455 35139
rect 2455 35105 2464 35139
rect 2412 35096 2464 35105
rect 1584 35071 1636 35080
rect 1584 35037 1593 35071
rect 1593 35037 1627 35071
rect 1627 35037 1636 35071
rect 1584 35028 1636 35037
rect 3884 35028 3936 35080
rect 5908 35028 5960 35080
rect 16856 35071 16908 35080
rect 16856 35037 16865 35071
rect 16865 35037 16899 35071
rect 16899 35037 16908 35071
rect 16856 35028 16908 35037
rect 20076 35028 20128 35080
rect 22376 35071 22428 35080
rect 22376 35037 22394 35071
rect 22394 35037 22428 35071
rect 22376 35028 22428 35037
rect 22560 35028 22612 35080
rect 23112 35071 23164 35080
rect 23112 35037 23121 35071
rect 23121 35037 23155 35071
rect 23155 35037 23164 35071
rect 23112 35028 23164 35037
rect 17592 34960 17644 35012
rect 19708 35003 19760 35012
rect 19708 34969 19742 35003
rect 19742 34969 19760 35003
rect 19708 34960 19760 34969
rect 22744 34960 22796 35012
rect 24124 34960 24176 35012
rect 24952 35028 25004 35080
rect 25964 35096 26016 35148
rect 26516 35139 26568 35148
rect 26516 35105 26525 35139
rect 26525 35105 26559 35139
rect 26559 35105 26568 35139
rect 26516 35096 26568 35105
rect 27528 35139 27580 35148
rect 27528 35105 27537 35139
rect 27537 35105 27571 35139
rect 27571 35105 27580 35139
rect 27528 35096 27580 35105
rect 17960 34892 18012 34944
rect 18880 34892 18932 34944
rect 27896 34892 27948 34944
rect 7896 34790 7948 34842
rect 7960 34790 8012 34842
rect 8024 34790 8076 34842
rect 8088 34790 8140 34842
rect 8152 34790 8204 34842
rect 14842 34790 14894 34842
rect 14906 34790 14958 34842
rect 14970 34790 15022 34842
rect 15034 34790 15086 34842
rect 15098 34790 15150 34842
rect 21788 34790 21840 34842
rect 21852 34790 21904 34842
rect 21916 34790 21968 34842
rect 21980 34790 22032 34842
rect 22044 34790 22096 34842
rect 28734 34790 28786 34842
rect 28798 34790 28850 34842
rect 28862 34790 28914 34842
rect 28926 34790 28978 34842
rect 28990 34790 29042 34842
rect 19340 34688 19392 34740
rect 26608 34731 26660 34740
rect 26608 34697 26617 34731
rect 26617 34697 26651 34731
rect 26651 34697 26660 34731
rect 26608 34688 26660 34697
rect 14740 34620 14792 34672
rect 24952 34620 25004 34672
rect 25688 34620 25740 34672
rect 19616 34552 19668 34604
rect 24860 34552 24912 34604
rect 1676 34527 1728 34536
rect 1676 34493 1685 34527
rect 1685 34493 1719 34527
rect 1719 34493 1728 34527
rect 1676 34484 1728 34493
rect 1860 34527 1912 34536
rect 1860 34493 1869 34527
rect 1869 34493 1903 34527
rect 1903 34493 1912 34527
rect 1860 34484 1912 34493
rect 2780 34527 2832 34536
rect 2780 34493 2789 34527
rect 2789 34493 2823 34527
rect 2823 34493 2832 34527
rect 2780 34484 2832 34493
rect 16672 34484 16724 34536
rect 19708 34484 19760 34536
rect 27160 34391 27212 34400
rect 27160 34357 27169 34391
rect 27169 34357 27203 34391
rect 27203 34357 27212 34391
rect 27160 34348 27212 34357
rect 4423 34246 4475 34298
rect 4487 34246 4539 34298
rect 4551 34246 4603 34298
rect 4615 34246 4667 34298
rect 4679 34246 4731 34298
rect 11369 34246 11421 34298
rect 11433 34246 11485 34298
rect 11497 34246 11549 34298
rect 11561 34246 11613 34298
rect 11625 34246 11677 34298
rect 18315 34246 18367 34298
rect 18379 34246 18431 34298
rect 18443 34246 18495 34298
rect 18507 34246 18559 34298
rect 18571 34246 18623 34298
rect 25261 34246 25313 34298
rect 25325 34246 25377 34298
rect 25389 34246 25441 34298
rect 25453 34246 25505 34298
rect 25517 34246 25569 34298
rect 1860 34144 1912 34196
rect 21456 34144 21508 34196
rect 26148 34076 26200 34128
rect 2320 33940 2372 33992
rect 4344 33940 4396 33992
rect 22468 33983 22520 33992
rect 22468 33949 22477 33983
rect 22477 33949 22511 33983
rect 22511 33949 22520 33983
rect 22468 33940 22520 33949
rect 23756 33940 23808 33992
rect 24676 33983 24728 33992
rect 24676 33949 24685 33983
rect 24685 33949 24719 33983
rect 24719 33949 24728 33983
rect 24676 33940 24728 33949
rect 26608 34008 26660 34060
rect 22192 33915 22244 33924
rect 22192 33881 22210 33915
rect 22210 33881 22244 33915
rect 22192 33872 22244 33881
rect 27252 33872 27304 33924
rect 20720 33804 20772 33856
rect 24952 33804 25004 33856
rect 26240 33804 26292 33856
rect 7896 33702 7948 33754
rect 7960 33702 8012 33754
rect 8024 33702 8076 33754
rect 8088 33702 8140 33754
rect 8152 33702 8204 33754
rect 14842 33702 14894 33754
rect 14906 33702 14958 33754
rect 14970 33702 15022 33754
rect 15034 33702 15086 33754
rect 15098 33702 15150 33754
rect 21788 33702 21840 33754
rect 21852 33702 21904 33754
rect 21916 33702 21968 33754
rect 21980 33702 22032 33754
rect 22044 33702 22096 33754
rect 28734 33702 28786 33754
rect 28798 33702 28850 33754
rect 28862 33702 28914 33754
rect 28926 33702 28978 33754
rect 28990 33702 29042 33754
rect 18696 33532 18748 33584
rect 19432 33532 19484 33584
rect 1676 33464 1728 33516
rect 17960 33507 18012 33516
rect 17960 33473 17969 33507
rect 17969 33473 18003 33507
rect 18003 33473 18012 33507
rect 17960 33464 18012 33473
rect 18144 33464 18196 33516
rect 18880 33464 18932 33516
rect 20904 33600 20956 33652
rect 21640 33600 21692 33652
rect 22192 33643 22244 33652
rect 22192 33609 22201 33643
rect 22201 33609 22235 33643
rect 22235 33609 22244 33643
rect 22192 33600 22244 33609
rect 27252 33643 27304 33652
rect 27252 33609 27261 33643
rect 27261 33609 27295 33643
rect 27295 33609 27304 33643
rect 27252 33600 27304 33609
rect 20720 33532 20772 33584
rect 24860 33532 24912 33584
rect 20444 33507 20496 33516
rect 20444 33473 20453 33507
rect 20453 33473 20487 33507
rect 20487 33473 20496 33507
rect 20444 33464 20496 33473
rect 19984 33396 20036 33448
rect 22284 33464 22336 33516
rect 23388 33507 23440 33516
rect 23388 33473 23397 33507
rect 23397 33473 23431 33507
rect 23431 33473 23440 33507
rect 23388 33464 23440 33473
rect 24032 33507 24084 33516
rect 24032 33473 24041 33507
rect 24041 33473 24075 33507
rect 24075 33473 24084 33507
rect 24032 33464 24084 33473
rect 26884 33464 26936 33516
rect 28172 33464 28224 33516
rect 27160 33396 27212 33448
rect 3516 33328 3568 33380
rect 9128 33328 9180 33380
rect 16764 33328 16816 33380
rect 18972 33328 19024 33380
rect 26700 33328 26752 33380
rect 26884 33328 26936 33380
rect 18144 33260 18196 33312
rect 19340 33303 19392 33312
rect 19340 33269 19349 33303
rect 19349 33269 19383 33303
rect 19383 33269 19392 33303
rect 19340 33260 19392 33269
rect 21916 33260 21968 33312
rect 23204 33303 23256 33312
rect 23204 33269 23213 33303
rect 23213 33269 23247 33303
rect 23247 33269 23256 33303
rect 23204 33260 23256 33269
rect 25044 33260 25096 33312
rect 28264 33260 28316 33312
rect 4423 33158 4475 33210
rect 4487 33158 4539 33210
rect 4551 33158 4603 33210
rect 4615 33158 4667 33210
rect 4679 33158 4731 33210
rect 11369 33158 11421 33210
rect 11433 33158 11485 33210
rect 11497 33158 11549 33210
rect 11561 33158 11613 33210
rect 11625 33158 11677 33210
rect 18315 33158 18367 33210
rect 18379 33158 18431 33210
rect 18443 33158 18495 33210
rect 18507 33158 18559 33210
rect 18571 33158 18623 33210
rect 25261 33158 25313 33210
rect 25325 33158 25377 33210
rect 25389 33158 25441 33210
rect 25453 33158 25505 33210
rect 25517 33158 25569 33210
rect 17868 33056 17920 33108
rect 17960 33056 18012 33108
rect 18236 33056 18288 33108
rect 19432 33099 19484 33108
rect 19432 33065 19441 33099
rect 19441 33065 19475 33099
rect 19475 33065 19484 33099
rect 19432 33056 19484 33065
rect 19892 33056 19944 33108
rect 20444 33056 20496 33108
rect 20720 33099 20772 33108
rect 20720 33065 20729 33099
rect 20729 33065 20763 33099
rect 20763 33065 20772 33099
rect 20720 33056 20772 33065
rect 24032 33099 24084 33108
rect 1676 32895 1728 32904
rect 1676 32861 1685 32895
rect 1685 32861 1719 32895
rect 1719 32861 1728 32895
rect 1676 32852 1728 32861
rect 15292 32895 15344 32904
rect 15292 32861 15301 32895
rect 15301 32861 15335 32895
rect 15335 32861 15344 32895
rect 15292 32852 15344 32861
rect 16764 32988 16816 33040
rect 16212 32963 16264 32972
rect 16212 32929 16221 32963
rect 16221 32929 16255 32963
rect 16255 32929 16264 32963
rect 16212 32920 16264 32929
rect 16764 32852 16816 32904
rect 18788 32988 18840 33040
rect 18696 32920 18748 32972
rect 19892 32963 19944 32972
rect 19892 32929 19901 32963
rect 19901 32929 19935 32963
rect 19935 32929 19944 32963
rect 19892 32920 19944 32929
rect 18052 32895 18104 32904
rect 15936 32827 15988 32836
rect 15936 32793 15945 32827
rect 15945 32793 15979 32827
rect 15979 32793 15988 32827
rect 15936 32784 15988 32793
rect 18052 32861 18061 32895
rect 18061 32861 18095 32895
rect 18095 32861 18104 32895
rect 18052 32852 18104 32861
rect 18328 32852 18380 32904
rect 19616 32895 19668 32904
rect 19616 32861 19625 32895
rect 19625 32861 19659 32895
rect 19659 32861 19668 32895
rect 19616 32852 19668 32861
rect 19800 32895 19852 32904
rect 19800 32861 19809 32895
rect 19809 32861 19843 32895
rect 19843 32861 19852 32895
rect 19800 32852 19852 32861
rect 19984 32895 20036 32904
rect 19984 32861 19993 32895
rect 19993 32861 20027 32895
rect 20027 32861 20036 32895
rect 19984 32852 20036 32861
rect 20352 32988 20404 33040
rect 20904 32988 20956 33040
rect 20812 32852 20864 32904
rect 24032 33065 24041 33099
rect 24041 33065 24075 33099
rect 24075 33065 24084 33099
rect 24032 33056 24084 33065
rect 24676 32988 24728 33040
rect 25136 32963 25188 32972
rect 25136 32929 25145 32963
rect 25145 32929 25179 32963
rect 25179 32929 25188 32963
rect 25136 32920 25188 32929
rect 27528 32963 27580 32972
rect 27528 32929 27537 32963
rect 27537 32929 27571 32963
rect 27571 32929 27580 32963
rect 27528 32920 27580 32929
rect 21916 32895 21968 32904
rect 21916 32861 21925 32895
rect 21925 32861 21959 32895
rect 21959 32861 21968 32895
rect 21916 32852 21968 32861
rect 22192 32852 22244 32904
rect 22468 32852 22520 32904
rect 23204 32852 23256 32904
rect 24860 32895 24912 32904
rect 24860 32861 24869 32895
rect 24869 32861 24903 32895
rect 24903 32861 24912 32895
rect 24860 32852 24912 32861
rect 25044 32852 25096 32904
rect 26516 32895 26568 32904
rect 26516 32861 26525 32895
rect 26525 32861 26559 32895
rect 26559 32861 26568 32895
rect 26516 32852 26568 32861
rect 15476 32759 15528 32768
rect 15476 32725 15485 32759
rect 15485 32725 15519 32759
rect 15519 32725 15528 32759
rect 15476 32716 15528 32725
rect 16580 32716 16632 32768
rect 18972 32784 19024 32836
rect 19156 32784 19208 32836
rect 28080 32784 28132 32836
rect 18052 32716 18104 32768
rect 20536 32716 20588 32768
rect 24676 32759 24728 32768
rect 24676 32725 24685 32759
rect 24685 32725 24719 32759
rect 24719 32725 24728 32759
rect 24676 32716 24728 32725
rect 7896 32614 7948 32666
rect 7960 32614 8012 32666
rect 8024 32614 8076 32666
rect 8088 32614 8140 32666
rect 8152 32614 8204 32666
rect 14842 32614 14894 32666
rect 14906 32614 14958 32666
rect 14970 32614 15022 32666
rect 15034 32614 15086 32666
rect 15098 32614 15150 32666
rect 21788 32614 21840 32666
rect 21852 32614 21904 32666
rect 21916 32614 21968 32666
rect 21980 32614 22032 32666
rect 22044 32614 22096 32666
rect 28734 32614 28786 32666
rect 28798 32614 28850 32666
rect 28862 32614 28914 32666
rect 28926 32614 28978 32666
rect 28990 32614 29042 32666
rect 15476 32512 15528 32564
rect 16212 32512 16264 32564
rect 20536 32555 20588 32564
rect 15292 32487 15344 32496
rect 15292 32453 15301 32487
rect 15301 32453 15335 32487
rect 15335 32453 15344 32487
rect 15292 32444 15344 32453
rect 15752 32487 15804 32496
rect 15752 32453 15761 32487
rect 15761 32453 15795 32487
rect 15795 32453 15804 32487
rect 15752 32444 15804 32453
rect 20536 32521 20545 32555
rect 20545 32521 20579 32555
rect 20579 32521 20588 32555
rect 20536 32512 20588 32521
rect 24032 32512 24084 32564
rect 28080 32555 28132 32564
rect 28080 32521 28089 32555
rect 28089 32521 28123 32555
rect 28123 32521 28132 32555
rect 28080 32512 28132 32521
rect 19156 32487 19208 32496
rect 19156 32453 19165 32487
rect 19165 32453 19199 32487
rect 19199 32453 19208 32487
rect 19156 32444 19208 32453
rect 1676 32419 1728 32428
rect 1676 32385 1685 32419
rect 1685 32385 1719 32419
rect 1719 32385 1728 32419
rect 1676 32376 1728 32385
rect 2044 32308 2096 32360
rect 2780 32351 2832 32360
rect 2780 32317 2789 32351
rect 2789 32317 2823 32351
rect 2823 32317 2832 32351
rect 2780 32308 2832 32317
rect 15936 32308 15988 32360
rect 18052 32419 18104 32428
rect 18052 32385 18061 32419
rect 18061 32385 18095 32419
rect 18095 32385 18104 32419
rect 18052 32376 18104 32385
rect 18144 32419 18196 32428
rect 18144 32385 18153 32419
rect 18153 32385 18187 32419
rect 18187 32385 18196 32419
rect 18144 32376 18196 32385
rect 19340 32376 19392 32428
rect 18696 32308 18748 32360
rect 18788 32351 18840 32360
rect 18788 32317 18797 32351
rect 18797 32317 18831 32351
rect 18831 32317 18840 32351
rect 20076 32419 20128 32428
rect 20076 32385 20085 32419
rect 20085 32385 20119 32419
rect 20119 32385 20128 32419
rect 20812 32444 20864 32496
rect 26424 32444 26476 32496
rect 20076 32376 20128 32385
rect 20352 32419 20404 32428
rect 20352 32385 20361 32419
rect 20361 32385 20395 32419
rect 20395 32385 20404 32419
rect 20352 32376 20404 32385
rect 22100 32376 22152 32428
rect 22652 32376 22704 32428
rect 26516 32376 26568 32428
rect 27068 32376 27120 32428
rect 27988 32419 28040 32428
rect 27988 32385 27997 32419
rect 27997 32385 28031 32419
rect 28031 32385 28040 32419
rect 27988 32376 28040 32385
rect 18788 32308 18840 32317
rect 20168 32308 20220 32360
rect 20996 32308 21048 32360
rect 24492 32351 24544 32360
rect 24492 32317 24501 32351
rect 24501 32317 24535 32351
rect 24535 32317 24544 32351
rect 24492 32308 24544 32317
rect 15844 32172 15896 32224
rect 17040 32215 17092 32224
rect 17040 32181 17049 32215
rect 17049 32181 17083 32215
rect 17083 32181 17092 32215
rect 17040 32172 17092 32181
rect 19064 32172 19116 32224
rect 21640 32172 21692 32224
rect 23480 32172 23532 32224
rect 23664 32172 23716 32224
rect 26700 32172 26752 32224
rect 4423 32070 4475 32122
rect 4487 32070 4539 32122
rect 4551 32070 4603 32122
rect 4615 32070 4667 32122
rect 4679 32070 4731 32122
rect 11369 32070 11421 32122
rect 11433 32070 11485 32122
rect 11497 32070 11549 32122
rect 11561 32070 11613 32122
rect 11625 32070 11677 32122
rect 18315 32070 18367 32122
rect 18379 32070 18431 32122
rect 18443 32070 18495 32122
rect 18507 32070 18559 32122
rect 18571 32070 18623 32122
rect 25261 32070 25313 32122
rect 25325 32070 25377 32122
rect 25389 32070 25441 32122
rect 25453 32070 25505 32122
rect 25517 32070 25569 32122
rect 2044 32011 2096 32020
rect 2044 31977 2053 32011
rect 2053 31977 2087 32011
rect 2087 31977 2096 32011
rect 2044 31968 2096 31977
rect 15936 31968 15988 32020
rect 18236 31968 18288 32020
rect 19800 31968 19852 32020
rect 20904 31968 20956 32020
rect 22284 31968 22336 32020
rect 23388 31968 23440 32020
rect 16580 31832 16632 31884
rect 16856 31832 16908 31884
rect 22744 31832 22796 31884
rect 25872 31900 25924 31952
rect 27712 31900 27764 31952
rect 26700 31875 26752 31884
rect 2596 31764 2648 31816
rect 4160 31764 4212 31816
rect 15292 31764 15344 31816
rect 17040 31764 17092 31816
rect 18880 31764 18932 31816
rect 20904 31764 20956 31816
rect 21548 31807 21600 31816
rect 21548 31773 21557 31807
rect 21557 31773 21591 31807
rect 21591 31773 21600 31807
rect 21548 31764 21600 31773
rect 21640 31764 21692 31816
rect 26700 31841 26709 31875
rect 26709 31841 26743 31875
rect 26743 31841 26752 31875
rect 26700 31832 26752 31841
rect 28356 31875 28408 31884
rect 28356 31841 28365 31875
rect 28365 31841 28399 31875
rect 28399 31841 28408 31875
rect 28356 31832 28408 31841
rect 23664 31807 23716 31816
rect 23664 31773 23673 31807
rect 23673 31773 23707 31807
rect 23707 31773 23716 31807
rect 23664 31764 23716 31773
rect 25136 31764 25188 31816
rect 25596 31739 25648 31748
rect 25596 31705 25605 31739
rect 25605 31705 25639 31739
rect 25639 31705 25648 31739
rect 25596 31696 25648 31705
rect 16028 31628 16080 31680
rect 18328 31671 18380 31680
rect 18328 31637 18337 31671
rect 18337 31637 18371 31671
rect 18371 31637 18380 31671
rect 18328 31628 18380 31637
rect 26332 31764 26384 31816
rect 26516 31628 26568 31680
rect 7896 31526 7948 31578
rect 7960 31526 8012 31578
rect 8024 31526 8076 31578
rect 8088 31526 8140 31578
rect 8152 31526 8204 31578
rect 14842 31526 14894 31578
rect 14906 31526 14958 31578
rect 14970 31526 15022 31578
rect 15034 31526 15086 31578
rect 15098 31526 15150 31578
rect 21788 31526 21840 31578
rect 21852 31526 21904 31578
rect 21916 31526 21968 31578
rect 21980 31526 22032 31578
rect 22044 31526 22096 31578
rect 28734 31526 28786 31578
rect 28798 31526 28850 31578
rect 28862 31526 28914 31578
rect 28926 31526 28978 31578
rect 28990 31526 29042 31578
rect 18236 31424 18288 31476
rect 22652 31467 22704 31476
rect 22652 31433 22661 31467
rect 22661 31433 22695 31467
rect 22695 31433 22704 31467
rect 22652 31424 22704 31433
rect 25044 31424 25096 31476
rect 25596 31356 25648 31408
rect 15844 31331 15896 31340
rect 15844 31297 15853 31331
rect 15853 31297 15887 31331
rect 15887 31297 15896 31331
rect 15844 31288 15896 31297
rect 16580 31288 16632 31340
rect 17868 31288 17920 31340
rect 18328 31331 18380 31340
rect 18328 31297 18337 31331
rect 18337 31297 18371 31331
rect 18371 31297 18380 31331
rect 18328 31288 18380 31297
rect 22652 31288 22704 31340
rect 23480 31288 23532 31340
rect 24400 31331 24452 31340
rect 24400 31297 24409 31331
rect 24409 31297 24443 31331
rect 24443 31297 24452 31331
rect 24400 31288 24452 31297
rect 26056 31288 26108 31340
rect 26516 31288 26568 31340
rect 27712 31288 27764 31340
rect 28356 31288 28408 31340
rect 24492 31220 24544 31272
rect 27344 31263 27396 31272
rect 15936 31127 15988 31136
rect 15936 31093 15945 31127
rect 15945 31093 15979 31127
rect 15979 31093 15988 31127
rect 15936 31084 15988 31093
rect 25596 31084 25648 31136
rect 25964 31084 26016 31136
rect 27344 31229 27353 31263
rect 27353 31229 27387 31263
rect 27387 31229 27396 31263
rect 27344 31220 27396 31229
rect 26700 31084 26752 31136
rect 28172 31084 28224 31136
rect 4423 30982 4475 31034
rect 4487 30982 4539 31034
rect 4551 30982 4603 31034
rect 4615 30982 4667 31034
rect 4679 30982 4731 31034
rect 11369 30982 11421 31034
rect 11433 30982 11485 31034
rect 11497 30982 11549 31034
rect 11561 30982 11613 31034
rect 11625 30982 11677 31034
rect 18315 30982 18367 31034
rect 18379 30982 18431 31034
rect 18443 30982 18495 31034
rect 18507 30982 18559 31034
rect 18571 30982 18623 31034
rect 25261 30982 25313 31034
rect 25325 30982 25377 31034
rect 25389 30982 25441 31034
rect 25453 30982 25505 31034
rect 25517 30982 25569 31034
rect 16028 30923 16080 30932
rect 16028 30889 16037 30923
rect 16037 30889 16071 30923
rect 16071 30889 16080 30923
rect 16028 30880 16080 30889
rect 17868 30923 17920 30932
rect 17868 30889 17877 30923
rect 17877 30889 17911 30923
rect 17911 30889 17920 30923
rect 17868 30880 17920 30889
rect 25136 30880 25188 30932
rect 26056 30923 26108 30932
rect 26056 30889 26065 30923
rect 26065 30889 26099 30923
rect 26099 30889 26108 30923
rect 26056 30880 26108 30889
rect 2136 30812 2188 30864
rect 28356 30880 28408 30932
rect 28264 30812 28316 30864
rect 27436 30787 27488 30796
rect 27436 30753 27445 30787
rect 27445 30753 27479 30787
rect 27479 30753 27488 30787
rect 27436 30744 27488 30753
rect 28172 30787 28224 30796
rect 28172 30753 28181 30787
rect 28181 30753 28215 30787
rect 28215 30753 28224 30787
rect 28172 30744 28224 30753
rect 9128 30719 9180 30728
rect 9128 30685 9137 30719
rect 9137 30685 9171 30719
rect 9171 30685 9180 30719
rect 9128 30676 9180 30685
rect 12624 30676 12676 30728
rect 17960 30719 18012 30728
rect 17960 30685 17969 30719
rect 17969 30685 18003 30719
rect 18003 30685 18012 30719
rect 17960 30676 18012 30685
rect 24860 30719 24912 30728
rect 24860 30685 24869 30719
rect 24869 30685 24903 30719
rect 24903 30685 24912 30719
rect 24860 30676 24912 30685
rect 25044 30719 25096 30728
rect 25044 30685 25053 30719
rect 25053 30685 25087 30719
rect 25087 30685 25096 30719
rect 25044 30676 25096 30685
rect 25872 30719 25924 30728
rect 9588 30608 9640 30660
rect 9956 30608 10008 30660
rect 15844 30651 15896 30660
rect 15844 30617 15853 30651
rect 15853 30617 15887 30651
rect 15887 30617 15896 30651
rect 15844 30608 15896 30617
rect 15936 30608 15988 30660
rect 22560 30651 22612 30660
rect 22560 30617 22569 30651
rect 22569 30617 22603 30651
rect 22603 30617 22612 30651
rect 22560 30608 22612 30617
rect 24400 30608 24452 30660
rect 25872 30685 25881 30719
rect 25881 30685 25915 30719
rect 25915 30685 25924 30719
rect 25872 30676 25924 30685
rect 26700 30676 26752 30728
rect 25780 30608 25832 30660
rect 16212 30583 16264 30592
rect 16212 30549 16221 30583
rect 16221 30549 16255 30583
rect 16255 30549 16264 30583
rect 16212 30540 16264 30549
rect 22192 30540 22244 30592
rect 7896 30438 7948 30490
rect 7960 30438 8012 30490
rect 8024 30438 8076 30490
rect 8088 30438 8140 30490
rect 8152 30438 8204 30490
rect 14842 30438 14894 30490
rect 14906 30438 14958 30490
rect 14970 30438 15022 30490
rect 15034 30438 15086 30490
rect 15098 30438 15150 30490
rect 21788 30438 21840 30490
rect 21852 30438 21904 30490
rect 21916 30438 21968 30490
rect 21980 30438 22032 30490
rect 22044 30438 22096 30490
rect 28734 30438 28786 30490
rect 28798 30438 28850 30490
rect 28862 30438 28914 30490
rect 28926 30438 28978 30490
rect 28990 30438 29042 30490
rect 17960 30336 18012 30388
rect 20536 30268 20588 30320
rect 1584 30243 1636 30252
rect 1584 30209 1593 30243
rect 1593 30209 1627 30243
rect 1627 30209 1636 30243
rect 1584 30200 1636 30209
rect 16212 30200 16264 30252
rect 16856 30243 16908 30252
rect 16856 30209 16865 30243
rect 16865 30209 16899 30243
rect 16899 30209 16908 30243
rect 16856 30200 16908 30209
rect 21180 30268 21232 30320
rect 22652 30268 22704 30320
rect 20168 30175 20220 30184
rect 20168 30141 20177 30175
rect 20177 30141 20211 30175
rect 20211 30141 20220 30175
rect 20168 30132 20220 30141
rect 20996 30243 21048 30252
rect 20996 30209 21005 30243
rect 21005 30209 21039 30243
rect 21039 30209 21048 30243
rect 20996 30200 21048 30209
rect 26608 30243 26660 30252
rect 26608 30209 26617 30243
rect 26617 30209 26651 30243
rect 26651 30209 26660 30243
rect 26608 30200 26660 30209
rect 22376 30132 22428 30184
rect 24584 30132 24636 30184
rect 26424 30107 26476 30116
rect 26424 30073 26433 30107
rect 26433 30073 26467 30107
rect 26467 30073 26476 30107
rect 26424 30064 26476 30073
rect 1860 29996 1912 30048
rect 19616 29996 19668 30048
rect 20812 29996 20864 30048
rect 28356 29996 28408 30048
rect 4423 29894 4475 29946
rect 4487 29894 4539 29946
rect 4551 29894 4603 29946
rect 4615 29894 4667 29946
rect 4679 29894 4731 29946
rect 11369 29894 11421 29946
rect 11433 29894 11485 29946
rect 11497 29894 11549 29946
rect 11561 29894 11613 29946
rect 11625 29894 11677 29946
rect 18315 29894 18367 29946
rect 18379 29894 18431 29946
rect 18443 29894 18495 29946
rect 18507 29894 18559 29946
rect 18571 29894 18623 29946
rect 25261 29894 25313 29946
rect 25325 29894 25377 29946
rect 25389 29894 25441 29946
rect 25453 29894 25505 29946
rect 25517 29894 25569 29946
rect 16764 29792 16816 29844
rect 18236 29792 18288 29844
rect 18788 29792 18840 29844
rect 25596 29792 25648 29844
rect 26056 29792 26108 29844
rect 15936 29588 15988 29640
rect 16672 29656 16724 29708
rect 18052 29656 18104 29708
rect 16580 29631 16632 29640
rect 16580 29597 16589 29631
rect 16589 29597 16623 29631
rect 16623 29597 16632 29631
rect 16580 29588 16632 29597
rect 18144 29588 18196 29640
rect 19524 29656 19576 29708
rect 20812 29699 20864 29708
rect 20812 29665 20821 29699
rect 20821 29665 20855 29699
rect 20855 29665 20864 29699
rect 20812 29656 20864 29665
rect 22652 29699 22704 29708
rect 22652 29665 22661 29699
rect 22661 29665 22695 29699
rect 22695 29665 22704 29699
rect 22652 29656 22704 29665
rect 19616 29631 19668 29640
rect 19616 29597 19625 29631
rect 19625 29597 19659 29631
rect 19659 29597 19668 29631
rect 19616 29588 19668 29597
rect 21180 29588 21232 29640
rect 22836 29631 22888 29640
rect 22836 29597 22845 29631
rect 22845 29597 22879 29631
rect 22879 29597 22888 29631
rect 22836 29588 22888 29597
rect 27528 29699 27580 29708
rect 27528 29665 27537 29699
rect 27537 29665 27571 29699
rect 27571 29665 27580 29699
rect 27528 29656 27580 29665
rect 28356 29699 28408 29708
rect 28356 29665 28365 29699
rect 28365 29665 28399 29699
rect 28399 29665 28408 29699
rect 28356 29656 28408 29665
rect 23940 29588 23992 29640
rect 23480 29520 23532 29572
rect 24860 29520 24912 29572
rect 15752 29452 15804 29504
rect 16764 29495 16816 29504
rect 16764 29461 16773 29495
rect 16773 29461 16807 29495
rect 16807 29461 16816 29495
rect 16764 29452 16816 29461
rect 19524 29495 19576 29504
rect 19524 29461 19533 29495
rect 19533 29461 19567 29495
rect 19567 29461 19576 29495
rect 19524 29452 19576 29461
rect 20904 29452 20956 29504
rect 22928 29495 22980 29504
rect 22928 29461 22937 29495
rect 22937 29461 22971 29495
rect 22971 29461 22980 29495
rect 22928 29452 22980 29461
rect 24952 29495 25004 29504
rect 24952 29461 24961 29495
rect 24961 29461 24995 29495
rect 24995 29461 25004 29495
rect 24952 29452 25004 29461
rect 26148 29520 26200 29572
rect 27712 29520 27764 29572
rect 25872 29452 25924 29504
rect 7896 29350 7948 29402
rect 7960 29350 8012 29402
rect 8024 29350 8076 29402
rect 8088 29350 8140 29402
rect 8152 29350 8204 29402
rect 14842 29350 14894 29402
rect 14906 29350 14958 29402
rect 14970 29350 15022 29402
rect 15034 29350 15086 29402
rect 15098 29350 15150 29402
rect 21788 29350 21840 29402
rect 21852 29350 21904 29402
rect 21916 29350 21968 29402
rect 21980 29350 22032 29402
rect 22044 29350 22096 29402
rect 28734 29350 28786 29402
rect 28798 29350 28850 29402
rect 28862 29350 28914 29402
rect 28926 29350 28978 29402
rect 28990 29350 29042 29402
rect 20996 29248 21048 29300
rect 22836 29248 22888 29300
rect 27712 29291 27764 29300
rect 27712 29257 27721 29291
rect 27721 29257 27755 29291
rect 27755 29257 27764 29291
rect 27712 29248 27764 29257
rect 22560 29180 22612 29232
rect 15936 29112 15988 29164
rect 16672 29112 16724 29164
rect 20904 29112 20956 29164
rect 21088 29155 21140 29164
rect 21088 29121 21097 29155
rect 21097 29121 21131 29155
rect 21131 29121 21140 29155
rect 21088 29112 21140 29121
rect 22100 29155 22152 29164
rect 22100 29121 22109 29155
rect 22109 29121 22143 29155
rect 22143 29121 22152 29155
rect 22100 29112 22152 29121
rect 22928 29112 22980 29164
rect 23480 29112 23532 29164
rect 24584 29155 24636 29164
rect 16856 29044 16908 29096
rect 19432 29044 19484 29096
rect 21640 29044 21692 29096
rect 24032 29044 24084 29096
rect 24584 29121 24593 29155
rect 24593 29121 24627 29155
rect 24627 29121 24636 29155
rect 24584 29112 24636 29121
rect 24952 29180 25004 29232
rect 26148 29223 26200 29232
rect 26148 29189 26157 29223
rect 26157 29189 26191 29223
rect 26191 29189 26200 29223
rect 26148 29180 26200 29189
rect 25872 29155 25924 29164
rect 25872 29121 25881 29155
rect 25881 29121 25915 29155
rect 25915 29121 25924 29155
rect 25872 29112 25924 29121
rect 26056 29112 26108 29164
rect 25136 29044 25188 29096
rect 23480 29019 23532 29028
rect 15936 28951 15988 28960
rect 15936 28917 15945 28951
rect 15945 28917 15979 28951
rect 15979 28917 15988 28951
rect 15936 28908 15988 28917
rect 23480 28985 23489 29019
rect 23489 28985 23523 29019
rect 23523 28985 23532 29019
rect 23480 28976 23532 28985
rect 27896 29112 27948 29164
rect 22284 28908 22336 28960
rect 25596 28908 25648 28960
rect 26240 28908 26292 28960
rect 4423 28806 4475 28858
rect 4487 28806 4539 28858
rect 4551 28806 4603 28858
rect 4615 28806 4667 28858
rect 4679 28806 4731 28858
rect 11369 28806 11421 28858
rect 11433 28806 11485 28858
rect 11497 28806 11549 28858
rect 11561 28806 11613 28858
rect 11625 28806 11677 28858
rect 18315 28806 18367 28858
rect 18379 28806 18431 28858
rect 18443 28806 18495 28858
rect 18507 28806 18559 28858
rect 18571 28806 18623 28858
rect 25261 28806 25313 28858
rect 25325 28806 25377 28858
rect 25389 28806 25441 28858
rect 25453 28806 25505 28858
rect 25517 28806 25569 28858
rect 15844 28704 15896 28756
rect 16580 28704 16632 28756
rect 18236 28747 18288 28756
rect 18236 28713 18245 28747
rect 18245 28713 18279 28747
rect 18279 28713 18288 28747
rect 18236 28704 18288 28713
rect 20168 28704 20220 28756
rect 21548 28704 21600 28756
rect 24584 28704 24636 28756
rect 25136 28747 25188 28756
rect 25136 28713 25145 28747
rect 25145 28713 25179 28747
rect 25179 28713 25188 28747
rect 25136 28704 25188 28713
rect 16672 28636 16724 28688
rect 16856 28611 16908 28620
rect 16856 28577 16865 28611
rect 16865 28577 16899 28611
rect 16899 28577 16908 28611
rect 16856 28568 16908 28577
rect 19432 28611 19484 28620
rect 19432 28577 19441 28611
rect 19441 28577 19475 28611
rect 19475 28577 19484 28611
rect 19432 28568 19484 28577
rect 22100 28568 22152 28620
rect 25964 28568 26016 28620
rect 15752 28543 15804 28552
rect 15752 28509 15761 28543
rect 15761 28509 15795 28543
rect 15795 28509 15804 28543
rect 15752 28500 15804 28509
rect 16764 28500 16816 28552
rect 19524 28500 19576 28552
rect 20536 28500 20588 28552
rect 23664 28543 23716 28552
rect 23664 28509 23673 28543
rect 23673 28509 23707 28543
rect 23707 28509 23716 28543
rect 23664 28500 23716 28509
rect 23848 28500 23900 28552
rect 24676 28500 24728 28552
rect 15936 28432 15988 28484
rect 23388 28432 23440 28484
rect 24400 28432 24452 28484
rect 24952 28543 25004 28552
rect 24952 28509 24961 28543
rect 24961 28509 24995 28543
rect 24995 28509 25004 28543
rect 24952 28500 25004 28509
rect 25596 28500 25648 28552
rect 25044 28432 25096 28484
rect 26148 28432 26200 28484
rect 18236 28364 18288 28416
rect 19064 28364 19116 28416
rect 25688 28364 25740 28416
rect 26056 28364 26108 28416
rect 7896 28262 7948 28314
rect 7960 28262 8012 28314
rect 8024 28262 8076 28314
rect 8088 28262 8140 28314
rect 8152 28262 8204 28314
rect 14842 28262 14894 28314
rect 14906 28262 14958 28314
rect 14970 28262 15022 28314
rect 15034 28262 15086 28314
rect 15098 28262 15150 28314
rect 21788 28262 21840 28314
rect 21852 28262 21904 28314
rect 21916 28262 21968 28314
rect 21980 28262 22032 28314
rect 22044 28262 22096 28314
rect 28734 28262 28786 28314
rect 28798 28262 28850 28314
rect 28862 28262 28914 28314
rect 28926 28262 28978 28314
rect 28990 28262 29042 28314
rect 20352 28160 20404 28212
rect 24492 28203 24544 28212
rect 24492 28169 24501 28203
rect 24501 28169 24535 28203
rect 24535 28169 24544 28203
rect 24492 28160 24544 28169
rect 26148 28203 26200 28212
rect 26148 28169 26157 28203
rect 26157 28169 26191 28203
rect 26191 28169 26200 28203
rect 26148 28160 26200 28169
rect 18236 28135 18288 28144
rect 18236 28101 18245 28135
rect 18245 28101 18279 28135
rect 18279 28101 18288 28135
rect 18236 28092 18288 28101
rect 1584 28067 1636 28076
rect 1584 28033 1593 28067
rect 1593 28033 1627 28067
rect 1627 28033 1636 28067
rect 1584 28024 1636 28033
rect 21088 28092 21140 28144
rect 25044 28092 25096 28144
rect 18880 28067 18932 28076
rect 18880 28033 18889 28067
rect 18889 28033 18923 28067
rect 18923 28033 18932 28067
rect 19064 28067 19116 28076
rect 18880 28024 18932 28033
rect 19064 28033 19073 28067
rect 19073 28033 19107 28067
rect 19107 28033 19116 28067
rect 19064 28024 19116 28033
rect 19156 28067 19208 28076
rect 19156 28033 19165 28067
rect 19165 28033 19199 28067
rect 19199 28033 19208 28067
rect 19892 28067 19944 28076
rect 19156 28024 19208 28033
rect 19892 28033 19901 28067
rect 19901 28033 19935 28067
rect 19935 28033 19944 28067
rect 19892 28024 19944 28033
rect 23388 28067 23440 28076
rect 23388 28033 23397 28067
rect 23397 28033 23431 28067
rect 23431 28033 23440 28067
rect 23388 28024 23440 28033
rect 23480 28024 23532 28076
rect 18880 27888 18932 27940
rect 23664 27888 23716 27940
rect 25136 28024 25188 28076
rect 25688 28067 25740 28076
rect 25688 28033 25697 28067
rect 25697 28033 25731 28067
rect 25731 28033 25740 28067
rect 25688 28024 25740 28033
rect 26516 28092 26568 28144
rect 26056 28024 26108 28076
rect 26608 27956 26660 28008
rect 26148 27888 26200 27940
rect 1768 27863 1820 27872
rect 1768 27829 1777 27863
rect 1777 27829 1811 27863
rect 1811 27829 1820 27863
rect 1768 27820 1820 27829
rect 18788 27820 18840 27872
rect 20536 27820 20588 27872
rect 23020 27820 23072 27872
rect 24860 27820 24912 27872
rect 25688 27820 25740 27872
rect 28172 27863 28224 27872
rect 28172 27829 28181 27863
rect 28181 27829 28215 27863
rect 28215 27829 28224 27863
rect 28172 27820 28224 27829
rect 4423 27718 4475 27770
rect 4487 27718 4539 27770
rect 4551 27718 4603 27770
rect 4615 27718 4667 27770
rect 4679 27718 4731 27770
rect 11369 27718 11421 27770
rect 11433 27718 11485 27770
rect 11497 27718 11549 27770
rect 11561 27718 11613 27770
rect 11625 27718 11677 27770
rect 18315 27718 18367 27770
rect 18379 27718 18431 27770
rect 18443 27718 18495 27770
rect 18507 27718 18559 27770
rect 18571 27718 18623 27770
rect 25261 27718 25313 27770
rect 25325 27718 25377 27770
rect 25389 27718 25441 27770
rect 25453 27718 25505 27770
rect 25517 27718 25569 27770
rect 24952 27616 25004 27668
rect 18052 27591 18104 27600
rect 18052 27557 18061 27591
rect 18061 27557 18095 27591
rect 18095 27557 18104 27591
rect 18052 27548 18104 27557
rect 21456 27548 21508 27600
rect 15384 27523 15436 27532
rect 15384 27489 15393 27523
rect 15393 27489 15427 27523
rect 15427 27489 15436 27523
rect 15384 27480 15436 27489
rect 16764 27412 16816 27464
rect 19432 27480 19484 27532
rect 27528 27523 27580 27532
rect 27528 27489 27537 27523
rect 27537 27489 27571 27523
rect 27571 27489 27580 27523
rect 27528 27480 27580 27489
rect 28172 27480 28224 27532
rect 1768 27344 1820 27396
rect 18788 27412 18840 27464
rect 23020 27412 23072 27464
rect 23848 27455 23900 27464
rect 23848 27421 23857 27455
rect 23857 27421 23891 27455
rect 23891 27421 23900 27455
rect 23848 27412 23900 27421
rect 24032 27455 24084 27464
rect 24032 27421 24041 27455
rect 24041 27421 24075 27455
rect 24075 27421 24084 27455
rect 24032 27412 24084 27421
rect 24860 27412 24912 27464
rect 17040 27344 17092 27396
rect 20812 27344 20864 27396
rect 22376 27344 22428 27396
rect 15660 27276 15712 27328
rect 21364 27319 21416 27328
rect 21364 27285 21373 27319
rect 21373 27285 21407 27319
rect 21407 27285 21416 27319
rect 21364 27276 21416 27285
rect 23940 27319 23992 27328
rect 23940 27285 23949 27319
rect 23949 27285 23983 27319
rect 23983 27285 23992 27319
rect 23940 27276 23992 27285
rect 25872 27412 25924 27464
rect 25688 27344 25740 27396
rect 27896 27344 27948 27396
rect 25596 27276 25648 27328
rect 7896 27174 7948 27226
rect 7960 27174 8012 27226
rect 8024 27174 8076 27226
rect 8088 27174 8140 27226
rect 8152 27174 8204 27226
rect 14842 27174 14894 27226
rect 14906 27174 14958 27226
rect 14970 27174 15022 27226
rect 15034 27174 15086 27226
rect 15098 27174 15150 27226
rect 21788 27174 21840 27226
rect 21852 27174 21904 27226
rect 21916 27174 21968 27226
rect 21980 27174 22032 27226
rect 22044 27174 22096 27226
rect 28734 27174 28786 27226
rect 28798 27174 28850 27226
rect 28862 27174 28914 27226
rect 28926 27174 28978 27226
rect 28990 27174 29042 27226
rect 17040 27115 17092 27124
rect 17040 27081 17049 27115
rect 17049 27081 17083 27115
rect 17083 27081 17092 27115
rect 17040 27072 17092 27081
rect 15660 27004 15712 27056
rect 16212 27004 16264 27056
rect 20720 27072 20772 27124
rect 22468 27072 22520 27124
rect 25872 27115 25924 27124
rect 25872 27081 25881 27115
rect 25881 27081 25915 27115
rect 25915 27081 25924 27115
rect 25872 27072 25924 27081
rect 27896 27115 27948 27124
rect 27896 27081 27905 27115
rect 27905 27081 27939 27115
rect 27939 27081 27948 27115
rect 27896 27072 27948 27081
rect 22284 27004 22336 27056
rect 22744 27004 22796 27056
rect 18788 26979 18840 26988
rect 18788 26945 18797 26979
rect 18797 26945 18831 26979
rect 18831 26945 18840 26979
rect 18788 26936 18840 26945
rect 20996 26936 21048 26988
rect 21180 26936 21232 26988
rect 21456 26979 21508 26988
rect 21456 26945 21465 26979
rect 21465 26945 21499 26979
rect 21499 26945 21508 26979
rect 21456 26936 21508 26945
rect 26148 26979 26200 26988
rect 26148 26945 26157 26979
rect 26157 26945 26191 26979
rect 26191 26945 26200 26979
rect 26148 26936 26200 26945
rect 27620 26936 27672 26988
rect 26056 26868 26108 26920
rect 21548 26800 21600 26852
rect 17040 26732 17092 26784
rect 21732 26732 21784 26784
rect 26608 26800 26660 26852
rect 26516 26732 26568 26784
rect 4423 26630 4475 26682
rect 4487 26630 4539 26682
rect 4551 26630 4603 26682
rect 4615 26630 4667 26682
rect 4679 26630 4731 26682
rect 11369 26630 11421 26682
rect 11433 26630 11485 26682
rect 11497 26630 11549 26682
rect 11561 26630 11613 26682
rect 11625 26630 11677 26682
rect 18315 26630 18367 26682
rect 18379 26630 18431 26682
rect 18443 26630 18495 26682
rect 18507 26630 18559 26682
rect 18571 26630 18623 26682
rect 25261 26630 25313 26682
rect 25325 26630 25377 26682
rect 25389 26630 25441 26682
rect 25453 26630 25505 26682
rect 25517 26630 25569 26682
rect 20076 26528 20128 26580
rect 16672 26460 16724 26512
rect 17408 26460 17460 26512
rect 21364 26392 21416 26444
rect 22192 26528 22244 26580
rect 23388 26528 23440 26580
rect 26516 26435 26568 26444
rect 26516 26401 26525 26435
rect 26525 26401 26559 26435
rect 26559 26401 26568 26435
rect 26516 26392 26568 26401
rect 28356 26435 28408 26444
rect 28356 26401 28365 26435
rect 28365 26401 28399 26435
rect 28399 26401 28408 26435
rect 28356 26392 28408 26401
rect 1676 26324 1728 26376
rect 17040 26324 17092 26376
rect 19432 26367 19484 26376
rect 19432 26333 19441 26367
rect 19441 26333 19475 26367
rect 19475 26333 19484 26367
rect 19432 26324 19484 26333
rect 21548 26324 21600 26376
rect 21732 26324 21784 26376
rect 24492 26324 24544 26376
rect 21640 26256 21692 26308
rect 26700 26299 26752 26308
rect 26700 26265 26709 26299
rect 26709 26265 26743 26299
rect 26743 26265 26752 26299
rect 26700 26256 26752 26265
rect 21272 26231 21324 26240
rect 21272 26197 21281 26231
rect 21281 26197 21315 26231
rect 21315 26197 21324 26231
rect 21272 26188 21324 26197
rect 24676 26231 24728 26240
rect 24676 26197 24685 26231
rect 24685 26197 24719 26231
rect 24719 26197 24728 26231
rect 24676 26188 24728 26197
rect 7896 26086 7948 26138
rect 7960 26086 8012 26138
rect 8024 26086 8076 26138
rect 8088 26086 8140 26138
rect 8152 26086 8204 26138
rect 14842 26086 14894 26138
rect 14906 26086 14958 26138
rect 14970 26086 15022 26138
rect 15034 26086 15086 26138
rect 15098 26086 15150 26138
rect 21788 26086 21840 26138
rect 21852 26086 21904 26138
rect 21916 26086 21968 26138
rect 21980 26086 22032 26138
rect 22044 26086 22096 26138
rect 28734 26086 28786 26138
rect 28798 26086 28850 26138
rect 28862 26086 28914 26138
rect 28926 26086 28978 26138
rect 28990 26086 29042 26138
rect 19892 25984 19944 26036
rect 21364 25984 21416 26036
rect 23848 25984 23900 26036
rect 24584 25984 24636 26036
rect 1676 25891 1728 25900
rect 1676 25857 1685 25891
rect 1685 25857 1719 25891
rect 1719 25857 1728 25891
rect 1676 25848 1728 25857
rect 16764 25848 16816 25900
rect 17132 25891 17184 25900
rect 17132 25857 17166 25891
rect 17166 25857 17184 25891
rect 24768 25916 24820 25968
rect 17132 25848 17184 25857
rect 18880 25848 18932 25900
rect 20168 25848 20220 25900
rect 24676 25891 24728 25900
rect 24676 25857 24685 25891
rect 24685 25857 24719 25891
rect 24719 25857 24728 25891
rect 24676 25848 24728 25857
rect 26700 25984 26752 26036
rect 2412 25780 2464 25832
rect 2780 25823 2832 25832
rect 2780 25789 2789 25823
rect 2789 25789 2823 25823
rect 2823 25789 2832 25823
rect 2780 25780 2832 25789
rect 15568 25780 15620 25832
rect 15844 25823 15896 25832
rect 15844 25789 15853 25823
rect 15853 25789 15887 25823
rect 15887 25789 15896 25823
rect 15844 25780 15896 25789
rect 19984 25780 20036 25832
rect 20904 25780 20956 25832
rect 23388 25780 23440 25832
rect 25780 25848 25832 25900
rect 26608 25891 26660 25900
rect 26608 25857 26617 25891
rect 26617 25857 26651 25891
rect 26651 25857 26660 25891
rect 26608 25848 26660 25857
rect 26884 25848 26936 25900
rect 25044 25780 25096 25832
rect 26148 25780 26200 25832
rect 27344 25712 27396 25764
rect 16120 25644 16172 25696
rect 20168 25687 20220 25696
rect 20168 25653 20177 25687
rect 20177 25653 20211 25687
rect 20211 25653 20220 25687
rect 20168 25644 20220 25653
rect 20628 25687 20680 25696
rect 20628 25653 20637 25687
rect 20637 25653 20671 25687
rect 20671 25653 20680 25687
rect 20628 25644 20680 25653
rect 22560 25644 22612 25696
rect 24032 25644 24084 25696
rect 24676 25644 24728 25696
rect 25596 25644 25648 25696
rect 26056 25644 26108 25696
rect 28356 25644 28408 25696
rect 4423 25542 4475 25594
rect 4487 25542 4539 25594
rect 4551 25542 4603 25594
rect 4615 25542 4667 25594
rect 4679 25542 4731 25594
rect 11369 25542 11421 25594
rect 11433 25542 11485 25594
rect 11497 25542 11549 25594
rect 11561 25542 11613 25594
rect 11625 25542 11677 25594
rect 18315 25542 18367 25594
rect 18379 25542 18431 25594
rect 18443 25542 18495 25594
rect 18507 25542 18559 25594
rect 18571 25542 18623 25594
rect 25261 25542 25313 25594
rect 25325 25542 25377 25594
rect 25389 25542 25441 25594
rect 25453 25542 25505 25594
rect 25517 25542 25569 25594
rect 2412 25483 2464 25492
rect 2412 25449 2421 25483
rect 2421 25449 2455 25483
rect 2455 25449 2464 25483
rect 2412 25440 2464 25449
rect 17132 25483 17184 25492
rect 17132 25449 17141 25483
rect 17141 25449 17175 25483
rect 17175 25449 17184 25483
rect 17132 25440 17184 25449
rect 18880 25483 18932 25492
rect 18880 25449 18889 25483
rect 18889 25449 18923 25483
rect 18923 25449 18932 25483
rect 18880 25440 18932 25449
rect 20812 25483 20864 25492
rect 20812 25449 20821 25483
rect 20821 25449 20855 25483
rect 20855 25449 20864 25483
rect 20812 25440 20864 25449
rect 23388 25483 23440 25492
rect 23388 25449 23397 25483
rect 23397 25449 23431 25483
rect 23431 25449 23440 25483
rect 23388 25440 23440 25449
rect 24584 25440 24636 25492
rect 25780 25440 25832 25492
rect 1584 25279 1636 25288
rect 1584 25245 1593 25279
rect 1593 25245 1627 25279
rect 1627 25245 1636 25279
rect 1584 25236 1636 25245
rect 4252 25236 4304 25288
rect 16120 25279 16172 25288
rect 16120 25245 16129 25279
rect 16129 25245 16163 25279
rect 16163 25245 16172 25279
rect 16120 25236 16172 25245
rect 20628 25304 20680 25356
rect 21272 25347 21324 25356
rect 21272 25313 21281 25347
rect 21281 25313 21315 25347
rect 21315 25313 21324 25347
rect 21272 25304 21324 25313
rect 22468 25304 22520 25356
rect 24768 25347 24820 25356
rect 24768 25313 24777 25347
rect 24777 25313 24811 25347
rect 24811 25313 24820 25347
rect 24768 25304 24820 25313
rect 24952 25304 25004 25356
rect 19708 25279 19760 25288
rect 19708 25245 19717 25279
rect 19717 25245 19751 25279
rect 19751 25245 19760 25279
rect 20996 25279 21048 25288
rect 19708 25236 19760 25245
rect 20996 25245 21005 25279
rect 21005 25245 21039 25279
rect 21039 25245 21048 25279
rect 20996 25236 21048 25245
rect 22376 25236 22428 25288
rect 24492 25236 24544 25288
rect 17132 25168 17184 25220
rect 24860 25236 24912 25288
rect 25964 25304 26016 25356
rect 27528 25347 27580 25356
rect 27528 25313 27537 25347
rect 27537 25313 27571 25347
rect 27571 25313 27580 25347
rect 27528 25304 27580 25313
rect 28356 25347 28408 25356
rect 28356 25313 28365 25347
rect 28365 25313 28399 25347
rect 28399 25313 28408 25347
rect 28356 25304 28408 25313
rect 25228 25168 25280 25220
rect 28172 25211 28224 25220
rect 28172 25177 28181 25211
rect 28181 25177 28215 25211
rect 28215 25177 28224 25211
rect 28172 25168 28224 25177
rect 1768 25143 1820 25152
rect 1768 25109 1777 25143
rect 1777 25109 1811 25143
rect 1811 25109 1820 25143
rect 1768 25100 1820 25109
rect 23848 25100 23900 25152
rect 25044 25143 25096 25152
rect 25044 25109 25053 25143
rect 25053 25109 25087 25143
rect 25087 25109 25096 25143
rect 25044 25100 25096 25109
rect 7896 24998 7948 25050
rect 7960 24998 8012 25050
rect 8024 24998 8076 25050
rect 8088 24998 8140 25050
rect 8152 24998 8204 25050
rect 14842 24998 14894 25050
rect 14906 24998 14958 25050
rect 14970 24998 15022 25050
rect 15034 24998 15086 25050
rect 15098 24998 15150 25050
rect 21788 24998 21840 25050
rect 21852 24998 21904 25050
rect 21916 24998 21968 25050
rect 21980 24998 22032 25050
rect 22044 24998 22096 25050
rect 28734 24998 28786 25050
rect 28798 24998 28850 25050
rect 28862 24998 28914 25050
rect 28926 24998 28978 25050
rect 28990 24998 29042 25050
rect 1768 24896 1820 24948
rect 15844 24896 15896 24948
rect 22376 24939 22428 24948
rect 22376 24905 22385 24939
rect 22385 24905 22419 24939
rect 22419 24905 22428 24939
rect 22376 24896 22428 24905
rect 28172 24939 28224 24948
rect 28172 24905 28181 24939
rect 28181 24905 28215 24939
rect 28215 24905 28224 24939
rect 28172 24896 28224 24905
rect 17132 24828 17184 24880
rect 20904 24828 20956 24880
rect 22744 24871 22796 24880
rect 17224 24760 17276 24812
rect 21640 24760 21692 24812
rect 21824 24760 21876 24812
rect 22744 24837 22753 24871
rect 22753 24837 22787 24871
rect 22787 24837 22796 24871
rect 22744 24828 22796 24837
rect 23388 24828 23440 24880
rect 23756 24803 23808 24812
rect 23756 24769 23765 24803
rect 23765 24769 23799 24803
rect 23799 24769 23808 24803
rect 23756 24760 23808 24769
rect 24400 24803 24452 24812
rect 24400 24769 24409 24803
rect 24409 24769 24443 24803
rect 24443 24769 24452 24803
rect 24400 24760 24452 24769
rect 25228 24803 25280 24812
rect 25228 24769 25237 24803
rect 25237 24769 25271 24803
rect 25271 24769 25280 24803
rect 25228 24760 25280 24769
rect 16856 24599 16908 24608
rect 16856 24565 16865 24599
rect 16865 24565 16899 24599
rect 16899 24565 16908 24599
rect 16856 24556 16908 24565
rect 23572 24624 23624 24676
rect 23296 24556 23348 24608
rect 24584 24624 24636 24676
rect 25504 24803 25556 24812
rect 25504 24769 25513 24803
rect 25513 24769 25547 24803
rect 25547 24769 25556 24803
rect 25504 24760 25556 24769
rect 25780 24760 25832 24812
rect 25872 24803 25924 24812
rect 25872 24769 25881 24803
rect 25881 24769 25915 24803
rect 25915 24769 25924 24803
rect 25872 24760 25924 24769
rect 27436 24803 27488 24812
rect 27436 24769 27445 24803
rect 27445 24769 27479 24803
rect 27479 24769 27488 24803
rect 27436 24760 27488 24769
rect 28080 24803 28132 24812
rect 28080 24769 28089 24803
rect 28089 24769 28123 24803
rect 28123 24769 28132 24803
rect 28080 24760 28132 24769
rect 26424 24692 26476 24744
rect 26700 24692 26752 24744
rect 26240 24624 26292 24676
rect 26608 24624 26660 24676
rect 24676 24556 24728 24608
rect 25688 24556 25740 24608
rect 26516 24599 26568 24608
rect 26516 24565 26525 24599
rect 26525 24565 26559 24599
rect 26559 24565 26568 24599
rect 26516 24556 26568 24565
rect 4423 24454 4475 24506
rect 4487 24454 4539 24506
rect 4551 24454 4603 24506
rect 4615 24454 4667 24506
rect 4679 24454 4731 24506
rect 11369 24454 11421 24506
rect 11433 24454 11485 24506
rect 11497 24454 11549 24506
rect 11561 24454 11613 24506
rect 11625 24454 11677 24506
rect 18315 24454 18367 24506
rect 18379 24454 18431 24506
rect 18443 24454 18495 24506
rect 18507 24454 18559 24506
rect 18571 24454 18623 24506
rect 25261 24454 25313 24506
rect 25325 24454 25377 24506
rect 25389 24454 25441 24506
rect 25453 24454 25505 24506
rect 25517 24454 25569 24506
rect 15568 24216 15620 24268
rect 19432 24352 19484 24404
rect 22744 24352 22796 24404
rect 24400 24352 24452 24404
rect 26424 24352 26476 24404
rect 27436 24352 27488 24404
rect 27896 24216 27948 24268
rect 28356 24259 28408 24268
rect 28356 24225 28365 24259
rect 28365 24225 28399 24259
rect 28399 24225 28408 24259
rect 28356 24216 28408 24225
rect 16764 24191 16816 24200
rect 16764 24157 16773 24191
rect 16773 24157 16807 24191
rect 16807 24157 16816 24191
rect 16764 24148 16816 24157
rect 16856 24148 16908 24200
rect 18788 24191 18840 24200
rect 18788 24157 18797 24191
rect 18797 24157 18831 24191
rect 18831 24157 18840 24191
rect 18788 24148 18840 24157
rect 20076 24148 20128 24200
rect 21548 24148 21600 24200
rect 21732 24148 21784 24200
rect 21364 24080 21416 24132
rect 9404 24012 9456 24064
rect 16856 24012 16908 24064
rect 18604 24055 18656 24064
rect 18604 24021 18613 24055
rect 18613 24021 18647 24055
rect 18647 24021 18656 24055
rect 18604 24012 18656 24021
rect 21456 24055 21508 24064
rect 21456 24021 21465 24055
rect 21465 24021 21499 24055
rect 21499 24021 21508 24055
rect 21456 24012 21508 24021
rect 22836 24123 22888 24132
rect 22836 24089 22870 24123
rect 22870 24089 22888 24123
rect 22836 24080 22888 24089
rect 27344 24080 27396 24132
rect 21824 24012 21876 24064
rect 23756 24012 23808 24064
rect 24216 24012 24268 24064
rect 7896 23910 7948 23962
rect 7960 23910 8012 23962
rect 8024 23910 8076 23962
rect 8088 23910 8140 23962
rect 8152 23910 8204 23962
rect 14842 23910 14894 23962
rect 14906 23910 14958 23962
rect 14970 23910 15022 23962
rect 15034 23910 15086 23962
rect 15098 23910 15150 23962
rect 21788 23910 21840 23962
rect 21852 23910 21904 23962
rect 21916 23910 21968 23962
rect 21980 23910 22032 23962
rect 22044 23910 22096 23962
rect 28734 23910 28786 23962
rect 28798 23910 28850 23962
rect 28862 23910 28914 23962
rect 28926 23910 28978 23962
rect 28990 23910 29042 23962
rect 17224 23851 17276 23860
rect 17224 23817 17233 23851
rect 17233 23817 17267 23851
rect 17267 23817 17276 23851
rect 17224 23808 17276 23817
rect 20076 23851 20128 23860
rect 20076 23817 20085 23851
rect 20085 23817 20119 23851
rect 20119 23817 20128 23851
rect 20076 23808 20128 23817
rect 22836 23851 22888 23860
rect 22836 23817 22845 23851
rect 22845 23817 22879 23851
rect 22879 23817 22888 23851
rect 22836 23808 22888 23817
rect 24952 23851 25004 23860
rect 24952 23817 24961 23851
rect 24961 23817 24995 23851
rect 24995 23817 25004 23851
rect 24952 23808 25004 23817
rect 25780 23851 25832 23860
rect 25780 23817 25789 23851
rect 25789 23817 25823 23851
rect 25823 23817 25832 23851
rect 25780 23808 25832 23817
rect 26240 23851 26292 23860
rect 26240 23817 26249 23851
rect 26249 23817 26283 23851
rect 26283 23817 26292 23851
rect 26240 23808 26292 23817
rect 16856 23783 16908 23792
rect 16856 23749 16865 23783
rect 16865 23749 16899 23783
rect 16899 23749 16908 23783
rect 16856 23740 16908 23749
rect 17132 23740 17184 23792
rect 18604 23740 18656 23792
rect 21364 23740 21416 23792
rect 22376 23783 22428 23792
rect 22376 23749 22385 23783
rect 22385 23749 22419 23783
rect 22419 23749 22428 23783
rect 22376 23740 22428 23749
rect 22744 23740 22796 23792
rect 21180 23715 21232 23724
rect 24216 23740 24268 23792
rect 21180 23681 21198 23715
rect 21198 23681 21232 23715
rect 21180 23672 21232 23681
rect 16764 23604 16816 23656
rect 21640 23604 21692 23656
rect 23296 23715 23348 23724
rect 23296 23681 23305 23715
rect 23305 23681 23339 23715
rect 23339 23681 23348 23715
rect 23296 23672 23348 23681
rect 25136 23740 25188 23792
rect 24768 23715 24820 23724
rect 24768 23681 24777 23715
rect 24777 23681 24811 23715
rect 24811 23681 24820 23715
rect 24768 23672 24820 23681
rect 26424 23715 26476 23724
rect 23940 23604 23992 23656
rect 24308 23604 24360 23656
rect 26424 23681 26433 23715
rect 26433 23681 26467 23715
rect 26467 23681 26476 23715
rect 26424 23672 26476 23681
rect 26516 23672 26568 23724
rect 26792 23672 26844 23724
rect 27068 23672 27120 23724
rect 23664 23536 23716 23588
rect 26700 23604 26752 23656
rect 19616 23511 19668 23520
rect 19616 23477 19625 23511
rect 19625 23477 19659 23511
rect 19659 23477 19668 23511
rect 19616 23468 19668 23477
rect 22008 23511 22060 23520
rect 22008 23477 22017 23511
rect 22017 23477 22051 23511
rect 22051 23477 22060 23511
rect 22008 23468 22060 23477
rect 24400 23468 24452 23520
rect 26700 23468 26752 23520
rect 27436 23468 27488 23520
rect 4423 23366 4475 23418
rect 4487 23366 4539 23418
rect 4551 23366 4603 23418
rect 4615 23366 4667 23418
rect 4679 23366 4731 23418
rect 11369 23366 11421 23418
rect 11433 23366 11485 23418
rect 11497 23366 11549 23418
rect 11561 23366 11613 23418
rect 11625 23366 11677 23418
rect 18315 23366 18367 23418
rect 18379 23366 18431 23418
rect 18443 23366 18495 23418
rect 18507 23366 18559 23418
rect 18571 23366 18623 23418
rect 25261 23366 25313 23418
rect 25325 23366 25377 23418
rect 25389 23366 25441 23418
rect 25453 23366 25505 23418
rect 25517 23366 25569 23418
rect 18788 23307 18840 23316
rect 18788 23273 18797 23307
rect 18797 23273 18831 23307
rect 18831 23273 18840 23307
rect 18788 23264 18840 23273
rect 21180 23264 21232 23316
rect 22008 23264 22060 23316
rect 16396 23103 16448 23112
rect 16396 23069 16405 23103
rect 16405 23069 16439 23103
rect 16439 23069 16448 23103
rect 16396 23060 16448 23069
rect 25228 23196 25280 23248
rect 19984 23171 20036 23180
rect 19984 23137 19993 23171
rect 19993 23137 20027 23171
rect 20027 23137 20036 23171
rect 19984 23128 20036 23137
rect 21456 23171 21508 23180
rect 21456 23137 21465 23171
rect 21465 23137 21499 23171
rect 21499 23137 21508 23171
rect 21456 23128 21508 23137
rect 25044 23128 25096 23180
rect 19616 23060 19668 23112
rect 20076 23060 20128 23112
rect 20996 23060 21048 23112
rect 25136 23060 25188 23112
rect 26148 23196 26200 23248
rect 27436 23196 27488 23248
rect 26700 23171 26752 23180
rect 26700 23137 26709 23171
rect 26709 23137 26743 23171
rect 26743 23137 26752 23171
rect 26700 23128 26752 23137
rect 29920 23128 29972 23180
rect 18788 22992 18840 23044
rect 19708 22992 19760 23044
rect 24308 22992 24360 23044
rect 16580 22967 16632 22976
rect 16580 22933 16589 22967
rect 16589 22933 16623 22967
rect 16623 22933 16632 22967
rect 16580 22924 16632 22933
rect 25872 22967 25924 22976
rect 25872 22933 25881 22967
rect 25881 22933 25915 22967
rect 25915 22933 25924 22967
rect 25872 22924 25924 22933
rect 7896 22822 7948 22874
rect 7960 22822 8012 22874
rect 8024 22822 8076 22874
rect 8088 22822 8140 22874
rect 8152 22822 8204 22874
rect 14842 22822 14894 22874
rect 14906 22822 14958 22874
rect 14970 22822 15022 22874
rect 15034 22822 15086 22874
rect 15098 22822 15150 22874
rect 21788 22822 21840 22874
rect 21852 22822 21904 22874
rect 21916 22822 21968 22874
rect 21980 22822 22032 22874
rect 22044 22822 22096 22874
rect 28734 22822 28786 22874
rect 28798 22822 28850 22874
rect 28862 22822 28914 22874
rect 28926 22822 28978 22874
rect 28990 22822 29042 22874
rect 18144 22720 18196 22772
rect 20536 22720 20588 22772
rect 24032 22720 24084 22772
rect 24768 22720 24820 22772
rect 26424 22720 26476 22772
rect 27344 22763 27396 22772
rect 27344 22729 27353 22763
rect 27353 22729 27387 22763
rect 27387 22729 27396 22763
rect 27344 22720 27396 22729
rect 16580 22652 16632 22704
rect 22376 22695 22428 22704
rect 22376 22661 22385 22695
rect 22385 22661 22419 22695
rect 22419 22661 22428 22695
rect 22376 22652 22428 22661
rect 24216 22695 24268 22704
rect 24216 22661 24225 22695
rect 24225 22661 24259 22695
rect 24259 22661 24268 22695
rect 24216 22652 24268 22661
rect 1860 22516 1912 22568
rect 23664 22584 23716 22636
rect 25872 22652 25924 22704
rect 27252 22584 27304 22636
rect 27896 22627 27948 22636
rect 27896 22593 27905 22627
rect 27905 22593 27939 22627
rect 27939 22593 27948 22627
rect 27896 22584 27948 22593
rect 15384 22516 15436 22568
rect 16672 22516 16724 22568
rect 16764 22516 16816 22568
rect 25044 22516 25096 22568
rect 23940 22448 23992 22500
rect 16120 22423 16172 22432
rect 16120 22389 16129 22423
rect 16129 22389 16163 22423
rect 16163 22389 16172 22423
rect 16120 22380 16172 22389
rect 21272 22380 21324 22432
rect 24308 22380 24360 22432
rect 24400 22423 24452 22432
rect 24400 22389 24409 22423
rect 24409 22389 24443 22423
rect 24443 22389 24452 22423
rect 24400 22380 24452 22389
rect 4423 22278 4475 22330
rect 4487 22278 4539 22330
rect 4551 22278 4603 22330
rect 4615 22278 4667 22330
rect 4679 22278 4731 22330
rect 11369 22278 11421 22330
rect 11433 22278 11485 22330
rect 11497 22278 11549 22330
rect 11561 22278 11613 22330
rect 11625 22278 11677 22330
rect 18315 22278 18367 22330
rect 18379 22278 18431 22330
rect 18443 22278 18495 22330
rect 18507 22278 18559 22330
rect 18571 22278 18623 22330
rect 25261 22278 25313 22330
rect 25325 22278 25377 22330
rect 25389 22278 25441 22330
rect 25453 22278 25505 22330
rect 25517 22278 25569 22330
rect 16396 22176 16448 22228
rect 22376 22176 22428 22228
rect 24860 22083 24912 22092
rect 24860 22049 24869 22083
rect 24869 22049 24903 22083
rect 24903 22049 24912 22083
rect 24860 22040 24912 22049
rect 16120 22015 16172 22024
rect 16120 21981 16129 22015
rect 16129 21981 16163 22015
rect 16163 21981 16172 22015
rect 16120 21972 16172 21981
rect 16580 22015 16632 22024
rect 16580 21981 16589 22015
rect 16589 21981 16623 22015
rect 16623 21981 16632 22015
rect 16580 21972 16632 21981
rect 19708 21972 19760 22024
rect 21456 21972 21508 22024
rect 23664 22015 23716 22024
rect 23664 21981 23673 22015
rect 23673 21981 23707 22015
rect 23707 21981 23716 22015
rect 23664 21972 23716 21981
rect 24584 22015 24636 22024
rect 24584 21981 24593 22015
rect 24593 21981 24627 22015
rect 24627 21981 24636 22015
rect 24584 21972 24636 21981
rect 16212 21904 16264 21956
rect 23940 21947 23992 21956
rect 16948 21836 17000 21888
rect 21180 21879 21232 21888
rect 21180 21845 21189 21879
rect 21189 21845 21223 21879
rect 21223 21845 21232 21879
rect 21180 21836 21232 21845
rect 21364 21836 21416 21888
rect 22284 21836 22336 21888
rect 22744 21879 22796 21888
rect 22744 21845 22753 21879
rect 22753 21845 22787 21879
rect 22787 21845 22796 21879
rect 22744 21836 22796 21845
rect 23940 21913 23949 21947
rect 23949 21913 23983 21947
rect 23983 21913 23992 21947
rect 23940 21904 23992 21913
rect 24492 21904 24544 21956
rect 25964 22040 26016 22092
rect 27528 22083 27580 22092
rect 27528 22049 27537 22083
rect 27537 22049 27571 22083
rect 27571 22049 27580 22083
rect 27528 22040 27580 22049
rect 28356 22015 28408 22024
rect 28356 21981 28365 22015
rect 28365 21981 28399 22015
rect 28399 21981 28408 22015
rect 28356 21972 28408 21981
rect 28172 21947 28224 21956
rect 28172 21913 28181 21947
rect 28181 21913 28215 21947
rect 28215 21913 28224 21947
rect 28172 21904 28224 21913
rect 23756 21879 23808 21888
rect 23756 21845 23765 21879
rect 23765 21845 23799 21879
rect 23799 21845 23808 21879
rect 23756 21836 23808 21845
rect 24216 21836 24268 21888
rect 24768 21836 24820 21888
rect 25136 21836 25188 21888
rect 7896 21734 7948 21786
rect 7960 21734 8012 21786
rect 8024 21734 8076 21786
rect 8088 21734 8140 21786
rect 8152 21734 8204 21786
rect 14842 21734 14894 21786
rect 14906 21734 14958 21786
rect 14970 21734 15022 21786
rect 15034 21734 15086 21786
rect 15098 21734 15150 21786
rect 21788 21734 21840 21786
rect 21852 21734 21904 21786
rect 21916 21734 21968 21786
rect 21980 21734 22032 21786
rect 22044 21734 22096 21786
rect 28734 21734 28786 21786
rect 28798 21734 28850 21786
rect 28862 21734 28914 21786
rect 28926 21734 28978 21786
rect 28990 21734 29042 21786
rect 19064 21632 19116 21684
rect 28172 21675 28224 21684
rect 28172 21641 28181 21675
rect 28181 21641 28215 21675
rect 28215 21641 28224 21675
rect 28172 21632 28224 21641
rect 15200 21496 15252 21548
rect 16764 21496 16816 21548
rect 16948 21496 17000 21548
rect 21088 21564 21140 21616
rect 18972 21539 19024 21548
rect 18972 21505 19006 21539
rect 19006 21505 19024 21539
rect 20996 21539 21048 21548
rect 18972 21496 19024 21505
rect 20996 21505 21005 21539
rect 21005 21505 21039 21539
rect 21039 21505 21048 21539
rect 20996 21496 21048 21505
rect 21180 21496 21232 21548
rect 22744 21539 22796 21548
rect 15660 21428 15712 21480
rect 16856 21360 16908 21412
rect 21272 21360 21324 21412
rect 22744 21505 22753 21539
rect 22753 21505 22787 21539
rect 22787 21505 22796 21539
rect 22744 21496 22796 21505
rect 25136 21539 25188 21548
rect 25136 21505 25145 21539
rect 25145 21505 25179 21539
rect 25179 21505 25188 21539
rect 25136 21496 25188 21505
rect 25228 21496 25280 21548
rect 25688 21496 25740 21548
rect 28356 21564 28408 21616
rect 22836 21471 22888 21480
rect 22836 21437 22845 21471
rect 22845 21437 22879 21471
rect 22879 21437 22888 21471
rect 22836 21428 22888 21437
rect 28264 21496 28316 21548
rect 24952 21360 25004 21412
rect 27620 21360 27672 21412
rect 16304 21335 16356 21344
rect 16304 21301 16313 21335
rect 16313 21301 16347 21335
rect 16347 21301 16356 21335
rect 16304 21292 16356 21301
rect 20076 21335 20128 21344
rect 20076 21301 20085 21335
rect 20085 21301 20119 21335
rect 20119 21301 20128 21335
rect 20076 21292 20128 21301
rect 20812 21335 20864 21344
rect 20812 21301 20821 21335
rect 20821 21301 20855 21335
rect 20855 21301 20864 21335
rect 20812 21292 20864 21301
rect 22376 21335 22428 21344
rect 22376 21301 22385 21335
rect 22385 21301 22419 21335
rect 22419 21301 22428 21335
rect 22376 21292 22428 21301
rect 25596 21292 25648 21344
rect 4423 21190 4475 21242
rect 4487 21190 4539 21242
rect 4551 21190 4603 21242
rect 4615 21190 4667 21242
rect 4679 21190 4731 21242
rect 11369 21190 11421 21242
rect 11433 21190 11485 21242
rect 11497 21190 11549 21242
rect 11561 21190 11613 21242
rect 11625 21190 11677 21242
rect 18315 21190 18367 21242
rect 18379 21190 18431 21242
rect 18443 21190 18495 21242
rect 18507 21190 18559 21242
rect 18571 21190 18623 21242
rect 25261 21190 25313 21242
rect 25325 21190 25377 21242
rect 25389 21190 25441 21242
rect 25453 21190 25505 21242
rect 25517 21190 25569 21242
rect 14740 21088 14792 21140
rect 16580 21088 16632 21140
rect 19708 21131 19760 21140
rect 19708 21097 19717 21131
rect 19717 21097 19751 21131
rect 19751 21097 19760 21131
rect 19708 21088 19760 21097
rect 18788 20952 18840 21004
rect 21088 20995 21140 21004
rect 21088 20961 21097 20995
rect 21097 20961 21131 20995
rect 21131 20961 21140 20995
rect 21088 20952 21140 20961
rect 21640 20952 21692 21004
rect 27528 20995 27580 21004
rect 27528 20961 27537 20995
rect 27537 20961 27571 20995
rect 27571 20961 27580 20995
rect 27528 20952 27580 20961
rect 16304 20927 16356 20936
rect 16304 20893 16313 20927
rect 16313 20893 16347 20927
rect 16347 20893 16356 20927
rect 16304 20884 16356 20893
rect 19524 20884 19576 20936
rect 20812 20927 20864 20936
rect 20812 20893 20830 20927
rect 20830 20893 20864 20927
rect 20812 20884 20864 20893
rect 22376 20884 22428 20936
rect 24952 20884 25004 20936
rect 25596 20927 25648 20936
rect 25596 20893 25605 20927
rect 25605 20893 25639 20927
rect 25639 20893 25648 20927
rect 25596 20884 25648 20893
rect 25688 20927 25740 20936
rect 25688 20893 25697 20927
rect 25697 20893 25731 20927
rect 25731 20893 25740 20927
rect 25688 20884 25740 20893
rect 25964 20884 26016 20936
rect 28356 20927 28408 20936
rect 28356 20893 28365 20927
rect 28365 20893 28399 20927
rect 28399 20893 28408 20927
rect 28356 20884 28408 20893
rect 14740 20816 14792 20868
rect 15384 20859 15436 20868
rect 15384 20825 15393 20859
rect 15393 20825 15427 20859
rect 15427 20825 15436 20859
rect 15384 20816 15436 20825
rect 16212 20816 16264 20868
rect 28172 20859 28224 20868
rect 28172 20825 28181 20859
rect 28181 20825 28215 20859
rect 28215 20825 28224 20859
rect 28172 20816 28224 20825
rect 18696 20748 18748 20800
rect 22468 20748 22520 20800
rect 26056 20791 26108 20800
rect 26056 20757 26065 20791
rect 26065 20757 26099 20791
rect 26099 20757 26108 20791
rect 26056 20748 26108 20757
rect 7896 20646 7948 20698
rect 7960 20646 8012 20698
rect 8024 20646 8076 20698
rect 8088 20646 8140 20698
rect 8152 20646 8204 20698
rect 14842 20646 14894 20698
rect 14906 20646 14958 20698
rect 14970 20646 15022 20698
rect 15034 20646 15086 20698
rect 15098 20646 15150 20698
rect 21788 20646 21840 20698
rect 21852 20646 21904 20698
rect 21916 20646 21968 20698
rect 21980 20646 22032 20698
rect 22044 20646 22096 20698
rect 28734 20646 28786 20698
rect 28798 20646 28850 20698
rect 28862 20646 28914 20698
rect 28926 20646 28978 20698
rect 28990 20646 29042 20698
rect 12624 20587 12676 20596
rect 12624 20553 12633 20587
rect 12633 20553 12667 20587
rect 12667 20553 12676 20587
rect 12624 20544 12676 20553
rect 18972 20544 19024 20596
rect 19524 20587 19576 20596
rect 19524 20553 19533 20587
rect 19533 20553 19567 20587
rect 19567 20553 19576 20587
rect 19524 20544 19576 20553
rect 19800 20544 19852 20596
rect 20076 20544 20128 20596
rect 22836 20544 22888 20596
rect 24676 20544 24728 20596
rect 28172 20587 28224 20596
rect 14464 20476 14516 20528
rect 19708 20476 19760 20528
rect 23664 20476 23716 20528
rect 24952 20476 25004 20528
rect 2504 20451 2556 20460
rect 2504 20417 2513 20451
rect 2513 20417 2547 20451
rect 2547 20417 2556 20451
rect 2504 20408 2556 20417
rect 12992 20451 13044 20460
rect 12992 20417 13001 20451
rect 13001 20417 13035 20451
rect 13035 20417 13044 20451
rect 12992 20408 13044 20417
rect 13084 20451 13136 20460
rect 13084 20417 13093 20451
rect 13093 20417 13127 20451
rect 13127 20417 13136 20451
rect 14648 20451 14700 20460
rect 13084 20408 13136 20417
rect 14648 20417 14657 20451
rect 14657 20417 14691 20451
rect 14691 20417 14700 20451
rect 14648 20408 14700 20417
rect 14832 20408 14884 20460
rect 18696 20451 18748 20460
rect 18696 20417 18705 20451
rect 18705 20417 18739 20451
rect 18739 20417 18748 20451
rect 18696 20408 18748 20417
rect 21456 20408 21508 20460
rect 22376 20451 22428 20460
rect 22376 20417 22385 20451
rect 22385 20417 22419 20451
rect 22419 20417 22428 20451
rect 22376 20408 22428 20417
rect 13820 20340 13872 20392
rect 19984 20340 20036 20392
rect 22468 20340 22520 20392
rect 23940 20408 23992 20460
rect 24584 20340 24636 20392
rect 25136 20408 25188 20460
rect 25688 20476 25740 20528
rect 28172 20553 28181 20587
rect 28181 20553 28215 20587
rect 28215 20553 28224 20587
rect 28172 20544 28224 20553
rect 28080 20451 28132 20460
rect 28080 20417 28089 20451
rect 28089 20417 28123 20451
rect 28123 20417 28132 20451
rect 28080 20408 28132 20417
rect 25964 20340 26016 20392
rect 28356 20340 28408 20392
rect 26332 20272 26384 20324
rect 1584 20204 1636 20256
rect 1768 20204 1820 20256
rect 25688 20247 25740 20256
rect 25688 20213 25697 20247
rect 25697 20213 25731 20247
rect 25731 20213 25740 20247
rect 25688 20204 25740 20213
rect 4423 20102 4475 20154
rect 4487 20102 4539 20154
rect 4551 20102 4603 20154
rect 4615 20102 4667 20154
rect 4679 20102 4731 20154
rect 11369 20102 11421 20154
rect 11433 20102 11485 20154
rect 11497 20102 11549 20154
rect 11561 20102 11613 20154
rect 11625 20102 11677 20154
rect 18315 20102 18367 20154
rect 18379 20102 18431 20154
rect 18443 20102 18495 20154
rect 18507 20102 18559 20154
rect 18571 20102 18623 20154
rect 25261 20102 25313 20154
rect 25325 20102 25377 20154
rect 25389 20102 25441 20154
rect 25453 20102 25505 20154
rect 25517 20102 25569 20154
rect 13084 20000 13136 20052
rect 14648 20043 14700 20052
rect 14648 20009 14657 20043
rect 14657 20009 14691 20043
rect 14691 20009 14700 20043
rect 14648 20000 14700 20009
rect 14740 20000 14792 20052
rect 15384 20000 15436 20052
rect 25136 20043 25188 20052
rect 25136 20009 25145 20043
rect 25145 20009 25179 20043
rect 25179 20009 25188 20043
rect 25136 20000 25188 20009
rect 25964 20000 26016 20052
rect 1584 19907 1636 19916
rect 1584 19873 1593 19907
rect 1593 19873 1627 19907
rect 1627 19873 1636 19907
rect 1584 19864 1636 19873
rect 1768 19907 1820 19916
rect 1768 19873 1777 19907
rect 1777 19873 1811 19907
rect 1811 19873 1820 19907
rect 1768 19864 1820 19873
rect 2780 19907 2832 19916
rect 2780 19873 2789 19907
rect 2789 19873 2823 19907
rect 2823 19873 2832 19907
rect 2780 19864 2832 19873
rect 23940 19864 23992 19916
rect 24492 19864 24544 19916
rect 24768 19864 24820 19916
rect 13728 19796 13780 19848
rect 14556 19796 14608 19848
rect 14648 19796 14700 19848
rect 16580 19796 16632 19848
rect 24860 19839 24912 19848
rect 14004 19728 14056 19780
rect 15936 19728 15988 19780
rect 24860 19805 24869 19839
rect 24869 19805 24903 19839
rect 24903 19805 24912 19839
rect 24860 19796 24912 19805
rect 25044 19864 25096 19916
rect 25596 19796 25648 19848
rect 26056 19839 26108 19848
rect 26056 19805 26090 19839
rect 26090 19805 26108 19839
rect 26056 19796 26108 19805
rect 27896 19839 27948 19848
rect 27896 19805 27905 19839
rect 27905 19805 27939 19839
rect 27939 19805 27948 19839
rect 27896 19796 27948 19805
rect 24676 19728 24728 19780
rect 14280 19660 14332 19712
rect 14740 19660 14792 19712
rect 17224 19660 17276 19712
rect 7896 19558 7948 19610
rect 7960 19558 8012 19610
rect 8024 19558 8076 19610
rect 8088 19558 8140 19610
rect 8152 19558 8204 19610
rect 14842 19558 14894 19610
rect 14906 19558 14958 19610
rect 14970 19558 15022 19610
rect 15034 19558 15086 19610
rect 15098 19558 15150 19610
rect 21788 19558 21840 19610
rect 21852 19558 21904 19610
rect 21916 19558 21968 19610
rect 21980 19558 22032 19610
rect 22044 19558 22096 19610
rect 28734 19558 28786 19610
rect 28798 19558 28850 19610
rect 28862 19558 28914 19610
rect 28926 19558 28978 19610
rect 28990 19558 29042 19610
rect 13820 19456 13872 19508
rect 14096 19456 14148 19508
rect 14464 19499 14516 19508
rect 14464 19465 14473 19499
rect 14473 19465 14507 19499
rect 14507 19465 14516 19499
rect 14464 19456 14516 19465
rect 14740 19456 14792 19508
rect 16948 19456 17000 19508
rect 12808 19388 12860 19440
rect 13728 19363 13780 19372
rect 13728 19329 13737 19363
rect 13737 19329 13771 19363
rect 13771 19329 13780 19363
rect 13728 19320 13780 19329
rect 14004 19320 14056 19372
rect 14556 19388 14608 19440
rect 19616 19499 19668 19508
rect 19616 19465 19625 19499
rect 19625 19465 19659 19499
rect 19659 19465 19668 19499
rect 19616 19456 19668 19465
rect 17224 19431 17276 19440
rect 17224 19397 17258 19431
rect 17258 19397 17276 19431
rect 17224 19388 17276 19397
rect 15936 19320 15988 19372
rect 16304 19320 16356 19372
rect 16764 19320 16816 19372
rect 19340 19320 19392 19372
rect 21180 19363 21232 19372
rect 21180 19329 21189 19363
rect 21189 19329 21223 19363
rect 21223 19329 21232 19363
rect 21180 19320 21232 19329
rect 1676 19295 1728 19304
rect 1676 19261 1685 19295
rect 1685 19261 1719 19295
rect 1719 19261 1728 19295
rect 1676 19252 1728 19261
rect 1860 19295 1912 19304
rect 1860 19261 1869 19295
rect 1869 19261 1903 19295
rect 1903 19261 1912 19295
rect 1860 19252 1912 19261
rect 2136 19295 2188 19304
rect 2136 19261 2145 19295
rect 2145 19261 2179 19295
rect 2179 19261 2188 19295
rect 2136 19252 2188 19261
rect 14280 19252 14332 19304
rect 14004 19184 14056 19236
rect 14740 19184 14792 19236
rect 20260 19252 20312 19304
rect 14556 19116 14608 19168
rect 17132 19116 17184 19168
rect 21088 19116 21140 19168
rect 28356 19116 28408 19168
rect 4423 19014 4475 19066
rect 4487 19014 4539 19066
rect 4551 19014 4603 19066
rect 4615 19014 4667 19066
rect 4679 19014 4731 19066
rect 11369 19014 11421 19066
rect 11433 19014 11485 19066
rect 11497 19014 11549 19066
rect 11561 19014 11613 19066
rect 11625 19014 11677 19066
rect 18315 19014 18367 19066
rect 18379 19014 18431 19066
rect 18443 19014 18495 19066
rect 18507 19014 18559 19066
rect 18571 19014 18623 19066
rect 25261 19014 25313 19066
rect 25325 19014 25377 19066
rect 25389 19014 25441 19066
rect 25453 19014 25505 19066
rect 25517 19014 25569 19066
rect 1676 18912 1728 18964
rect 1860 18912 1912 18964
rect 12992 18912 13044 18964
rect 13820 18912 13872 18964
rect 16580 18912 16632 18964
rect 17040 18912 17092 18964
rect 24860 18912 24912 18964
rect 24216 18844 24268 18896
rect 2596 18751 2648 18760
rect 2596 18717 2605 18751
rect 2605 18717 2639 18751
rect 2639 18717 2648 18751
rect 2596 18708 2648 18717
rect 12256 18708 12308 18760
rect 14556 18776 14608 18828
rect 18052 18776 18104 18828
rect 24676 18819 24728 18828
rect 24676 18785 24685 18819
rect 24685 18785 24719 18819
rect 24719 18785 24728 18819
rect 24676 18776 24728 18785
rect 26148 18776 26200 18828
rect 28356 18819 28408 18828
rect 28356 18785 28365 18819
rect 28365 18785 28399 18819
rect 28399 18785 28408 18819
rect 28356 18776 28408 18785
rect 12808 18708 12860 18760
rect 13728 18708 13780 18760
rect 15660 18751 15712 18760
rect 15660 18717 15669 18751
rect 15669 18717 15703 18751
rect 15703 18717 15712 18751
rect 15660 18708 15712 18717
rect 16764 18708 16816 18760
rect 16948 18751 17000 18760
rect 16948 18717 16982 18751
rect 16982 18717 17000 18751
rect 16948 18708 17000 18717
rect 18696 18751 18748 18760
rect 18696 18717 18705 18751
rect 18705 18717 18739 18751
rect 18739 18717 18748 18751
rect 18696 18708 18748 18717
rect 19800 18751 19852 18760
rect 19800 18717 19809 18751
rect 19809 18717 19843 18751
rect 19843 18717 19852 18751
rect 19800 18708 19852 18717
rect 21088 18751 21140 18760
rect 21088 18717 21122 18751
rect 21122 18717 21140 18751
rect 21088 18708 21140 18717
rect 22376 18708 22428 18760
rect 23388 18708 23440 18760
rect 23756 18708 23808 18760
rect 24860 18708 24912 18760
rect 14004 18640 14056 18692
rect 14280 18683 14332 18692
rect 14280 18649 14289 18683
rect 14289 18649 14323 18683
rect 14323 18649 14332 18683
rect 14280 18640 14332 18649
rect 14740 18640 14792 18692
rect 15936 18640 15988 18692
rect 20260 18640 20312 18692
rect 20904 18640 20956 18692
rect 23112 18640 23164 18692
rect 23296 18640 23348 18692
rect 27988 18640 28040 18692
rect 13452 18615 13504 18624
rect 13452 18581 13461 18615
rect 13461 18581 13495 18615
rect 13495 18581 13504 18615
rect 13452 18572 13504 18581
rect 14648 18615 14700 18624
rect 14648 18581 14657 18615
rect 14657 18581 14691 18615
rect 14691 18581 14700 18615
rect 14648 18572 14700 18581
rect 17224 18572 17276 18624
rect 17960 18572 18012 18624
rect 18236 18572 18288 18624
rect 20812 18572 20864 18624
rect 22192 18615 22244 18624
rect 22192 18581 22201 18615
rect 22201 18581 22235 18615
rect 22235 18581 22244 18615
rect 22192 18572 22244 18581
rect 23020 18615 23072 18624
rect 23020 18581 23029 18615
rect 23029 18581 23063 18615
rect 23063 18581 23072 18615
rect 23020 18572 23072 18581
rect 23572 18572 23624 18624
rect 26700 18572 26752 18624
rect 7896 18470 7948 18522
rect 7960 18470 8012 18522
rect 8024 18470 8076 18522
rect 8088 18470 8140 18522
rect 8152 18470 8204 18522
rect 14842 18470 14894 18522
rect 14906 18470 14958 18522
rect 14970 18470 15022 18522
rect 15034 18470 15086 18522
rect 15098 18470 15150 18522
rect 21788 18470 21840 18522
rect 21852 18470 21904 18522
rect 21916 18470 21968 18522
rect 21980 18470 22032 18522
rect 22044 18470 22096 18522
rect 28734 18470 28786 18522
rect 28798 18470 28850 18522
rect 28862 18470 28914 18522
rect 28926 18470 28978 18522
rect 28990 18470 29042 18522
rect 16304 18411 16356 18420
rect 16304 18377 16313 18411
rect 16313 18377 16347 18411
rect 16347 18377 16356 18411
rect 16304 18368 16356 18377
rect 17224 18411 17276 18420
rect 17224 18377 17233 18411
rect 17233 18377 17267 18411
rect 17267 18377 17276 18411
rect 17224 18368 17276 18377
rect 21180 18368 21232 18420
rect 22192 18368 22244 18420
rect 22468 18411 22520 18420
rect 22468 18377 22477 18411
rect 22477 18377 22511 18411
rect 22511 18377 22520 18411
rect 22468 18368 22520 18377
rect 23020 18368 23072 18420
rect 24676 18368 24728 18420
rect 27988 18411 28040 18420
rect 27988 18377 27997 18411
rect 27997 18377 28031 18411
rect 28031 18377 28040 18411
rect 27988 18368 28040 18377
rect 14464 18300 14516 18352
rect 16120 18343 16172 18352
rect 1584 18275 1636 18284
rect 1584 18241 1593 18275
rect 1593 18241 1627 18275
rect 1627 18241 1636 18275
rect 1584 18232 1636 18241
rect 12256 18275 12308 18284
rect 12256 18241 12265 18275
rect 12265 18241 12299 18275
rect 12299 18241 12308 18275
rect 12256 18232 12308 18241
rect 11888 18164 11940 18216
rect 12900 18275 12952 18284
rect 12900 18241 12909 18275
rect 12909 18241 12943 18275
rect 12943 18241 12952 18275
rect 12900 18232 12952 18241
rect 13452 18232 13504 18284
rect 13820 18275 13872 18284
rect 13820 18241 13829 18275
rect 13829 18241 13863 18275
rect 13863 18241 13872 18275
rect 13820 18232 13872 18241
rect 14004 18275 14056 18284
rect 14004 18241 14012 18275
rect 14012 18241 14046 18275
rect 14046 18241 14056 18275
rect 14004 18232 14056 18241
rect 14096 18275 14148 18284
rect 14096 18241 14105 18275
rect 14105 18241 14139 18275
rect 14139 18241 14148 18275
rect 14556 18275 14608 18284
rect 14096 18232 14148 18241
rect 14556 18241 14565 18275
rect 14565 18241 14599 18275
rect 14599 18241 14608 18275
rect 14556 18232 14608 18241
rect 14740 18275 14792 18284
rect 14740 18241 14749 18275
rect 14749 18241 14783 18275
rect 14783 18241 14792 18275
rect 14740 18232 14792 18241
rect 16120 18309 16129 18343
rect 16129 18309 16163 18343
rect 16163 18309 16172 18343
rect 16120 18300 16172 18309
rect 16764 18300 16816 18352
rect 18052 18300 18104 18352
rect 22560 18300 22612 18352
rect 23112 18300 23164 18352
rect 25688 18300 25740 18352
rect 15752 18275 15804 18284
rect 15752 18241 15761 18275
rect 15761 18241 15795 18275
rect 15795 18241 15804 18275
rect 15752 18232 15804 18241
rect 17040 18275 17092 18284
rect 17040 18241 17049 18275
rect 17049 18241 17083 18275
rect 17083 18241 17092 18275
rect 17040 18232 17092 18241
rect 20904 18207 20956 18216
rect 20904 18173 20913 18207
rect 20913 18173 20947 18207
rect 20947 18173 20956 18207
rect 20904 18164 20956 18173
rect 15200 18096 15252 18148
rect 13452 18071 13504 18080
rect 13452 18037 13461 18071
rect 13461 18037 13495 18071
rect 13495 18037 13504 18071
rect 13452 18028 13504 18037
rect 14556 18071 14608 18080
rect 14556 18037 14565 18071
rect 14565 18037 14599 18071
rect 14599 18037 14608 18071
rect 14556 18028 14608 18037
rect 16856 18028 16908 18080
rect 17408 18028 17460 18080
rect 19984 18028 20036 18080
rect 23296 18164 23348 18216
rect 24216 18275 24268 18284
rect 24216 18241 24225 18275
rect 24225 18241 24259 18275
rect 24259 18241 24268 18275
rect 24216 18232 24268 18241
rect 25044 18232 25096 18284
rect 24584 18164 24636 18216
rect 23940 18096 23992 18148
rect 27620 18232 27672 18284
rect 23204 18071 23256 18080
rect 23204 18037 23213 18071
rect 23213 18037 23247 18071
rect 23247 18037 23256 18071
rect 23204 18028 23256 18037
rect 24400 18028 24452 18080
rect 4423 17926 4475 17978
rect 4487 17926 4539 17978
rect 4551 17926 4603 17978
rect 4615 17926 4667 17978
rect 4679 17926 4731 17978
rect 11369 17926 11421 17978
rect 11433 17926 11485 17978
rect 11497 17926 11549 17978
rect 11561 17926 11613 17978
rect 11625 17926 11677 17978
rect 18315 17926 18367 17978
rect 18379 17926 18431 17978
rect 18443 17926 18495 17978
rect 18507 17926 18559 17978
rect 18571 17926 18623 17978
rect 25261 17926 25313 17978
rect 25325 17926 25377 17978
rect 25389 17926 25441 17978
rect 25453 17926 25505 17978
rect 25517 17926 25569 17978
rect 2780 17731 2832 17740
rect 2780 17697 2789 17731
rect 2789 17697 2823 17731
rect 2823 17697 2832 17731
rect 2780 17688 2832 17697
rect 1584 17663 1636 17672
rect 1584 17629 1593 17663
rect 1593 17629 1627 17663
rect 1627 17629 1636 17663
rect 1584 17620 1636 17629
rect 16120 17824 16172 17876
rect 18696 17824 18748 17876
rect 21640 17824 21692 17876
rect 23112 17824 23164 17876
rect 23848 17824 23900 17876
rect 24032 17824 24084 17876
rect 14648 17756 14700 17808
rect 14740 17756 14792 17808
rect 16212 17688 16264 17740
rect 20168 17688 20220 17740
rect 23204 17731 23256 17740
rect 23204 17697 23213 17731
rect 23213 17697 23247 17731
rect 23247 17697 23256 17731
rect 23204 17688 23256 17697
rect 23388 17731 23440 17740
rect 23388 17697 23397 17731
rect 23397 17697 23431 17731
rect 23431 17697 23440 17731
rect 23388 17688 23440 17697
rect 13728 17663 13780 17672
rect 13728 17629 13737 17663
rect 13737 17629 13771 17663
rect 13771 17629 13780 17663
rect 13728 17620 13780 17629
rect 13820 17620 13872 17672
rect 14740 17663 14792 17672
rect 14740 17629 14749 17663
rect 14749 17629 14783 17663
rect 14783 17629 14792 17663
rect 14740 17620 14792 17629
rect 15844 17620 15896 17672
rect 2412 17552 2464 17604
rect 7748 17484 7800 17536
rect 16580 17552 16632 17604
rect 18788 17663 18840 17672
rect 18788 17629 18797 17663
rect 18797 17629 18831 17663
rect 18831 17629 18840 17663
rect 18788 17620 18840 17629
rect 19892 17620 19944 17672
rect 20904 17620 20956 17672
rect 22560 17663 22612 17672
rect 22560 17629 22569 17663
rect 22569 17629 22603 17663
rect 22603 17629 22612 17663
rect 22560 17620 22612 17629
rect 23112 17620 23164 17672
rect 27896 17756 27948 17808
rect 23848 17620 23900 17672
rect 19800 17552 19852 17604
rect 20076 17527 20128 17536
rect 20076 17493 20085 17527
rect 20085 17493 20119 17527
rect 20119 17493 20128 17527
rect 20076 17484 20128 17493
rect 23388 17552 23440 17604
rect 26700 17731 26752 17740
rect 26700 17697 26709 17731
rect 26709 17697 26743 17731
rect 26743 17697 26752 17731
rect 26700 17688 26752 17697
rect 28632 17688 28684 17740
rect 20260 17484 20312 17536
rect 22652 17484 22704 17536
rect 23480 17484 23532 17536
rect 24584 17527 24636 17536
rect 24584 17493 24593 17527
rect 24593 17493 24627 17527
rect 24627 17493 24636 17527
rect 24584 17484 24636 17493
rect 25504 17484 25556 17536
rect 7896 17382 7948 17434
rect 7960 17382 8012 17434
rect 8024 17382 8076 17434
rect 8088 17382 8140 17434
rect 8152 17382 8204 17434
rect 14842 17382 14894 17434
rect 14906 17382 14958 17434
rect 14970 17382 15022 17434
rect 15034 17382 15086 17434
rect 15098 17382 15150 17434
rect 21788 17382 21840 17434
rect 21852 17382 21904 17434
rect 21916 17382 21968 17434
rect 21980 17382 22032 17434
rect 22044 17382 22096 17434
rect 28734 17382 28786 17434
rect 28798 17382 28850 17434
rect 28862 17382 28914 17434
rect 28926 17382 28978 17434
rect 28990 17382 29042 17434
rect 2412 17323 2464 17332
rect 2412 17289 2421 17323
rect 2421 17289 2455 17323
rect 2455 17289 2464 17323
rect 2412 17280 2464 17289
rect 15752 17323 15804 17332
rect 15752 17289 15761 17323
rect 15761 17289 15795 17323
rect 15795 17289 15804 17323
rect 15752 17280 15804 17289
rect 20076 17280 20128 17332
rect 23020 17280 23072 17332
rect 14004 17212 14056 17264
rect 1584 17144 1636 17196
rect 2504 17187 2556 17196
rect 2504 17153 2513 17187
rect 2513 17153 2547 17187
rect 2547 17153 2556 17187
rect 2504 17144 2556 17153
rect 4344 17144 4396 17196
rect 14556 17187 14608 17196
rect 14556 17153 14565 17187
rect 14565 17153 14599 17187
rect 14599 17153 14608 17187
rect 14556 17144 14608 17153
rect 15844 17144 15896 17196
rect 18052 17187 18104 17196
rect 18052 17153 18061 17187
rect 18061 17153 18095 17187
rect 18095 17153 18104 17187
rect 18052 17144 18104 17153
rect 18328 17255 18380 17264
rect 18328 17221 18362 17255
rect 18362 17221 18380 17255
rect 18328 17212 18380 17221
rect 22192 17212 22244 17264
rect 22560 17255 22612 17264
rect 22560 17221 22569 17255
rect 22569 17221 22603 17255
rect 22603 17221 22612 17255
rect 22560 17212 22612 17221
rect 22652 17255 22704 17264
rect 22652 17221 22661 17255
rect 22661 17221 22695 17255
rect 22695 17221 22704 17255
rect 24124 17280 24176 17332
rect 25504 17323 25556 17332
rect 25504 17289 25513 17323
rect 25513 17289 25547 17323
rect 25547 17289 25556 17323
rect 25504 17280 25556 17289
rect 22652 17212 22704 17221
rect 21640 17144 21692 17196
rect 25044 17212 25096 17264
rect 24400 17187 24452 17196
rect 24400 17153 24434 17187
rect 24434 17153 24452 17187
rect 24400 17144 24452 17153
rect 26240 17187 26292 17196
rect 26240 17153 26249 17187
rect 26249 17153 26283 17187
rect 26283 17153 26292 17187
rect 26240 17144 26292 17153
rect 16580 17076 16632 17128
rect 19984 17076 20036 17128
rect 20444 17119 20496 17128
rect 20444 17085 20453 17119
rect 20453 17085 20487 17119
rect 20487 17085 20496 17119
rect 20444 17076 20496 17085
rect 14556 17051 14608 17060
rect 14556 17017 14565 17051
rect 14565 17017 14599 17051
rect 14599 17017 14608 17051
rect 14556 17008 14608 17017
rect 14740 17008 14792 17060
rect 19800 17008 19852 17060
rect 28264 17144 28316 17196
rect 20536 16940 20588 16992
rect 25872 16940 25924 16992
rect 26700 16940 26752 16992
rect 27896 16983 27948 16992
rect 27896 16949 27905 16983
rect 27905 16949 27939 16983
rect 27939 16949 27948 16983
rect 27896 16940 27948 16949
rect 4423 16838 4475 16890
rect 4487 16838 4539 16890
rect 4551 16838 4603 16890
rect 4615 16838 4667 16890
rect 4679 16838 4731 16890
rect 11369 16838 11421 16890
rect 11433 16838 11485 16890
rect 11497 16838 11549 16890
rect 11561 16838 11613 16890
rect 11625 16838 11677 16890
rect 18315 16838 18367 16890
rect 18379 16838 18431 16890
rect 18443 16838 18495 16890
rect 18507 16838 18559 16890
rect 18571 16838 18623 16890
rect 25261 16838 25313 16890
rect 25325 16838 25377 16890
rect 25389 16838 25441 16890
rect 25453 16838 25505 16890
rect 25517 16838 25569 16890
rect 15660 16736 15712 16788
rect 16580 16736 16632 16788
rect 17684 16736 17736 16788
rect 17960 16736 18012 16788
rect 24952 16711 25004 16720
rect 1676 16532 1728 16584
rect 19248 16532 19300 16584
rect 21456 16532 21508 16584
rect 24952 16677 24961 16711
rect 24961 16677 24995 16711
rect 24995 16677 25004 16711
rect 24952 16668 25004 16677
rect 23848 16600 23900 16652
rect 27896 16668 27948 16720
rect 26700 16643 26752 16652
rect 26700 16609 26709 16643
rect 26709 16609 26743 16643
rect 26743 16609 26752 16643
rect 26700 16600 26752 16609
rect 23020 16575 23072 16584
rect 23020 16541 23029 16575
rect 23029 16541 23063 16575
rect 23063 16541 23072 16575
rect 23020 16532 23072 16541
rect 23480 16575 23532 16584
rect 15844 16464 15896 16516
rect 17040 16464 17092 16516
rect 18880 16464 18932 16516
rect 20720 16464 20772 16516
rect 23480 16541 23489 16575
rect 23489 16541 23523 16575
rect 23523 16541 23532 16575
rect 23480 16532 23532 16541
rect 24584 16464 24636 16516
rect 25872 16464 25924 16516
rect 26240 16464 26292 16516
rect 28632 16464 28684 16516
rect 22560 16396 22612 16448
rect 23664 16439 23716 16448
rect 23664 16405 23673 16439
rect 23673 16405 23707 16439
rect 23707 16405 23716 16439
rect 23664 16396 23716 16405
rect 7896 16294 7948 16346
rect 7960 16294 8012 16346
rect 8024 16294 8076 16346
rect 8088 16294 8140 16346
rect 8152 16294 8204 16346
rect 14842 16294 14894 16346
rect 14906 16294 14958 16346
rect 14970 16294 15022 16346
rect 15034 16294 15086 16346
rect 15098 16294 15150 16346
rect 21788 16294 21840 16346
rect 21852 16294 21904 16346
rect 21916 16294 21968 16346
rect 21980 16294 22032 16346
rect 22044 16294 22096 16346
rect 28734 16294 28786 16346
rect 28798 16294 28850 16346
rect 28862 16294 28914 16346
rect 28926 16294 28978 16346
rect 28990 16294 29042 16346
rect 11980 16192 12032 16244
rect 1676 16099 1728 16108
rect 1676 16065 1685 16099
rect 1685 16065 1719 16099
rect 1719 16065 1728 16099
rect 1676 16056 1728 16065
rect 18052 16124 18104 16176
rect 20720 16192 20772 16244
rect 26240 16192 26292 16244
rect 24860 16124 24912 16176
rect 17132 16099 17184 16108
rect 17132 16065 17166 16099
rect 17166 16065 17184 16099
rect 17132 16056 17184 16065
rect 21272 16099 21324 16108
rect 21272 16065 21281 16099
rect 21281 16065 21315 16099
rect 21315 16065 21324 16099
rect 21272 16056 21324 16065
rect 21456 16099 21508 16108
rect 21456 16065 21465 16099
rect 21465 16065 21499 16099
rect 21499 16065 21508 16099
rect 21456 16056 21508 16065
rect 26240 16099 26292 16108
rect 26240 16065 26249 16099
rect 26249 16065 26283 16099
rect 26283 16065 26292 16099
rect 26240 16056 26292 16065
rect 29920 16056 29972 16108
rect 2228 15988 2280 16040
rect 2780 16031 2832 16040
rect 2780 15997 2789 16031
rect 2789 15997 2823 16031
rect 2823 15997 2832 16031
rect 2780 15988 2832 15997
rect 25964 15988 26016 16040
rect 17224 15852 17276 15904
rect 27160 15895 27212 15904
rect 27160 15861 27169 15895
rect 27169 15861 27203 15895
rect 27203 15861 27212 15895
rect 27160 15852 27212 15861
rect 4423 15750 4475 15802
rect 4487 15750 4539 15802
rect 4551 15750 4603 15802
rect 4615 15750 4667 15802
rect 4679 15750 4731 15802
rect 11369 15750 11421 15802
rect 11433 15750 11485 15802
rect 11497 15750 11549 15802
rect 11561 15750 11613 15802
rect 11625 15750 11677 15802
rect 18315 15750 18367 15802
rect 18379 15750 18431 15802
rect 18443 15750 18495 15802
rect 18507 15750 18559 15802
rect 18571 15750 18623 15802
rect 25261 15750 25313 15802
rect 25325 15750 25377 15802
rect 25389 15750 25441 15802
rect 25453 15750 25505 15802
rect 25517 15750 25569 15802
rect 2228 15691 2280 15700
rect 2228 15657 2237 15691
rect 2237 15657 2271 15691
rect 2271 15657 2280 15691
rect 2228 15648 2280 15657
rect 20812 15691 20864 15700
rect 20812 15657 20821 15691
rect 20821 15657 20855 15691
rect 20855 15657 20864 15691
rect 20812 15648 20864 15657
rect 13452 15512 13504 15564
rect 21640 15555 21692 15564
rect 21640 15521 21649 15555
rect 21649 15521 21683 15555
rect 21683 15521 21692 15555
rect 21640 15512 21692 15521
rect 25044 15512 25096 15564
rect 26056 15512 26108 15564
rect 2320 15487 2372 15496
rect 2320 15453 2329 15487
rect 2329 15453 2363 15487
rect 2363 15453 2372 15487
rect 2320 15444 2372 15453
rect 10692 15487 10744 15496
rect 10692 15453 10701 15487
rect 10701 15453 10735 15487
rect 10735 15453 10744 15487
rect 10692 15444 10744 15453
rect 11060 15376 11112 15428
rect 18052 15444 18104 15496
rect 19248 15444 19300 15496
rect 25504 15487 25556 15496
rect 25504 15453 25513 15487
rect 25513 15453 25547 15487
rect 25547 15453 25556 15487
rect 25504 15444 25556 15453
rect 27160 15444 27212 15496
rect 28080 15444 28132 15496
rect 11980 15376 12032 15428
rect 17316 15376 17368 15428
rect 19708 15419 19760 15428
rect 19708 15385 19742 15419
rect 19742 15385 19760 15419
rect 19708 15376 19760 15385
rect 21548 15376 21600 15428
rect 18696 15308 18748 15360
rect 23020 15351 23072 15360
rect 23020 15317 23029 15351
rect 23029 15317 23063 15351
rect 23063 15317 23072 15351
rect 23020 15308 23072 15317
rect 27344 15308 27396 15360
rect 27436 15308 27488 15360
rect 28172 15308 28224 15360
rect 7896 15206 7948 15258
rect 7960 15206 8012 15258
rect 8024 15206 8076 15258
rect 8088 15206 8140 15258
rect 8152 15206 8204 15258
rect 14842 15206 14894 15258
rect 14906 15206 14958 15258
rect 14970 15206 15022 15258
rect 15034 15206 15086 15258
rect 15098 15206 15150 15258
rect 21788 15206 21840 15258
rect 21852 15206 21904 15258
rect 21916 15206 21968 15258
rect 21980 15206 22032 15258
rect 22044 15206 22096 15258
rect 28734 15206 28786 15258
rect 28798 15206 28850 15258
rect 28862 15206 28914 15258
rect 28926 15206 28978 15258
rect 28990 15206 29042 15258
rect 20444 15104 20496 15156
rect 20628 15104 20680 15156
rect 19248 15036 19300 15088
rect 21272 15104 21324 15156
rect 22560 15104 22612 15156
rect 23112 15104 23164 15156
rect 26240 15104 26292 15156
rect 27344 15104 27396 15156
rect 17960 15011 18012 15020
rect 17960 14977 17978 15011
rect 17978 14977 18012 15011
rect 17960 14968 18012 14977
rect 18144 14968 18196 15020
rect 20352 15011 20404 15020
rect 20352 14977 20370 15011
rect 20370 14977 20404 15011
rect 20352 14968 20404 14977
rect 23664 15036 23716 15088
rect 26056 15036 26108 15088
rect 25044 14968 25096 15020
rect 25136 14968 25188 15020
rect 27436 14968 27488 15020
rect 19340 14832 19392 14884
rect 27344 14900 27396 14952
rect 22744 14832 22796 14884
rect 23296 14832 23348 14884
rect 16212 14764 16264 14816
rect 21456 14764 21508 14816
rect 24216 14764 24268 14816
rect 4423 14662 4475 14714
rect 4487 14662 4539 14714
rect 4551 14662 4603 14714
rect 4615 14662 4667 14714
rect 4679 14662 4731 14714
rect 11369 14662 11421 14714
rect 11433 14662 11485 14714
rect 11497 14662 11549 14714
rect 11561 14662 11613 14714
rect 11625 14662 11677 14714
rect 18315 14662 18367 14714
rect 18379 14662 18431 14714
rect 18443 14662 18495 14714
rect 18507 14662 18559 14714
rect 18571 14662 18623 14714
rect 25261 14662 25313 14714
rect 25325 14662 25377 14714
rect 25389 14662 25441 14714
rect 25453 14662 25505 14714
rect 25517 14662 25569 14714
rect 17960 14560 18012 14612
rect 19708 14560 19760 14612
rect 3424 14399 3476 14408
rect 3424 14365 3433 14399
rect 3433 14365 3467 14399
rect 3467 14365 3476 14399
rect 3424 14356 3476 14365
rect 15660 14356 15712 14408
rect 16120 14356 16172 14408
rect 1584 14331 1636 14340
rect 1584 14297 1593 14331
rect 1593 14297 1627 14331
rect 1627 14297 1636 14331
rect 1584 14288 1636 14297
rect 2872 14288 2924 14340
rect 16212 14331 16264 14340
rect 16212 14297 16221 14331
rect 16221 14297 16255 14331
rect 16255 14297 16264 14331
rect 16212 14288 16264 14297
rect 16856 14331 16908 14340
rect 16856 14297 16865 14331
rect 16865 14297 16899 14331
rect 16899 14297 16908 14331
rect 16856 14288 16908 14297
rect 16304 14220 16356 14272
rect 17408 14424 17460 14476
rect 26056 14467 26108 14476
rect 26056 14433 26065 14467
rect 26065 14433 26099 14467
rect 26099 14433 26108 14467
rect 26056 14424 26108 14433
rect 27528 14467 27580 14476
rect 27528 14433 27537 14467
rect 27537 14433 27571 14467
rect 27571 14433 27580 14467
rect 27528 14424 27580 14433
rect 28172 14467 28224 14476
rect 28172 14433 28181 14467
rect 28181 14433 28215 14467
rect 28215 14433 28224 14467
rect 28172 14424 28224 14433
rect 19432 14399 19484 14408
rect 19432 14365 19441 14399
rect 19441 14365 19475 14399
rect 19475 14365 19484 14399
rect 19432 14356 19484 14365
rect 28356 14399 28408 14408
rect 28356 14365 28365 14399
rect 28365 14365 28399 14399
rect 28399 14365 28408 14399
rect 28356 14356 28408 14365
rect 25780 14331 25832 14340
rect 25780 14297 25798 14331
rect 25798 14297 25832 14331
rect 25780 14288 25832 14297
rect 24308 14220 24360 14272
rect 26240 14220 26292 14272
rect 7896 14118 7948 14170
rect 7960 14118 8012 14170
rect 8024 14118 8076 14170
rect 8088 14118 8140 14170
rect 8152 14118 8204 14170
rect 14842 14118 14894 14170
rect 14906 14118 14958 14170
rect 14970 14118 15022 14170
rect 15034 14118 15086 14170
rect 15098 14118 15150 14170
rect 21788 14118 21840 14170
rect 21852 14118 21904 14170
rect 21916 14118 21968 14170
rect 21980 14118 22032 14170
rect 22044 14118 22096 14170
rect 28734 14118 28786 14170
rect 28798 14118 28850 14170
rect 28862 14118 28914 14170
rect 28926 14118 28978 14170
rect 28990 14118 29042 14170
rect 2872 14059 2924 14068
rect 2872 14025 2881 14059
rect 2881 14025 2915 14059
rect 2915 14025 2924 14059
rect 2872 14016 2924 14025
rect 16304 14059 16356 14068
rect 16304 14025 16313 14059
rect 16313 14025 16347 14059
rect 16347 14025 16356 14059
rect 16304 14016 16356 14025
rect 17316 14016 17368 14068
rect 19432 14059 19484 14068
rect 19432 14025 19441 14059
rect 19441 14025 19475 14059
rect 19475 14025 19484 14059
rect 19432 14016 19484 14025
rect 20352 14016 20404 14068
rect 22744 14016 22796 14068
rect 23480 14016 23532 14068
rect 23756 14016 23808 14068
rect 24032 14016 24084 14068
rect 25136 14016 25188 14068
rect 25780 14059 25832 14068
rect 25780 14025 25789 14059
rect 25789 14025 25823 14059
rect 25823 14025 25832 14059
rect 25780 14016 25832 14025
rect 3424 13948 3476 14000
rect 23020 13948 23072 14000
rect 2964 13923 3016 13932
rect 2964 13889 2973 13923
rect 2973 13889 3007 13923
rect 3007 13889 3016 13923
rect 2964 13880 3016 13889
rect 16120 13923 16172 13932
rect 16120 13889 16129 13923
rect 16129 13889 16163 13923
rect 16163 13889 16172 13923
rect 16120 13880 16172 13889
rect 16212 13880 16264 13932
rect 16856 13855 16908 13864
rect 16856 13821 16865 13855
rect 16865 13821 16899 13855
rect 16899 13821 16908 13855
rect 16856 13812 16908 13821
rect 17040 13880 17092 13932
rect 17408 13880 17460 13932
rect 18696 13880 18748 13932
rect 19616 13923 19668 13932
rect 19616 13889 19625 13923
rect 19625 13889 19659 13923
rect 19659 13889 19668 13923
rect 19616 13880 19668 13889
rect 19892 13880 19944 13932
rect 20444 13923 20496 13932
rect 20444 13889 20453 13923
rect 20453 13889 20487 13923
rect 20487 13889 20496 13923
rect 20444 13880 20496 13889
rect 23756 13923 23808 13932
rect 23756 13889 23765 13923
rect 23765 13889 23799 13923
rect 23799 13889 23808 13923
rect 23756 13880 23808 13889
rect 21640 13812 21692 13864
rect 22468 13855 22520 13864
rect 22468 13821 22477 13855
rect 22477 13821 22511 13855
rect 22511 13821 22520 13855
rect 22468 13812 22520 13821
rect 23664 13812 23716 13864
rect 24216 13880 24268 13932
rect 24584 13923 24636 13932
rect 24584 13889 24593 13923
rect 24593 13889 24627 13923
rect 24627 13889 24636 13923
rect 24584 13880 24636 13889
rect 25596 13923 25648 13932
rect 25596 13889 25605 13923
rect 25605 13889 25639 13923
rect 25639 13889 25648 13923
rect 25596 13880 25648 13889
rect 28356 13880 28408 13932
rect 18144 13744 18196 13796
rect 22284 13744 22336 13796
rect 3424 13719 3476 13728
rect 3424 13685 3433 13719
rect 3433 13685 3467 13719
rect 3467 13685 3476 13719
rect 3424 13676 3476 13685
rect 17960 13719 18012 13728
rect 17960 13685 17969 13719
rect 17969 13685 18003 13719
rect 18003 13685 18012 13719
rect 17960 13676 18012 13685
rect 18052 13676 18104 13728
rect 24308 13744 24360 13796
rect 23112 13719 23164 13728
rect 23112 13685 23121 13719
rect 23121 13685 23155 13719
rect 23155 13685 23164 13719
rect 23112 13676 23164 13685
rect 23296 13719 23348 13728
rect 23296 13685 23305 13719
rect 23305 13685 23339 13719
rect 23339 13685 23348 13719
rect 23296 13676 23348 13685
rect 24676 13676 24728 13728
rect 4423 13574 4475 13626
rect 4487 13574 4539 13626
rect 4551 13574 4603 13626
rect 4615 13574 4667 13626
rect 4679 13574 4731 13626
rect 11369 13574 11421 13626
rect 11433 13574 11485 13626
rect 11497 13574 11549 13626
rect 11561 13574 11613 13626
rect 11625 13574 11677 13626
rect 18315 13574 18367 13626
rect 18379 13574 18431 13626
rect 18443 13574 18495 13626
rect 18507 13574 18559 13626
rect 18571 13574 18623 13626
rect 25261 13574 25313 13626
rect 25325 13574 25377 13626
rect 25389 13574 25441 13626
rect 25453 13574 25505 13626
rect 25517 13574 25569 13626
rect 18052 13515 18104 13524
rect 18052 13481 18061 13515
rect 18061 13481 18095 13515
rect 18095 13481 18104 13515
rect 18052 13472 18104 13481
rect 19616 13472 19668 13524
rect 22284 13515 22336 13524
rect 22284 13481 22293 13515
rect 22293 13481 22327 13515
rect 22327 13481 22336 13515
rect 22284 13472 22336 13481
rect 23296 13472 23348 13524
rect 24584 13515 24636 13524
rect 1584 13379 1636 13388
rect 1584 13345 1593 13379
rect 1593 13345 1627 13379
rect 1627 13345 1636 13379
rect 1584 13336 1636 13345
rect 3424 13379 3476 13388
rect 3424 13345 3433 13379
rect 3433 13345 3467 13379
rect 3467 13345 3476 13379
rect 3424 13336 3476 13345
rect 20628 13336 20680 13388
rect 17040 13268 17092 13320
rect 18144 13268 18196 13320
rect 1952 13200 2004 13252
rect 18328 13311 18380 13320
rect 18328 13277 18337 13311
rect 18337 13277 18371 13311
rect 18371 13277 18380 13311
rect 18328 13268 18380 13277
rect 18972 13268 19024 13320
rect 20812 13268 20864 13320
rect 21456 13311 21508 13320
rect 21456 13277 21465 13311
rect 21465 13277 21499 13311
rect 21499 13277 21508 13311
rect 21456 13268 21508 13277
rect 23020 13336 23072 13388
rect 23664 13404 23716 13456
rect 24584 13481 24593 13515
rect 24593 13481 24627 13515
rect 24627 13481 24636 13515
rect 24584 13472 24636 13481
rect 24676 13472 24728 13524
rect 25596 13515 25648 13524
rect 25596 13481 25605 13515
rect 25605 13481 25639 13515
rect 25639 13481 25648 13515
rect 25596 13472 25648 13481
rect 23572 13311 23624 13320
rect 23112 13200 23164 13252
rect 23572 13277 23581 13311
rect 23581 13277 23615 13311
rect 23615 13277 23624 13311
rect 23572 13268 23624 13277
rect 23480 13200 23532 13252
rect 17960 13132 18012 13184
rect 18788 13132 18840 13184
rect 21088 13175 21140 13184
rect 21088 13141 21097 13175
rect 21097 13141 21131 13175
rect 21131 13141 21140 13175
rect 21088 13132 21140 13141
rect 22744 13175 22796 13184
rect 22744 13141 22753 13175
rect 22753 13141 22787 13175
rect 22787 13141 22796 13175
rect 22744 13132 22796 13141
rect 22836 13175 22888 13184
rect 22836 13141 22845 13175
rect 22845 13141 22879 13175
rect 22879 13141 22888 13175
rect 24032 13268 24084 13320
rect 25872 13268 25924 13320
rect 25964 13311 26016 13320
rect 25964 13277 25973 13311
rect 25973 13277 26007 13311
rect 26007 13277 26016 13311
rect 25964 13268 26016 13277
rect 24952 13243 25004 13252
rect 24952 13209 24961 13243
rect 24961 13209 24995 13243
rect 24995 13209 25004 13243
rect 24952 13200 25004 13209
rect 22836 13132 22888 13141
rect 7896 13030 7948 13082
rect 7960 13030 8012 13082
rect 8024 13030 8076 13082
rect 8088 13030 8140 13082
rect 8152 13030 8204 13082
rect 14842 13030 14894 13082
rect 14906 13030 14958 13082
rect 14970 13030 15022 13082
rect 15034 13030 15086 13082
rect 15098 13030 15150 13082
rect 21788 13030 21840 13082
rect 21852 13030 21904 13082
rect 21916 13030 21968 13082
rect 21980 13030 22032 13082
rect 22044 13030 22096 13082
rect 28734 13030 28786 13082
rect 28798 13030 28850 13082
rect 28862 13030 28914 13082
rect 28926 13030 28978 13082
rect 28990 13030 29042 13082
rect 1952 12971 2004 12980
rect 1952 12937 1961 12971
rect 1961 12937 1995 12971
rect 1995 12937 2004 12971
rect 1952 12928 2004 12937
rect 20444 12928 20496 12980
rect 22468 12928 22520 12980
rect 23756 12971 23808 12980
rect 2044 12835 2096 12844
rect 2044 12801 2053 12835
rect 2053 12801 2087 12835
rect 2087 12801 2096 12835
rect 2044 12792 2096 12801
rect 4988 12792 5040 12844
rect 16672 12792 16724 12844
rect 18052 12792 18104 12844
rect 18880 12792 18932 12844
rect 19892 12792 19944 12844
rect 20168 12835 20220 12844
rect 20168 12801 20177 12835
rect 20177 12801 20211 12835
rect 20211 12801 20220 12835
rect 20168 12792 20220 12801
rect 21088 12792 21140 12844
rect 23756 12937 23765 12971
rect 23765 12937 23799 12971
rect 23799 12937 23808 12971
rect 23756 12928 23808 12937
rect 25872 12971 25924 12980
rect 25872 12937 25881 12971
rect 25881 12937 25915 12971
rect 25915 12937 25924 12971
rect 25872 12928 25924 12937
rect 26240 12971 26292 12980
rect 26240 12937 26249 12971
rect 26249 12937 26283 12971
rect 26283 12937 26292 12971
rect 26240 12928 26292 12937
rect 23296 12860 23348 12912
rect 23940 12860 23992 12912
rect 23480 12792 23532 12844
rect 26976 12792 27028 12844
rect 27620 12792 27672 12844
rect 16948 12724 17000 12776
rect 22744 12767 22796 12776
rect 22744 12733 22753 12767
rect 22753 12733 22787 12767
rect 22787 12733 22796 12767
rect 22744 12724 22796 12733
rect 23848 12724 23900 12776
rect 17500 12656 17552 12708
rect 27344 12724 27396 12776
rect 26516 12656 26568 12708
rect 18236 12631 18288 12640
rect 18236 12597 18245 12631
rect 18245 12597 18279 12631
rect 18279 12597 18288 12631
rect 18236 12588 18288 12597
rect 18696 12588 18748 12640
rect 20260 12588 20312 12640
rect 26700 12588 26752 12640
rect 4423 12486 4475 12538
rect 4487 12486 4539 12538
rect 4551 12486 4603 12538
rect 4615 12486 4667 12538
rect 4679 12486 4731 12538
rect 11369 12486 11421 12538
rect 11433 12486 11485 12538
rect 11497 12486 11549 12538
rect 11561 12486 11613 12538
rect 11625 12486 11677 12538
rect 18315 12486 18367 12538
rect 18379 12486 18431 12538
rect 18443 12486 18495 12538
rect 18507 12486 18559 12538
rect 18571 12486 18623 12538
rect 25261 12486 25313 12538
rect 25325 12486 25377 12538
rect 25389 12486 25441 12538
rect 25453 12486 25505 12538
rect 25517 12486 25569 12538
rect 3516 12384 3568 12436
rect 11060 12384 11112 12436
rect 17132 12384 17184 12436
rect 21548 12384 21600 12436
rect 20168 12248 20220 12300
rect 1676 12223 1728 12232
rect 1676 12189 1685 12223
rect 1685 12189 1719 12223
rect 1719 12189 1728 12223
rect 1676 12180 1728 12189
rect 16672 12223 16724 12232
rect 16672 12189 16681 12223
rect 16681 12189 16715 12223
rect 16715 12189 16724 12223
rect 16672 12180 16724 12189
rect 24952 12248 25004 12300
rect 26516 12291 26568 12300
rect 26516 12257 26525 12291
rect 26525 12257 26559 12291
rect 26559 12257 26568 12291
rect 26516 12248 26568 12257
rect 26700 12291 26752 12300
rect 26700 12257 26709 12291
rect 26709 12257 26743 12291
rect 26743 12257 26752 12291
rect 26700 12248 26752 12257
rect 28356 12291 28408 12300
rect 28356 12257 28365 12291
rect 28365 12257 28399 12291
rect 28399 12257 28408 12291
rect 28356 12248 28408 12257
rect 21640 12180 21692 12232
rect 7896 11942 7948 11994
rect 7960 11942 8012 11994
rect 8024 11942 8076 11994
rect 8088 11942 8140 11994
rect 8152 11942 8204 11994
rect 14842 11942 14894 11994
rect 14906 11942 14958 11994
rect 14970 11942 15022 11994
rect 15034 11942 15086 11994
rect 15098 11942 15150 11994
rect 21788 11942 21840 11994
rect 21852 11942 21904 11994
rect 21916 11942 21968 11994
rect 21980 11942 22032 11994
rect 22044 11942 22096 11994
rect 28734 11942 28786 11994
rect 28798 11942 28850 11994
rect 28862 11942 28914 11994
rect 28926 11942 28978 11994
rect 28990 11942 29042 11994
rect 16672 11840 16724 11892
rect 18880 11840 18932 11892
rect 18236 11815 18288 11824
rect 18236 11781 18245 11815
rect 18245 11781 18279 11815
rect 18279 11781 18288 11815
rect 18236 11772 18288 11781
rect 1676 11747 1728 11756
rect 1676 11713 1685 11747
rect 1685 11713 1719 11747
rect 1719 11713 1728 11747
rect 1676 11704 1728 11713
rect 17224 11747 17276 11756
rect 17224 11713 17233 11747
rect 17233 11713 17267 11747
rect 17267 11713 17276 11747
rect 17224 11704 17276 11713
rect 18052 11704 18104 11756
rect 18788 11747 18840 11756
rect 18788 11713 18797 11747
rect 18797 11713 18831 11747
rect 18831 11713 18840 11747
rect 18788 11704 18840 11713
rect 27068 11704 27120 11756
rect 1860 11679 1912 11688
rect 1860 11645 1869 11679
rect 1869 11645 1903 11679
rect 1903 11645 1912 11679
rect 1860 11636 1912 11645
rect 2780 11679 2832 11688
rect 2780 11645 2789 11679
rect 2789 11645 2823 11679
rect 2823 11645 2832 11679
rect 2780 11636 2832 11645
rect 17500 11679 17552 11688
rect 17500 11645 17509 11679
rect 17509 11645 17543 11679
rect 17543 11645 17552 11679
rect 17500 11636 17552 11645
rect 18880 11679 18932 11688
rect 18880 11645 18889 11679
rect 18889 11645 18923 11679
rect 18923 11645 18932 11679
rect 18880 11636 18932 11645
rect 26700 11500 26752 11552
rect 4423 11398 4475 11450
rect 4487 11398 4539 11450
rect 4551 11398 4603 11450
rect 4615 11398 4667 11450
rect 4679 11398 4731 11450
rect 11369 11398 11421 11450
rect 11433 11398 11485 11450
rect 11497 11398 11549 11450
rect 11561 11398 11613 11450
rect 11625 11398 11677 11450
rect 18315 11398 18367 11450
rect 18379 11398 18431 11450
rect 18443 11398 18495 11450
rect 18507 11398 18559 11450
rect 18571 11398 18623 11450
rect 25261 11398 25313 11450
rect 25325 11398 25377 11450
rect 25389 11398 25441 11450
rect 25453 11398 25505 11450
rect 25517 11398 25569 11450
rect 1860 11339 1912 11348
rect 1860 11305 1869 11339
rect 1869 11305 1903 11339
rect 1903 11305 1912 11339
rect 1860 11296 1912 11305
rect 18788 11296 18840 11348
rect 19156 11296 19208 11348
rect 4344 11203 4396 11212
rect 4344 11169 4353 11203
rect 4353 11169 4387 11203
rect 4387 11169 4396 11203
rect 4344 11160 4396 11169
rect 26700 11203 26752 11212
rect 26700 11169 26709 11203
rect 26709 11169 26743 11203
rect 26743 11169 26752 11203
rect 26700 11160 26752 11169
rect 1492 11092 1544 11144
rect 2964 11092 3016 11144
rect 17684 11135 17736 11144
rect 17684 11101 17693 11135
rect 17693 11101 17727 11135
rect 17727 11101 17736 11135
rect 17684 11092 17736 11101
rect 26516 11135 26568 11144
rect 26516 11101 26525 11135
rect 26525 11101 26559 11135
rect 26559 11101 26568 11135
rect 26516 11092 26568 11101
rect 18328 11024 18380 11076
rect 29920 11024 29972 11076
rect 17776 10999 17828 11008
rect 17776 10965 17785 10999
rect 17785 10965 17819 10999
rect 17819 10965 17828 10999
rect 17776 10956 17828 10965
rect 19248 10956 19300 11008
rect 7896 10854 7948 10906
rect 7960 10854 8012 10906
rect 8024 10854 8076 10906
rect 8088 10854 8140 10906
rect 8152 10854 8204 10906
rect 14842 10854 14894 10906
rect 14906 10854 14958 10906
rect 14970 10854 15022 10906
rect 15034 10854 15086 10906
rect 15098 10854 15150 10906
rect 21788 10854 21840 10906
rect 21852 10854 21904 10906
rect 21916 10854 21968 10906
rect 21980 10854 22032 10906
rect 22044 10854 22096 10906
rect 28734 10854 28786 10906
rect 28798 10854 28850 10906
rect 28862 10854 28914 10906
rect 28926 10854 28978 10906
rect 28990 10854 29042 10906
rect 18236 10795 18288 10804
rect 18236 10761 18245 10795
rect 18245 10761 18279 10795
rect 18279 10761 18288 10795
rect 18236 10752 18288 10761
rect 18880 10752 18932 10804
rect 17776 10684 17828 10736
rect 18880 10659 18932 10668
rect 18880 10625 18889 10659
rect 18889 10625 18923 10659
rect 18923 10625 18932 10659
rect 18880 10616 18932 10625
rect 19156 10659 19208 10668
rect 17224 10548 17276 10600
rect 17960 10548 18012 10600
rect 19156 10625 19165 10659
rect 19165 10625 19199 10659
rect 19199 10625 19208 10659
rect 19156 10616 19208 10625
rect 19248 10659 19300 10668
rect 19248 10625 19257 10659
rect 19257 10625 19291 10659
rect 19291 10625 19300 10659
rect 19248 10616 19300 10625
rect 20260 10659 20312 10668
rect 20260 10625 20269 10659
rect 20269 10625 20303 10659
rect 20303 10625 20312 10659
rect 20260 10616 20312 10625
rect 26516 10616 26568 10668
rect 20168 10591 20220 10600
rect 20168 10557 20177 10591
rect 20177 10557 20211 10591
rect 20211 10557 20220 10591
rect 20168 10548 20220 10557
rect 27436 10548 27488 10600
rect 18144 10412 18196 10464
rect 28356 10412 28408 10464
rect 4423 10310 4475 10362
rect 4487 10310 4539 10362
rect 4551 10310 4603 10362
rect 4615 10310 4667 10362
rect 4679 10310 4731 10362
rect 11369 10310 11421 10362
rect 11433 10310 11485 10362
rect 11497 10310 11549 10362
rect 11561 10310 11613 10362
rect 11625 10310 11677 10362
rect 18315 10310 18367 10362
rect 18379 10310 18431 10362
rect 18443 10310 18495 10362
rect 18507 10310 18559 10362
rect 18571 10310 18623 10362
rect 25261 10310 25313 10362
rect 25325 10310 25377 10362
rect 25389 10310 25441 10362
rect 25453 10310 25505 10362
rect 25517 10310 25569 10362
rect 18236 10251 18288 10260
rect 18236 10217 18245 10251
rect 18245 10217 18279 10251
rect 18279 10217 18288 10251
rect 18236 10208 18288 10217
rect 19156 10140 19208 10192
rect 18144 10115 18196 10124
rect 18144 10081 18153 10115
rect 18153 10081 18187 10115
rect 18187 10081 18196 10115
rect 18144 10072 18196 10081
rect 20260 10072 20312 10124
rect 27528 10115 27580 10124
rect 27528 10081 27537 10115
rect 27537 10081 27571 10115
rect 27571 10081 27580 10115
rect 27528 10072 27580 10081
rect 28356 10115 28408 10124
rect 28356 10081 28365 10115
rect 28365 10081 28399 10115
rect 28399 10081 28408 10115
rect 28356 10072 28408 10081
rect 1676 10047 1728 10056
rect 1676 10013 1685 10047
rect 1685 10013 1719 10047
rect 1719 10013 1728 10047
rect 1676 10004 1728 10013
rect 2964 10004 3016 10056
rect 17960 10047 18012 10056
rect 17960 10013 17969 10047
rect 17969 10013 18003 10047
rect 18003 10013 18012 10047
rect 17960 10004 18012 10013
rect 20168 10004 20220 10056
rect 18880 9936 18932 9988
rect 28172 9979 28224 9988
rect 28172 9945 28181 9979
rect 28181 9945 28215 9979
rect 28215 9945 28224 9979
rect 28172 9936 28224 9945
rect 4068 9868 4120 9920
rect 7896 9766 7948 9818
rect 7960 9766 8012 9818
rect 8024 9766 8076 9818
rect 8088 9766 8140 9818
rect 8152 9766 8204 9818
rect 14842 9766 14894 9818
rect 14906 9766 14958 9818
rect 14970 9766 15022 9818
rect 15034 9766 15086 9818
rect 15098 9766 15150 9818
rect 21788 9766 21840 9818
rect 21852 9766 21904 9818
rect 21916 9766 21968 9818
rect 21980 9766 22032 9818
rect 22044 9766 22096 9818
rect 28734 9766 28786 9818
rect 28798 9766 28850 9818
rect 28862 9766 28914 9818
rect 28926 9766 28978 9818
rect 28990 9766 29042 9818
rect 28172 9664 28224 9716
rect 1676 9571 1728 9580
rect 1676 9537 1685 9571
rect 1685 9537 1719 9571
rect 1719 9537 1728 9571
rect 1676 9528 1728 9537
rect 20536 9528 20588 9580
rect 27344 9528 27396 9580
rect 27620 9528 27672 9580
rect 1860 9503 1912 9512
rect 1860 9469 1869 9503
rect 1869 9469 1903 9503
rect 1903 9469 1912 9503
rect 1860 9460 1912 9469
rect 2780 9503 2832 9512
rect 2780 9469 2789 9503
rect 2789 9469 2823 9503
rect 2823 9469 2832 9503
rect 2780 9460 2832 9469
rect 4252 9324 4304 9376
rect 20628 9324 20680 9376
rect 4423 9222 4475 9274
rect 4487 9222 4539 9274
rect 4551 9222 4603 9274
rect 4615 9222 4667 9274
rect 4679 9222 4731 9274
rect 11369 9222 11421 9274
rect 11433 9222 11485 9274
rect 11497 9222 11549 9274
rect 11561 9222 11613 9274
rect 11625 9222 11677 9274
rect 18315 9222 18367 9274
rect 18379 9222 18431 9274
rect 18443 9222 18495 9274
rect 18507 9222 18559 9274
rect 18571 9222 18623 9274
rect 25261 9222 25313 9274
rect 25325 9222 25377 9274
rect 25389 9222 25441 9274
rect 25453 9222 25505 9274
rect 25517 9222 25569 9274
rect 2964 9027 3016 9036
rect 2964 8993 2973 9027
rect 2973 8993 3007 9027
rect 3007 8993 3016 9027
rect 2964 8984 3016 8993
rect 1584 8959 1636 8968
rect 1584 8925 1593 8959
rect 1593 8925 1627 8959
rect 1627 8925 1636 8959
rect 1584 8916 1636 8925
rect 26516 8959 26568 8968
rect 26516 8925 26525 8959
rect 26525 8925 26559 8959
rect 26559 8925 26568 8959
rect 26516 8916 26568 8925
rect 28356 8959 28408 8968
rect 28356 8925 28365 8959
rect 28365 8925 28399 8959
rect 28399 8925 28408 8959
rect 28356 8916 28408 8925
rect 1768 8891 1820 8900
rect 1768 8857 1777 8891
rect 1777 8857 1811 8891
rect 1811 8857 1820 8891
rect 1768 8848 1820 8857
rect 27252 8848 27304 8900
rect 7896 8678 7948 8730
rect 7960 8678 8012 8730
rect 8024 8678 8076 8730
rect 8088 8678 8140 8730
rect 8152 8678 8204 8730
rect 14842 8678 14894 8730
rect 14906 8678 14958 8730
rect 14970 8678 15022 8730
rect 15034 8678 15086 8730
rect 15098 8678 15150 8730
rect 21788 8678 21840 8730
rect 21852 8678 21904 8730
rect 21916 8678 21968 8730
rect 21980 8678 22032 8730
rect 22044 8678 22096 8730
rect 28734 8678 28786 8730
rect 28798 8678 28850 8730
rect 28862 8678 28914 8730
rect 28926 8678 28978 8730
rect 28990 8678 29042 8730
rect 1860 8619 1912 8628
rect 1860 8585 1869 8619
rect 1869 8585 1903 8619
rect 1903 8585 1912 8619
rect 1860 8576 1912 8585
rect 4344 8576 4396 8628
rect 27252 8619 27304 8628
rect 4068 8551 4120 8560
rect 4068 8517 4077 8551
rect 4077 8517 4111 8551
rect 4111 8517 4120 8551
rect 4068 8508 4120 8517
rect 4252 8483 4304 8492
rect 4252 8449 4261 8483
rect 4261 8449 4295 8483
rect 4295 8449 4304 8483
rect 27252 8585 27261 8619
rect 27261 8585 27295 8619
rect 27295 8585 27304 8619
rect 27252 8576 27304 8585
rect 26516 8508 26568 8560
rect 4252 8440 4304 8449
rect 3332 8415 3384 8424
rect 3332 8381 3341 8415
rect 3341 8381 3375 8415
rect 3375 8381 3384 8415
rect 3332 8372 3384 8381
rect 27804 8304 27856 8356
rect 26608 8279 26660 8288
rect 26608 8245 26617 8279
rect 26617 8245 26651 8279
rect 26651 8245 26660 8279
rect 26608 8236 26660 8245
rect 4423 8134 4475 8186
rect 4487 8134 4539 8186
rect 4551 8134 4603 8186
rect 4615 8134 4667 8186
rect 4679 8134 4731 8186
rect 11369 8134 11421 8186
rect 11433 8134 11485 8186
rect 11497 8134 11549 8186
rect 11561 8134 11613 8186
rect 11625 8134 11677 8186
rect 18315 8134 18367 8186
rect 18379 8134 18431 8186
rect 18443 8134 18495 8186
rect 18507 8134 18559 8186
rect 18571 8134 18623 8186
rect 25261 8134 25313 8186
rect 25325 8134 25377 8186
rect 25389 8134 25441 8186
rect 25453 8134 25505 8186
rect 25517 8134 25569 8186
rect 1584 8032 1636 8084
rect 1768 8032 1820 8084
rect 1492 7828 1544 7880
rect 2504 7871 2556 7880
rect 2504 7837 2513 7871
rect 2513 7837 2547 7871
rect 2547 7837 2556 7871
rect 2504 7828 2556 7837
rect 3884 7828 3936 7880
rect 25688 7828 25740 7880
rect 27712 7896 27764 7948
rect 4896 7760 4948 7812
rect 4712 7692 4764 7744
rect 26424 7692 26476 7744
rect 26700 7803 26752 7812
rect 26700 7769 26709 7803
rect 26709 7769 26743 7803
rect 26743 7769 26752 7803
rect 26700 7760 26752 7769
rect 29920 7760 29972 7812
rect 27804 7692 27856 7744
rect 7896 7590 7948 7642
rect 7960 7590 8012 7642
rect 8024 7590 8076 7642
rect 8088 7590 8140 7642
rect 8152 7590 8204 7642
rect 14842 7590 14894 7642
rect 14906 7590 14958 7642
rect 14970 7590 15022 7642
rect 15034 7590 15086 7642
rect 15098 7590 15150 7642
rect 21788 7590 21840 7642
rect 21852 7590 21904 7642
rect 21916 7590 21968 7642
rect 21980 7590 22032 7642
rect 22044 7590 22096 7642
rect 28734 7590 28786 7642
rect 28798 7590 28850 7642
rect 28862 7590 28914 7642
rect 28926 7590 28978 7642
rect 28990 7590 29042 7642
rect 3056 7463 3108 7472
rect 3056 7429 3065 7463
rect 3065 7429 3099 7463
rect 3099 7429 3108 7463
rect 3056 7420 3108 7429
rect 4712 7463 4764 7472
rect 4712 7429 4721 7463
rect 4721 7429 4755 7463
rect 4755 7429 4764 7463
rect 4712 7420 4764 7429
rect 26424 7463 26476 7472
rect 26424 7429 26433 7463
rect 26433 7429 26467 7463
rect 26467 7429 26476 7463
rect 26424 7420 26476 7429
rect 4896 7395 4948 7404
rect 4896 7361 4905 7395
rect 4905 7361 4939 7395
rect 4939 7361 4948 7395
rect 4896 7352 4948 7361
rect 26608 7395 26660 7404
rect 26608 7361 26617 7395
rect 26617 7361 26651 7395
rect 26651 7361 26660 7395
rect 27804 7395 27856 7404
rect 26608 7352 26660 7361
rect 27804 7361 27813 7395
rect 27813 7361 27847 7395
rect 27847 7361 27856 7395
rect 27804 7352 27856 7361
rect 26148 7327 26200 7336
rect 26148 7293 26157 7327
rect 26157 7293 26191 7327
rect 26191 7293 26200 7327
rect 26148 7284 26200 7293
rect 1676 7148 1728 7200
rect 27160 7191 27212 7200
rect 27160 7157 27169 7191
rect 27169 7157 27203 7191
rect 27203 7157 27212 7191
rect 27160 7148 27212 7157
rect 4423 7046 4475 7098
rect 4487 7046 4539 7098
rect 4551 7046 4603 7098
rect 4615 7046 4667 7098
rect 4679 7046 4731 7098
rect 11369 7046 11421 7098
rect 11433 7046 11485 7098
rect 11497 7046 11549 7098
rect 11561 7046 11613 7098
rect 11625 7046 11677 7098
rect 18315 7046 18367 7098
rect 18379 7046 18431 7098
rect 18443 7046 18495 7098
rect 18507 7046 18559 7098
rect 18571 7046 18623 7098
rect 25261 7046 25313 7098
rect 25325 7046 25377 7098
rect 25389 7046 25441 7098
rect 25453 7046 25505 7098
rect 25517 7046 25569 7098
rect 3976 6944 4028 6996
rect 5356 6944 5408 6996
rect 7748 6876 7800 6928
rect 1584 6783 1636 6792
rect 1584 6749 1593 6783
rect 1593 6749 1627 6783
rect 1627 6749 1636 6783
rect 1584 6740 1636 6749
rect 3976 6808 4028 6860
rect 4068 6808 4120 6860
rect 2872 6783 2924 6792
rect 2872 6749 2881 6783
rect 2881 6749 2915 6783
rect 2915 6749 2924 6783
rect 2872 6740 2924 6749
rect 2596 6672 2648 6724
rect 5356 6783 5408 6792
rect 5356 6749 5365 6783
rect 5365 6749 5399 6783
rect 5399 6749 5408 6783
rect 5356 6740 5408 6749
rect 5540 6740 5592 6792
rect 3056 6604 3108 6656
rect 4160 6604 4212 6656
rect 26424 6808 26476 6860
rect 27160 6808 27212 6860
rect 28356 6851 28408 6860
rect 28356 6817 28365 6851
rect 28365 6817 28399 6851
rect 28399 6817 28408 6851
rect 28356 6808 28408 6817
rect 25780 6740 25832 6792
rect 7896 6502 7948 6554
rect 7960 6502 8012 6554
rect 8024 6502 8076 6554
rect 8088 6502 8140 6554
rect 8152 6502 8204 6554
rect 14842 6502 14894 6554
rect 14906 6502 14958 6554
rect 14970 6502 15022 6554
rect 15034 6502 15086 6554
rect 15098 6502 15150 6554
rect 21788 6502 21840 6554
rect 21852 6502 21904 6554
rect 21916 6502 21968 6554
rect 21980 6502 22032 6554
rect 22044 6502 22096 6554
rect 28734 6502 28786 6554
rect 28798 6502 28850 6554
rect 28862 6502 28914 6554
rect 28926 6502 28978 6554
rect 28990 6502 29042 6554
rect 26700 6400 26752 6452
rect 4160 6375 4212 6384
rect 4160 6341 4169 6375
rect 4169 6341 4203 6375
rect 4203 6341 4212 6375
rect 4160 6332 4212 6341
rect 1676 6307 1728 6316
rect 1676 6273 1685 6307
rect 1685 6273 1719 6307
rect 1719 6273 1728 6307
rect 1676 6264 1728 6273
rect 26424 6264 26476 6316
rect 27988 6307 28040 6316
rect 27988 6273 27997 6307
rect 27997 6273 28031 6307
rect 28031 6273 28040 6307
rect 27988 6264 28040 6273
rect 1860 6239 1912 6248
rect 1860 6205 1869 6239
rect 1869 6205 1903 6239
rect 1903 6205 1912 6239
rect 1860 6196 1912 6205
rect 3148 6239 3200 6248
rect 3148 6205 3157 6239
rect 3157 6205 3191 6239
rect 3191 6205 3200 6239
rect 3148 6196 3200 6205
rect 3976 6239 4028 6248
rect 3976 6205 3985 6239
rect 3985 6205 4019 6239
rect 4019 6205 4028 6239
rect 3976 6196 4028 6205
rect 4344 6196 4396 6248
rect 28172 6060 28224 6112
rect 4423 5958 4475 6010
rect 4487 5958 4539 6010
rect 4551 5958 4603 6010
rect 4615 5958 4667 6010
rect 4679 5958 4731 6010
rect 11369 5958 11421 6010
rect 11433 5958 11485 6010
rect 11497 5958 11549 6010
rect 11561 5958 11613 6010
rect 11625 5958 11677 6010
rect 18315 5958 18367 6010
rect 18379 5958 18431 6010
rect 18443 5958 18495 6010
rect 18507 5958 18559 6010
rect 18571 5958 18623 6010
rect 25261 5958 25313 6010
rect 25325 5958 25377 6010
rect 25389 5958 25441 6010
rect 25453 5958 25505 6010
rect 25517 5958 25569 6010
rect 3976 5856 4028 5908
rect 1584 5763 1636 5772
rect 1584 5729 1593 5763
rect 1593 5729 1627 5763
rect 1627 5729 1636 5763
rect 1584 5720 1636 5729
rect 2780 5763 2832 5772
rect 2780 5729 2789 5763
rect 2789 5729 2823 5763
rect 2823 5729 2832 5763
rect 2780 5720 2832 5729
rect 27528 5763 27580 5772
rect 27528 5729 27537 5763
rect 27537 5729 27571 5763
rect 27571 5729 27580 5763
rect 27528 5720 27580 5729
rect 28172 5763 28224 5772
rect 28172 5729 28181 5763
rect 28181 5729 28215 5763
rect 28215 5729 28224 5763
rect 28172 5720 28224 5729
rect 28356 5695 28408 5704
rect 28356 5661 28365 5695
rect 28365 5661 28399 5695
rect 28399 5661 28408 5695
rect 28356 5652 28408 5661
rect 1768 5627 1820 5636
rect 1768 5593 1777 5627
rect 1777 5593 1811 5627
rect 1811 5593 1820 5627
rect 1768 5584 1820 5593
rect 7896 5414 7948 5466
rect 7960 5414 8012 5466
rect 8024 5414 8076 5466
rect 8088 5414 8140 5466
rect 8152 5414 8204 5466
rect 14842 5414 14894 5466
rect 14906 5414 14958 5466
rect 14970 5414 15022 5466
rect 15034 5414 15086 5466
rect 15098 5414 15150 5466
rect 21788 5414 21840 5466
rect 21852 5414 21904 5466
rect 21916 5414 21968 5466
rect 21980 5414 22032 5466
rect 22044 5414 22096 5466
rect 28734 5414 28786 5466
rect 28798 5414 28850 5466
rect 28862 5414 28914 5466
rect 28926 5414 28978 5466
rect 28990 5414 29042 5466
rect 1768 5312 1820 5364
rect 2504 5312 2556 5364
rect 3056 5287 3108 5296
rect 3056 5253 3065 5287
rect 3065 5253 3099 5287
rect 3099 5253 3108 5287
rect 3056 5244 3108 5253
rect 2044 5219 2096 5228
rect 2044 5185 2053 5219
rect 2053 5185 2087 5219
rect 2087 5185 2096 5219
rect 2044 5176 2096 5185
rect 2872 5219 2924 5228
rect 2872 5185 2881 5219
rect 2881 5185 2915 5219
rect 2915 5185 2924 5219
rect 2872 5176 2924 5185
rect 28356 5176 28408 5228
rect 4804 5108 4856 5160
rect 4252 4972 4304 5024
rect 12992 4972 13044 5024
rect 4423 4870 4475 4922
rect 4487 4870 4539 4922
rect 4551 4870 4603 4922
rect 4615 4870 4667 4922
rect 4679 4870 4731 4922
rect 11369 4870 11421 4922
rect 11433 4870 11485 4922
rect 11497 4870 11549 4922
rect 11561 4870 11613 4922
rect 11625 4870 11677 4922
rect 18315 4870 18367 4922
rect 18379 4870 18431 4922
rect 18443 4870 18495 4922
rect 18507 4870 18559 4922
rect 18571 4870 18623 4922
rect 25261 4870 25313 4922
rect 25325 4870 25377 4922
rect 25389 4870 25441 4922
rect 25453 4870 25505 4922
rect 25517 4870 25569 4922
rect 1860 4768 1912 4820
rect 2044 4607 2096 4616
rect 2044 4573 2053 4607
rect 2053 4573 2087 4607
rect 2087 4573 2096 4607
rect 2044 4564 2096 4573
rect 3148 4607 3200 4616
rect 3148 4573 3157 4607
rect 3157 4573 3191 4607
rect 3191 4573 3200 4607
rect 3148 4564 3200 4573
rect 3976 4607 4028 4616
rect 3976 4573 3985 4607
rect 3985 4573 4019 4607
rect 4019 4573 4028 4607
rect 3976 4564 4028 4573
rect 4988 4632 5040 4684
rect 5724 4632 5776 4684
rect 20628 4675 20680 4684
rect 20628 4641 20637 4675
rect 20637 4641 20671 4675
rect 20671 4641 20680 4675
rect 20628 4632 20680 4641
rect 21272 4675 21324 4684
rect 21272 4641 21281 4675
rect 21281 4641 21315 4675
rect 21315 4641 21324 4675
rect 21272 4632 21324 4641
rect 27528 4675 27580 4684
rect 27528 4641 27537 4675
rect 27537 4641 27571 4675
rect 27571 4641 27580 4675
rect 27528 4632 27580 4641
rect 4896 4564 4948 4616
rect 5540 4564 5592 4616
rect 12808 4564 12860 4616
rect 20444 4607 20496 4616
rect 20444 4573 20453 4607
rect 20453 4573 20487 4607
rect 20487 4573 20496 4607
rect 20444 4564 20496 4573
rect 25780 4607 25832 4616
rect 25780 4573 25789 4607
rect 25789 4573 25823 4607
rect 25823 4573 25832 4607
rect 25780 4564 25832 4573
rect 26516 4607 26568 4616
rect 26516 4573 26525 4607
rect 26525 4573 26559 4607
rect 26559 4573 26568 4607
rect 26516 4564 26568 4573
rect 16764 4496 16816 4548
rect 26700 4539 26752 4548
rect 26700 4505 26709 4539
rect 26709 4505 26743 4539
rect 26743 4505 26752 4539
rect 26700 4496 26752 4505
rect 4160 4428 4212 4480
rect 6736 4428 6788 4480
rect 25872 4471 25924 4480
rect 25872 4437 25881 4471
rect 25881 4437 25915 4471
rect 25915 4437 25924 4471
rect 25872 4428 25924 4437
rect 7896 4326 7948 4378
rect 7960 4326 8012 4378
rect 8024 4326 8076 4378
rect 8088 4326 8140 4378
rect 8152 4326 8204 4378
rect 14842 4326 14894 4378
rect 14906 4326 14958 4378
rect 14970 4326 15022 4378
rect 15034 4326 15086 4378
rect 15098 4326 15150 4378
rect 21788 4326 21840 4378
rect 21852 4326 21904 4378
rect 21916 4326 21968 4378
rect 21980 4326 22032 4378
rect 22044 4326 22096 4378
rect 28734 4326 28786 4378
rect 28798 4326 28850 4378
rect 28862 4326 28914 4378
rect 28926 4326 28978 4378
rect 28990 4326 29042 4378
rect 26700 4224 26752 4276
rect 4160 4199 4212 4208
rect 4160 4165 4169 4199
rect 4169 4165 4203 4199
rect 4203 4165 4212 4199
rect 4160 4156 4212 4165
rect 12992 4199 13044 4208
rect 12992 4165 13001 4199
rect 13001 4165 13035 4199
rect 13035 4165 13044 4199
rect 12992 4156 13044 4165
rect 3976 4131 4028 4140
rect 3976 4097 3985 4131
rect 3985 4097 4019 4131
rect 4019 4097 4028 4131
rect 3976 4088 4028 4097
rect 11980 4131 12032 4140
rect 11980 4097 11989 4131
rect 11989 4097 12023 4131
rect 12023 4097 12032 4131
rect 11980 4088 12032 4097
rect 12808 4131 12860 4140
rect 12808 4097 12817 4131
rect 12817 4097 12851 4131
rect 12851 4097 12860 4131
rect 12808 4088 12860 4097
rect 17132 4131 17184 4140
rect 17132 4097 17141 4131
rect 17141 4097 17175 4131
rect 17175 4097 17184 4131
rect 17132 4088 17184 4097
rect 20444 4088 20496 4140
rect 27620 4088 27672 4140
rect 664 4020 716 4072
rect 1860 4020 1912 4072
rect 4896 4020 4948 4072
rect 7748 4063 7800 4072
rect 3240 3952 3292 4004
rect 7748 4029 7757 4063
rect 7757 4029 7791 4063
rect 7791 4029 7800 4063
rect 7748 4020 7800 4029
rect 8392 4063 8444 4072
rect 7656 3952 7708 4004
rect 8392 4029 8401 4063
rect 8401 4029 8435 4063
rect 8435 4029 8444 4063
rect 8392 4020 8444 4029
rect 13544 4063 13596 4072
rect 13544 4029 13553 4063
rect 13553 4029 13587 4063
rect 13587 4029 13596 4063
rect 13544 4020 13596 4029
rect 16764 4020 16816 4072
rect 25780 4020 25832 4072
rect 26148 4063 26200 4072
rect 26148 4029 26157 4063
rect 26157 4029 26191 4063
rect 26191 4029 26200 4063
rect 26148 4020 26200 4029
rect 26424 4063 26476 4072
rect 26424 4029 26433 4063
rect 26433 4029 26467 4063
rect 26467 4029 26476 4063
rect 26424 4020 26476 4029
rect 14188 3952 14240 4004
rect 14556 3952 14608 4004
rect 18696 3952 18748 4004
rect 6552 3927 6604 3936
rect 6552 3893 6561 3927
rect 6561 3893 6595 3927
rect 6595 3893 6604 3927
rect 6552 3884 6604 3893
rect 12072 3927 12124 3936
rect 12072 3893 12081 3927
rect 12081 3893 12115 3927
rect 12115 3893 12124 3927
rect 12072 3884 12124 3893
rect 17224 3927 17276 3936
rect 17224 3893 17233 3927
rect 17233 3893 17267 3927
rect 17267 3893 17276 3927
rect 17224 3884 17276 3893
rect 4423 3782 4475 3834
rect 4487 3782 4539 3834
rect 4551 3782 4603 3834
rect 4615 3782 4667 3834
rect 4679 3782 4731 3834
rect 11369 3782 11421 3834
rect 11433 3782 11485 3834
rect 11497 3782 11549 3834
rect 11561 3782 11613 3834
rect 11625 3782 11677 3834
rect 18315 3782 18367 3834
rect 18379 3782 18431 3834
rect 18443 3782 18495 3834
rect 18507 3782 18559 3834
rect 18571 3782 18623 3834
rect 25261 3782 25313 3834
rect 25325 3782 25377 3834
rect 25389 3782 25441 3834
rect 25453 3782 25505 3834
rect 25517 3782 25569 3834
rect 7748 3680 7800 3732
rect 18052 3723 18104 3732
rect 18052 3689 18061 3723
rect 18061 3689 18095 3723
rect 18095 3689 18104 3723
rect 18052 3680 18104 3689
rect 3148 3544 3200 3596
rect 5816 3587 5868 3596
rect 5816 3553 5825 3587
rect 5825 3553 5859 3587
rect 5859 3553 5868 3587
rect 5816 3544 5868 3553
rect 11888 3587 11940 3596
rect 11888 3553 11897 3587
rect 11897 3553 11931 3587
rect 11931 3553 11940 3587
rect 11888 3544 11940 3553
rect 12072 3587 12124 3596
rect 12072 3553 12081 3587
rect 12081 3553 12115 3587
rect 12115 3553 12124 3587
rect 12072 3544 12124 3553
rect 12440 3587 12492 3596
rect 12440 3553 12449 3587
rect 12449 3553 12483 3587
rect 12483 3553 12492 3587
rect 25688 3680 25740 3732
rect 26424 3680 26476 3732
rect 18696 3612 18748 3664
rect 12440 3544 12492 3553
rect 8944 3476 8996 3528
rect 9956 3519 10008 3528
rect 9956 3485 9965 3519
rect 9965 3485 9999 3519
rect 9999 3485 10008 3519
rect 9956 3476 10008 3485
rect 10600 3519 10652 3528
rect 10600 3485 10609 3519
rect 10609 3485 10643 3519
rect 10643 3485 10652 3519
rect 10600 3476 10652 3485
rect 1584 3451 1636 3460
rect 1584 3417 1593 3451
rect 1593 3417 1627 3451
rect 1627 3417 1636 3451
rect 1584 3408 1636 3417
rect 2504 3408 2556 3460
rect 5264 3451 5316 3460
rect 5264 3417 5273 3451
rect 5273 3417 5307 3451
rect 5307 3417 5316 3451
rect 5264 3408 5316 3417
rect 11704 3476 11756 3528
rect 14280 3476 14332 3528
rect 16304 3519 16356 3528
rect 16304 3485 16313 3519
rect 16313 3485 16347 3519
rect 16347 3485 16356 3519
rect 16304 3476 16356 3485
rect 16764 3519 16816 3528
rect 16764 3485 16773 3519
rect 16773 3485 16807 3519
rect 16807 3485 16816 3519
rect 16764 3476 16816 3485
rect 17408 3519 17460 3528
rect 17408 3485 17417 3519
rect 17417 3485 17451 3519
rect 17451 3485 17460 3519
rect 17408 3476 17460 3485
rect 17500 3476 17552 3528
rect 9128 3340 9180 3392
rect 11888 3340 11940 3392
rect 17040 3340 17092 3392
rect 17132 3340 17184 3392
rect 19248 3476 19300 3528
rect 21548 3519 21600 3528
rect 21548 3485 21557 3519
rect 21557 3485 21591 3519
rect 21591 3485 21600 3519
rect 21548 3476 21600 3485
rect 25872 3587 25924 3596
rect 25872 3553 25881 3587
rect 25881 3553 25915 3587
rect 25915 3553 25924 3587
rect 25872 3544 25924 3553
rect 23848 3519 23900 3528
rect 23848 3485 23857 3519
rect 23857 3485 23891 3519
rect 23891 3485 23900 3519
rect 23848 3476 23900 3485
rect 24308 3476 24360 3528
rect 27620 3476 27672 3528
rect 27896 3476 27948 3528
rect 27436 3408 27488 3460
rect 19432 3340 19484 3392
rect 22192 3340 22244 3392
rect 24492 3340 24544 3392
rect 7896 3238 7948 3290
rect 7960 3238 8012 3290
rect 8024 3238 8076 3290
rect 8088 3238 8140 3290
rect 8152 3238 8204 3290
rect 14842 3238 14894 3290
rect 14906 3238 14958 3290
rect 14970 3238 15022 3290
rect 15034 3238 15086 3290
rect 15098 3238 15150 3290
rect 21788 3238 21840 3290
rect 21852 3238 21904 3290
rect 21916 3238 21968 3290
rect 21980 3238 22032 3290
rect 22044 3238 22096 3290
rect 28734 3238 28786 3290
rect 28798 3238 28850 3290
rect 28862 3238 28914 3290
rect 28926 3238 28978 3290
rect 28990 3238 29042 3290
rect 1860 3179 1912 3188
rect 1860 3145 1869 3179
rect 1869 3145 1903 3179
rect 1903 3145 1912 3179
rect 1860 3136 1912 3145
rect 2504 3179 2556 3188
rect 2504 3145 2513 3179
rect 2513 3145 2547 3179
rect 2547 3145 2556 3179
rect 2504 3136 2556 3145
rect 9956 3136 10008 3188
rect 14188 3136 14240 3188
rect 17132 3136 17184 3188
rect 9128 3111 9180 3120
rect 9128 3077 9137 3111
rect 9137 3077 9171 3111
rect 9171 3077 9180 3111
rect 9128 3068 9180 3077
rect 11888 3111 11940 3120
rect 11888 3077 11897 3111
rect 11897 3077 11931 3111
rect 11931 3077 11940 3111
rect 11888 3068 11940 3077
rect 17040 3111 17092 3120
rect 17040 3077 17049 3111
rect 17049 3077 17083 3111
rect 17083 3077 17092 3111
rect 17040 3068 17092 3077
rect 19432 3111 19484 3120
rect 19432 3077 19441 3111
rect 19441 3077 19475 3111
rect 19475 3077 19484 3111
rect 19432 3068 19484 3077
rect 22192 3111 22244 3120
rect 22192 3077 22201 3111
rect 22201 3077 22235 3111
rect 22235 3077 22244 3111
rect 22192 3068 22244 3077
rect 24492 3111 24544 3120
rect 24492 3077 24501 3111
rect 24501 3077 24535 3111
rect 24535 3077 24544 3111
rect 24492 3068 24544 3077
rect 6552 3043 6604 3052
rect 6552 3009 6561 3043
rect 6561 3009 6595 3043
rect 6595 3009 6604 3043
rect 6552 3000 6604 3009
rect 8944 3043 8996 3052
rect 8944 3009 8953 3043
rect 8953 3009 8987 3043
rect 8987 3009 8996 3043
rect 8944 3000 8996 3009
rect 11704 3043 11756 3052
rect 11704 3009 11713 3043
rect 11713 3009 11747 3043
rect 11747 3009 11756 3043
rect 11704 3000 11756 3009
rect 14280 3043 14332 3052
rect 14280 3009 14289 3043
rect 14289 3009 14323 3043
rect 14323 3009 14332 3043
rect 14280 3000 14332 3009
rect 16304 3000 16356 3052
rect 19248 3043 19300 3052
rect 19248 3009 19257 3043
rect 19257 3009 19291 3043
rect 19291 3009 19300 3043
rect 19248 3000 19300 3009
rect 21548 3000 21600 3052
rect 24308 3043 24360 3052
rect 24308 3009 24317 3043
rect 24317 3009 24351 3043
rect 24351 3009 24360 3043
rect 24308 3000 24360 3009
rect 26516 3000 26568 3052
rect 27896 3000 27948 3052
rect 3884 2975 3936 2984
rect 3884 2941 3893 2975
rect 3893 2941 3927 2975
rect 3927 2941 3936 2975
rect 3884 2932 3936 2941
rect 3976 2932 4028 2984
rect 6736 2975 6788 2984
rect 6736 2941 6745 2975
rect 6745 2941 6779 2975
rect 6779 2941 6788 2975
rect 6736 2932 6788 2941
rect 6460 2864 6512 2916
rect 9680 2975 9732 2984
rect 9680 2941 9689 2975
rect 9689 2941 9723 2975
rect 9723 2941 9732 2975
rect 9680 2932 9732 2941
rect 10968 2932 11020 2984
rect 14464 2975 14516 2984
rect 14464 2941 14473 2975
rect 14473 2941 14507 2975
rect 14507 2941 14516 2975
rect 14464 2932 14516 2941
rect 14740 2975 14792 2984
rect 14740 2941 14749 2975
rect 14749 2941 14783 2975
rect 14783 2941 14792 2975
rect 14740 2932 14792 2941
rect 16764 2932 16816 2984
rect 19984 2975 20036 2984
rect 19984 2941 19993 2975
rect 19993 2941 20027 2975
rect 20027 2941 20036 2975
rect 19984 2932 20036 2941
rect 21640 2864 21692 2916
rect 25136 2975 25188 2984
rect 25136 2941 25145 2975
rect 25145 2941 25179 2975
rect 25179 2941 25188 2975
rect 25136 2932 25188 2941
rect 2596 2796 2648 2848
rect 4804 2796 4856 2848
rect 26424 2796 26476 2848
rect 4423 2694 4475 2746
rect 4487 2694 4539 2746
rect 4551 2694 4603 2746
rect 4615 2694 4667 2746
rect 4679 2694 4731 2746
rect 11369 2694 11421 2746
rect 11433 2694 11485 2746
rect 11497 2694 11549 2746
rect 11561 2694 11613 2746
rect 11625 2694 11677 2746
rect 18315 2694 18367 2746
rect 18379 2694 18431 2746
rect 18443 2694 18495 2746
rect 18507 2694 18559 2746
rect 18571 2694 18623 2746
rect 25261 2694 25313 2746
rect 25325 2694 25377 2746
rect 25389 2694 25441 2746
rect 25453 2694 25505 2746
rect 25517 2694 25569 2746
rect 3884 2592 3936 2644
rect 5264 2635 5316 2644
rect 5264 2601 5273 2635
rect 5273 2601 5307 2635
rect 5307 2601 5316 2635
rect 5264 2592 5316 2601
rect 7656 2592 7708 2644
rect 14464 2592 14516 2644
rect 16856 2592 16908 2644
rect 2320 2524 2372 2576
rect 23848 2592 23900 2644
rect 27068 2592 27120 2644
rect 2780 2499 2832 2508
rect 2780 2465 2789 2499
rect 2789 2465 2823 2499
rect 2823 2465 2832 2499
rect 2780 2456 2832 2465
rect 3792 2456 3844 2508
rect 4160 2431 4212 2440
rect 4160 2397 4169 2431
rect 4169 2397 4203 2431
rect 4203 2397 4212 2431
rect 4160 2388 4212 2397
rect 9404 2499 9456 2508
rect 9404 2465 9413 2499
rect 9413 2465 9447 2499
rect 9447 2465 9456 2499
rect 9404 2456 9456 2465
rect 17408 2524 17460 2576
rect 17224 2499 17276 2508
rect 17224 2465 17233 2499
rect 17233 2465 17267 2499
rect 17267 2465 17276 2499
rect 17224 2456 17276 2465
rect 18052 2499 18104 2508
rect 18052 2465 18061 2499
rect 18061 2465 18095 2499
rect 18095 2465 18104 2499
rect 18052 2456 18104 2465
rect 26148 2499 26200 2508
rect 26148 2465 26157 2499
rect 26157 2465 26191 2499
rect 26191 2465 26200 2499
rect 26148 2456 26200 2465
rect 26424 2499 26476 2508
rect 26424 2465 26433 2499
rect 26433 2465 26467 2499
rect 26467 2465 26476 2499
rect 26424 2456 26476 2465
rect 5724 2388 5776 2440
rect 9036 2388 9088 2440
rect 14188 2388 14240 2440
rect 27068 2388 27120 2440
rect 16120 2363 16172 2372
rect 16120 2329 16129 2363
rect 16129 2329 16163 2363
rect 16163 2329 16172 2363
rect 16120 2320 16172 2329
rect 4068 2252 4120 2304
rect 12440 2252 12492 2304
rect 7896 2150 7948 2202
rect 7960 2150 8012 2202
rect 8024 2150 8076 2202
rect 8088 2150 8140 2202
rect 8152 2150 8204 2202
rect 14842 2150 14894 2202
rect 14906 2150 14958 2202
rect 14970 2150 15022 2202
rect 15034 2150 15086 2202
rect 15098 2150 15150 2202
rect 21788 2150 21840 2202
rect 21852 2150 21904 2202
rect 21916 2150 21968 2202
rect 21980 2150 22032 2202
rect 22044 2150 22096 2202
rect 28734 2150 28786 2202
rect 28798 2150 28850 2202
rect 28862 2150 28914 2202
rect 28926 2150 28978 2202
rect 28990 2150 29042 2202
rect 4160 2048 4212 2100
rect 10600 2048 10652 2100
<< metal2 >>
rect -10 49200 102 49800
rect 634 49200 746 49800
rect 1278 49314 1390 49800
rect 952 49286 1390 49314
rect 20 47456 72 47462
rect 20 47398 72 47404
rect 32 43382 60 47398
rect 676 45554 704 49200
rect 952 47462 980 49286
rect 1278 49200 1390 49286
rect 1922 49200 2034 49800
rect 2566 49200 2678 49800
rect 2962 49736 3018 49745
rect 2962 49671 3018 49680
rect 940 47456 992 47462
rect 940 47398 992 47404
rect 1964 47122 1992 49200
rect 1952 47116 2004 47122
rect 1952 47058 2004 47064
rect 2608 46442 2636 49200
rect 2596 46436 2648 46442
rect 2596 46378 2648 46384
rect 1584 46368 1636 46374
rect 1584 46310 1636 46316
rect 1596 46034 1624 46310
rect 2976 46034 3004 49671
rect 3210 49200 3322 49800
rect 4498 49200 4610 49800
rect 5142 49200 5254 49800
rect 5786 49200 5898 49800
rect 6430 49200 6542 49800
rect 7074 49200 7186 49800
rect 7718 49200 7830 49800
rect 8362 49200 8474 49800
rect 9650 49200 9762 49800
rect 10294 49200 10406 49800
rect 10938 49200 11050 49800
rect 11582 49200 11694 49800
rect 12226 49200 12338 49800
rect 12870 49200 12982 49800
rect 13514 49200 13626 49800
rect 14802 49200 14914 49800
rect 15446 49200 15558 49800
rect 16090 49200 16202 49800
rect 16734 49200 16846 49800
rect 17378 49200 17490 49800
rect 18022 49200 18134 49800
rect 18666 49200 18778 49800
rect 19954 49200 20066 49800
rect 20598 49200 20710 49800
rect 21242 49200 21354 49800
rect 21886 49200 21998 49800
rect 22530 49200 22642 49800
rect 23174 49200 23286 49800
rect 23818 49200 23930 49800
rect 25106 49200 25218 49800
rect 25750 49200 25862 49800
rect 26394 49200 26506 49800
rect 27038 49200 27150 49800
rect 27682 49200 27794 49800
rect 28326 49200 28438 49800
rect 28970 49200 29082 49800
rect 29614 49200 29726 49800
rect 4423 47356 4731 47365
rect 4423 47354 4429 47356
rect 4485 47354 4509 47356
rect 4565 47354 4589 47356
rect 4645 47354 4669 47356
rect 4725 47354 4731 47356
rect 4485 47302 4487 47354
rect 4667 47302 4669 47354
rect 4423 47300 4429 47302
rect 4485 47300 4509 47302
rect 4565 47300 4589 47302
rect 4645 47300 4669 47302
rect 4725 47300 4731 47302
rect 4423 47291 4731 47300
rect 5828 47054 5856 49200
rect 6472 47054 6500 49200
rect 3516 47048 3568 47054
rect 3516 46990 3568 46996
rect 5816 47048 5868 47054
rect 5816 46990 5868 46996
rect 6460 47048 6512 47054
rect 6460 46990 6512 46996
rect 7012 47048 7064 47054
rect 7012 46990 7064 46996
rect 3240 46980 3292 46986
rect 3240 46922 3292 46928
rect 1584 46028 1636 46034
rect 1584 45970 1636 45976
rect 2964 46028 3016 46034
rect 2964 45970 3016 45976
rect 1952 45892 2004 45898
rect 1952 45834 2004 45840
rect 1964 45626 1992 45834
rect 1952 45620 2004 45626
rect 1952 45562 2004 45568
rect 3252 45558 3280 46922
rect 124 45526 704 45554
rect 2412 45552 2464 45558
rect 124 43858 152 45526
rect 3240 45552 3292 45558
rect 2464 45500 2544 45506
rect 2412 45494 2544 45500
rect 3240 45494 3292 45500
rect 2424 45478 2544 45494
rect 3528 45490 3556 46990
rect 6000 46912 6052 46918
rect 6000 46854 6052 46860
rect 6736 46912 6788 46918
rect 6736 46854 6788 46860
rect 4068 46504 4120 46510
rect 4068 46446 4120 46452
rect 4080 46170 4108 46446
rect 4423 46268 4731 46277
rect 4423 46266 4429 46268
rect 4485 46266 4509 46268
rect 4565 46266 4589 46268
rect 4645 46266 4669 46268
rect 4725 46266 4731 46268
rect 4485 46214 4487 46266
rect 4667 46214 4669 46266
rect 4423 46212 4429 46214
rect 4485 46212 4509 46214
rect 4565 46212 4589 46214
rect 4645 46212 4669 46214
rect 4725 46212 4731 46214
rect 4423 46203 4731 46212
rect 4068 46164 4120 46170
rect 4068 46106 4120 46112
rect 4804 45960 4856 45966
rect 4804 45902 4856 45908
rect 2320 45416 2372 45422
rect 2320 45358 2372 45364
rect 112 43852 164 43858
rect 112 43794 164 43800
rect 20 43376 72 43382
rect 20 43318 72 43324
rect 1582 42256 1638 42265
rect 1582 42191 1638 42200
rect 1596 41682 1624 42191
rect 1676 42016 1728 42022
rect 1676 41958 1728 41964
rect 1584 41676 1636 41682
rect 1584 41618 1636 41624
rect 1688 41138 1716 41958
rect 1676 41132 1728 41138
rect 1676 41074 1728 41080
rect 2228 41064 2280 41070
rect 2228 41006 2280 41012
rect 2240 40730 2268 41006
rect 2228 40724 2280 40730
rect 2228 40666 2280 40672
rect 2332 40526 2360 45358
rect 2412 44396 2464 44402
rect 2412 44338 2464 44344
rect 2424 42702 2452 44338
rect 2412 42696 2464 42702
rect 2412 42638 2464 42644
rect 2320 40520 2372 40526
rect 2320 40462 2372 40468
rect 1676 39840 1728 39846
rect 1676 39782 1728 39788
rect 1584 38752 1636 38758
rect 1584 38694 1636 38700
rect 1492 37256 1544 37262
rect 1492 37198 1544 37204
rect 1504 11150 1532 37198
rect 1596 35086 1624 38694
rect 1688 38486 1716 39782
rect 1768 39296 1820 39302
rect 1768 39238 1820 39244
rect 1676 38480 1728 38486
rect 1676 38422 1728 38428
rect 1780 38418 1808 39238
rect 1768 38412 1820 38418
rect 1768 38354 1820 38360
rect 1676 37800 1728 37806
rect 1676 37742 1728 37748
rect 1688 37505 1716 37742
rect 1674 37496 1730 37505
rect 1674 37431 1730 37440
rect 2424 36718 2452 42638
rect 2516 42226 2544 45478
rect 3516 45484 3568 45490
rect 3516 45426 3568 45432
rect 4423 45180 4731 45189
rect 4423 45178 4429 45180
rect 4485 45178 4509 45180
rect 4565 45178 4589 45180
rect 4645 45178 4669 45180
rect 4725 45178 4731 45180
rect 4485 45126 4487 45178
rect 4667 45126 4669 45178
rect 4423 45124 4429 45126
rect 4485 45124 4509 45126
rect 4565 45124 4589 45126
rect 4645 45124 4669 45126
rect 4725 45124 4731 45126
rect 4423 45115 4731 45124
rect 4816 45014 4844 45902
rect 4804 45008 4856 45014
rect 4250 44976 4306 44985
rect 4804 44950 4856 44956
rect 4250 44911 4306 44920
rect 3056 44872 3108 44878
rect 3056 44814 3108 44820
rect 3148 44872 3200 44878
rect 3148 44814 3200 44820
rect 3068 43858 3096 44814
rect 3160 44402 3188 44814
rect 3148 44396 3200 44402
rect 3148 44338 3200 44344
rect 3332 44328 3384 44334
rect 3608 44328 3660 44334
rect 3332 44270 3384 44276
rect 3606 44296 3608 44305
rect 3660 44296 3662 44305
rect 3344 43994 3372 44270
rect 3606 44231 3662 44240
rect 3608 44192 3660 44198
rect 3608 44134 3660 44140
rect 3332 43988 3384 43994
rect 3332 43930 3384 43936
rect 3056 43852 3108 43858
rect 3056 43794 3108 43800
rect 3240 43716 3292 43722
rect 3240 43658 3292 43664
rect 3252 42770 3280 43658
rect 3620 43382 3648 44134
rect 4160 43784 4212 43790
rect 4160 43726 4212 43732
rect 3608 43376 3660 43382
rect 3608 43318 3660 43324
rect 3240 42764 3292 42770
rect 3240 42706 3292 42712
rect 3424 42628 3476 42634
rect 3424 42570 3476 42576
rect 2504 42220 2556 42226
rect 2504 42162 2556 42168
rect 2136 36712 2188 36718
rect 2136 36654 2188 36660
rect 2412 36712 2464 36718
rect 2412 36654 2464 36660
rect 1674 36136 1730 36145
rect 1674 36071 1730 36080
rect 1688 35766 1716 36071
rect 1676 35760 1728 35766
rect 1676 35702 1728 35708
rect 1584 35080 1636 35086
rect 1584 35022 1636 35028
rect 1676 34536 1728 34542
rect 1676 34478 1728 34484
rect 1860 34536 1912 34542
rect 1860 34478 1912 34484
rect 1688 33522 1716 34478
rect 1872 34202 1900 34478
rect 1860 34196 1912 34202
rect 1860 34138 1912 34144
rect 1676 33516 1728 33522
rect 1676 33458 1728 33464
rect 1676 32904 1728 32910
rect 1676 32846 1728 32852
rect 1688 32434 1716 32846
rect 1676 32428 1728 32434
rect 1676 32370 1728 32376
rect 2044 32360 2096 32366
rect 2044 32302 2096 32308
rect 2056 32026 2084 32302
rect 2044 32020 2096 32026
rect 2044 31962 2096 31968
rect 2148 30870 2176 36654
rect 2412 36168 2464 36174
rect 2412 36110 2464 36116
rect 2424 35154 2452 36110
rect 2412 35148 2464 35154
rect 2412 35090 2464 35096
rect 2320 33992 2372 33998
rect 2320 33934 2372 33940
rect 2136 30864 2188 30870
rect 2136 30806 2188 30812
rect 1584 30252 1636 30258
rect 1584 30194 1636 30200
rect 1596 30025 1624 30194
rect 1860 30048 1912 30054
rect 1582 30016 1638 30025
rect 1860 29990 1912 29996
rect 1582 29951 1638 29960
rect 1584 28076 1636 28082
rect 1584 28018 1636 28024
rect 1596 27985 1624 28018
rect 1582 27976 1638 27985
rect 1582 27911 1638 27920
rect 1768 27872 1820 27878
rect 1768 27814 1820 27820
rect 1780 27402 1808 27814
rect 1768 27396 1820 27402
rect 1768 27338 1820 27344
rect 1676 26376 1728 26382
rect 1676 26318 1728 26324
rect 1688 25906 1716 26318
rect 1676 25900 1728 25906
rect 1676 25842 1728 25848
rect 1584 25288 1636 25294
rect 1582 25256 1584 25265
rect 1636 25256 1638 25265
rect 1582 25191 1638 25200
rect 1768 25152 1820 25158
rect 1768 25094 1820 25100
rect 1780 24954 1808 25094
rect 1768 24948 1820 24954
rect 1768 24890 1820 24896
rect 1872 22574 1900 29990
rect 2148 26234 2176 30806
rect 2056 26206 2176 26234
rect 1860 22568 1912 22574
rect 1860 22510 1912 22516
rect 1584 20256 1636 20262
rect 1584 20198 1636 20204
rect 1768 20256 1820 20262
rect 1768 20198 1820 20204
rect 1596 19922 1624 20198
rect 1780 19922 1808 20198
rect 1584 19916 1636 19922
rect 1584 19858 1636 19864
rect 1768 19916 1820 19922
rect 1768 19858 1820 19864
rect 1676 19304 1728 19310
rect 1676 19246 1728 19252
rect 1860 19304 1912 19310
rect 1860 19246 1912 19252
rect 1688 18970 1716 19246
rect 1872 18970 1900 19246
rect 1676 18964 1728 18970
rect 1676 18906 1728 18912
rect 1860 18964 1912 18970
rect 1860 18906 1912 18912
rect 1582 18456 1638 18465
rect 1582 18391 1638 18400
rect 1596 18290 1624 18391
rect 1584 18284 1636 18290
rect 1584 18226 1636 18232
rect 1584 17672 1636 17678
rect 1584 17614 1636 17620
rect 1596 17202 1624 17614
rect 1584 17196 1636 17202
rect 1584 17138 1636 17144
rect 1676 16584 1728 16590
rect 1676 16526 1728 16532
rect 1688 16114 1716 16526
rect 1676 16108 1728 16114
rect 1676 16050 1728 16056
rect 1582 14376 1638 14385
rect 1582 14311 1584 14320
rect 1636 14311 1638 14320
rect 1584 14282 1636 14288
rect 1582 13696 1638 13705
rect 1582 13631 1638 13640
rect 1596 13394 1624 13631
rect 1584 13388 1636 13394
rect 1584 13330 1636 13336
rect 1952 13252 2004 13258
rect 1952 13194 2004 13200
rect 1964 12986 1992 13194
rect 1952 12980 2004 12986
rect 1952 12922 2004 12928
rect 2056 12850 2084 26206
rect 2136 19304 2188 19310
rect 2136 19246 2188 19252
rect 2148 19145 2176 19246
rect 2134 19136 2190 19145
rect 2134 19071 2190 19080
rect 2228 16040 2280 16046
rect 2228 15982 2280 15988
rect 2240 15706 2268 15982
rect 2228 15700 2280 15706
rect 2228 15642 2280 15648
rect 2332 15502 2360 33934
rect 2412 25832 2464 25838
rect 2412 25774 2464 25780
rect 2424 25498 2452 25774
rect 2412 25492 2464 25498
rect 2412 25434 2464 25440
rect 2516 20466 2544 42162
rect 3240 42016 3292 42022
rect 3240 41958 3292 41964
rect 3252 41682 3280 41958
rect 3436 41682 3464 42570
rect 3240 41676 3292 41682
rect 3240 41618 3292 41624
rect 3424 41676 3476 41682
rect 3424 41618 3476 41624
rect 2778 41576 2834 41585
rect 2778 41511 2834 41520
rect 2792 41070 2820 41511
rect 2780 41064 2832 41070
rect 2780 41006 2832 41012
rect 2780 39432 2832 39438
rect 2780 39374 2832 39380
rect 3240 39432 3292 39438
rect 3240 39374 3292 39380
rect 2792 38962 2820 39374
rect 2964 39296 3016 39302
rect 2964 39238 3016 39244
rect 2976 39030 3004 39238
rect 2964 39024 3016 39030
rect 2964 38966 3016 38972
rect 2780 38956 2832 38962
rect 2780 38898 2832 38904
rect 2778 38856 2834 38865
rect 2778 38791 2834 38800
rect 2872 38820 2924 38826
rect 2792 38418 2820 38791
rect 2872 38762 2924 38768
rect 2780 38412 2832 38418
rect 2780 38354 2832 38360
rect 2780 37800 2832 37806
rect 2780 37742 2832 37748
rect 2792 37262 2820 37742
rect 2780 37256 2832 37262
rect 2780 37198 2832 37204
rect 2688 37188 2740 37194
rect 2688 37130 2740 37136
rect 2700 37074 2728 37130
rect 2608 37046 2728 37074
rect 2608 36786 2636 37046
rect 2884 36825 2912 38762
rect 2870 36816 2926 36825
rect 2596 36780 2648 36786
rect 2870 36751 2926 36760
rect 2596 36722 2648 36728
rect 2608 36174 2636 36722
rect 2596 36168 2648 36174
rect 2596 36110 2648 36116
rect 3252 36106 3280 39374
rect 4172 36718 4200 43726
rect 4264 38894 4292 44911
rect 4423 44092 4731 44101
rect 4423 44090 4429 44092
rect 4485 44090 4509 44092
rect 4565 44090 4589 44092
rect 4645 44090 4669 44092
rect 4725 44090 4731 44092
rect 4485 44038 4487 44090
rect 4667 44038 4669 44090
rect 4423 44036 4429 44038
rect 4485 44036 4509 44038
rect 4565 44036 4589 44038
rect 4645 44036 4669 44038
rect 4725 44036 4731 44038
rect 4423 44027 4731 44036
rect 4620 43784 4672 43790
rect 4620 43726 4672 43732
rect 4632 43314 4660 43726
rect 4620 43308 4672 43314
rect 4620 43250 4672 43256
rect 4423 43004 4731 43013
rect 4423 43002 4429 43004
rect 4485 43002 4509 43004
rect 4565 43002 4589 43004
rect 4645 43002 4669 43004
rect 4725 43002 4731 43004
rect 4485 42950 4487 43002
rect 4667 42950 4669 43002
rect 4423 42948 4429 42950
rect 4485 42948 4509 42950
rect 4565 42948 4589 42950
rect 4645 42948 4669 42950
rect 4725 42948 4731 42950
rect 4423 42939 4731 42948
rect 4423 41916 4731 41925
rect 4423 41914 4429 41916
rect 4485 41914 4509 41916
rect 4565 41914 4589 41916
rect 4645 41914 4669 41916
rect 4725 41914 4731 41916
rect 4485 41862 4487 41914
rect 4667 41862 4669 41914
rect 4423 41860 4429 41862
rect 4485 41860 4509 41862
rect 4565 41860 4589 41862
rect 4645 41860 4669 41862
rect 4725 41860 4731 41862
rect 4423 41851 4731 41860
rect 4423 40828 4731 40837
rect 4423 40826 4429 40828
rect 4485 40826 4509 40828
rect 4565 40826 4589 40828
rect 4645 40826 4669 40828
rect 4725 40826 4731 40828
rect 4485 40774 4487 40826
rect 4667 40774 4669 40826
rect 4423 40772 4429 40774
rect 4485 40772 4509 40774
rect 4565 40772 4589 40774
rect 4645 40772 4669 40774
rect 4725 40772 4731 40774
rect 4423 40763 4731 40772
rect 4423 39740 4731 39749
rect 4423 39738 4429 39740
rect 4485 39738 4509 39740
rect 4565 39738 4589 39740
rect 4645 39738 4669 39740
rect 4725 39738 4731 39740
rect 4485 39686 4487 39738
rect 4667 39686 4669 39738
rect 4423 39684 4429 39686
rect 4485 39684 4509 39686
rect 4565 39684 4589 39686
rect 4645 39684 4669 39686
rect 4725 39684 4731 39686
rect 4423 39675 4731 39684
rect 4344 39364 4396 39370
rect 4344 39306 4396 39312
rect 4252 38888 4304 38894
rect 4252 38830 4304 38836
rect 4356 37194 4384 39306
rect 4423 38652 4731 38661
rect 4423 38650 4429 38652
rect 4485 38650 4509 38652
rect 4565 38650 4589 38652
rect 4645 38650 4669 38652
rect 4725 38650 4731 38652
rect 4485 38598 4487 38650
rect 4667 38598 4669 38650
rect 4423 38596 4429 38598
rect 4485 38596 4509 38598
rect 4565 38596 4589 38598
rect 4645 38596 4669 38598
rect 4725 38596 4731 38598
rect 4423 38587 4731 38596
rect 4423 37564 4731 37573
rect 4423 37562 4429 37564
rect 4485 37562 4509 37564
rect 4565 37562 4589 37564
rect 4645 37562 4669 37564
rect 4725 37562 4731 37564
rect 4485 37510 4487 37562
rect 4667 37510 4669 37562
rect 4423 37508 4429 37510
rect 4485 37508 4509 37510
rect 4565 37508 4589 37510
rect 4645 37508 4669 37510
rect 4725 37508 4731 37510
rect 4423 37499 4731 37508
rect 4344 37188 4396 37194
rect 4344 37130 4396 37136
rect 4356 36854 4384 37130
rect 4344 36848 4396 36854
rect 4344 36790 4396 36796
rect 4160 36712 4212 36718
rect 4160 36654 4212 36660
rect 4356 36530 4384 36790
rect 4172 36502 4384 36530
rect 3516 36236 3568 36242
rect 3516 36178 3568 36184
rect 2964 36100 3016 36106
rect 2964 36042 3016 36048
rect 3240 36100 3292 36106
rect 3240 36042 3292 36048
rect 2778 34776 2834 34785
rect 2778 34711 2834 34720
rect 2792 34542 2820 34711
rect 2780 34536 2832 34542
rect 2780 34478 2832 34484
rect 2780 32360 2832 32366
rect 2780 32302 2832 32308
rect 2792 32065 2820 32302
rect 2778 32056 2834 32065
rect 2778 31991 2834 32000
rect 2596 31816 2648 31822
rect 2596 31758 2648 31764
rect 2504 20460 2556 20466
rect 2504 20402 2556 20408
rect 2412 17604 2464 17610
rect 2412 17546 2464 17552
rect 2424 17338 2452 17546
rect 2412 17332 2464 17338
rect 2412 17274 2464 17280
rect 2516 17202 2544 20402
rect 2608 18766 2636 31758
rect 2778 25936 2834 25945
rect 2778 25871 2834 25880
rect 2792 25838 2820 25871
rect 2780 25832 2832 25838
rect 2780 25774 2832 25780
rect 2780 19916 2832 19922
rect 2780 19858 2832 19864
rect 2792 19825 2820 19858
rect 2778 19816 2834 19825
rect 2778 19751 2834 19760
rect 2596 18760 2648 18766
rect 2596 18702 2648 18708
rect 2504 17196 2556 17202
rect 2504 17138 2556 17144
rect 2320 15496 2372 15502
rect 2320 15438 2372 15444
rect 2044 12844 2096 12850
rect 2044 12786 2096 12792
rect 1676 12232 1728 12238
rect 1676 12174 1728 12180
rect 1688 11762 1716 12174
rect 1676 11756 1728 11762
rect 1676 11698 1728 11704
rect 1860 11688 1912 11694
rect 1860 11630 1912 11636
rect 1872 11354 1900 11630
rect 1860 11348 1912 11354
rect 1860 11290 1912 11296
rect 1492 11144 1544 11150
rect 1492 11086 1544 11092
rect 1504 7886 1532 11086
rect 1676 10056 1728 10062
rect 1676 9998 1728 10004
rect 1688 9586 1716 9998
rect 1676 9580 1728 9586
rect 1676 9522 1728 9528
rect 1860 9512 1912 9518
rect 1860 9454 1912 9460
rect 1584 8968 1636 8974
rect 1584 8910 1636 8916
rect 1596 8090 1624 8910
rect 1768 8900 1820 8906
rect 1768 8842 1820 8848
rect 1780 8090 1808 8842
rect 1872 8634 1900 9454
rect 1860 8628 1912 8634
rect 1860 8570 1912 8576
rect 1584 8084 1636 8090
rect 1584 8026 1636 8032
rect 1768 8084 1820 8090
rect 1768 8026 1820 8032
rect 1492 7880 1544 7886
rect 1492 7822 1544 7828
rect 1676 7200 1728 7206
rect 1676 7142 1728 7148
rect 1584 6792 1636 6798
rect 1584 6734 1636 6740
rect 1596 5778 1624 6734
rect 1688 6322 1716 7142
rect 1676 6316 1728 6322
rect 1676 6258 1728 6264
rect 1860 6248 1912 6254
rect 1860 6190 1912 6196
rect 1584 5772 1636 5778
rect 1584 5714 1636 5720
rect 1768 5636 1820 5642
rect 1768 5578 1820 5584
rect 1780 5370 1808 5578
rect 1768 5364 1820 5370
rect 1768 5306 1820 5312
rect 1872 4826 1900 6190
rect 2044 5228 2096 5234
rect 2044 5170 2096 5176
rect 1860 4820 1912 4826
rect 1860 4762 1912 4768
rect 2056 4622 2084 5170
rect 2044 4616 2096 4622
rect 2044 4558 2096 4564
rect 664 4072 716 4078
rect 664 4014 716 4020
rect 1860 4072 1912 4078
rect 1860 4014 1912 4020
rect 676 800 704 4014
rect 1584 3460 1636 3466
rect 1584 3402 1636 3408
rect 1596 2825 1624 3402
rect 1872 3194 1900 4014
rect 1860 3188 1912 3194
rect 1860 3130 1912 3136
rect 1582 2816 1638 2825
rect 1582 2751 1638 2760
rect 2332 2582 2360 15438
rect 2504 7880 2556 7886
rect 2504 7822 2556 7828
rect 2516 5370 2544 7822
rect 2608 6730 2636 18702
rect 2778 17776 2834 17785
rect 2778 17711 2780 17720
rect 2832 17711 2834 17720
rect 2780 17682 2832 17688
rect 2780 16040 2832 16046
rect 2780 15982 2832 15988
rect 2792 15745 2820 15982
rect 2778 15736 2834 15745
rect 2778 15671 2834 15680
rect 2872 14340 2924 14346
rect 2872 14282 2924 14288
rect 2884 14074 2912 14282
rect 2872 14068 2924 14074
rect 2872 14010 2924 14016
rect 2976 13938 3004 36042
rect 3528 35698 3556 36178
rect 3976 36168 4028 36174
rect 3976 36110 4028 36116
rect 3988 35698 4016 36110
rect 3516 35692 3568 35698
rect 3516 35634 3568 35640
rect 3976 35692 4028 35698
rect 3976 35634 4028 35640
rect 3056 35624 3108 35630
rect 3056 35566 3108 35572
rect 3068 35290 3096 35566
rect 3056 35284 3108 35290
rect 3056 35226 3108 35232
rect 3884 35080 3936 35086
rect 3884 35022 3936 35028
rect 3514 33416 3570 33425
rect 3514 33351 3516 33360
rect 3568 33351 3570 33360
rect 3516 33322 3568 33328
rect 3424 14408 3476 14414
rect 3424 14350 3476 14356
rect 3436 14006 3464 14350
rect 3424 14000 3476 14006
rect 3424 13942 3476 13948
rect 2964 13932 3016 13938
rect 2964 13874 3016 13880
rect 2780 11688 2832 11694
rect 2778 11656 2780 11665
rect 2832 11656 2834 11665
rect 2778 11591 2834 11600
rect 2976 11150 3004 13874
rect 3424 13728 3476 13734
rect 3424 13670 3476 13676
rect 3436 13394 3464 13670
rect 3424 13388 3476 13394
rect 3424 13330 3476 13336
rect 3516 12436 3568 12442
rect 3516 12378 3568 12384
rect 3528 12345 3556 12378
rect 3514 12336 3570 12345
rect 3514 12271 3570 12280
rect 2964 11144 3016 11150
rect 2964 11086 3016 11092
rect 2976 10062 3004 11086
rect 2964 10056 3016 10062
rect 2964 9998 3016 10004
rect 2780 9512 2832 9518
rect 2780 9454 2832 9460
rect 2792 8945 2820 9454
rect 2964 9036 3016 9042
rect 2964 8978 3016 8984
rect 2778 8936 2834 8945
rect 2778 8871 2834 8880
rect 2976 8265 3004 8978
rect 3332 8424 3384 8430
rect 3332 8366 3384 8372
rect 2962 8256 3018 8265
rect 2962 8191 3018 8200
rect 3054 7576 3110 7585
rect 3054 7511 3110 7520
rect 3068 7478 3096 7511
rect 3056 7472 3108 7478
rect 3056 7414 3108 7420
rect 2872 6792 2924 6798
rect 2872 6734 2924 6740
rect 2596 6724 2648 6730
rect 2596 6666 2648 6672
rect 2780 5772 2832 5778
rect 2780 5714 2832 5720
rect 2504 5364 2556 5370
rect 2504 5306 2556 5312
rect 2792 4185 2820 5714
rect 2884 5234 2912 6734
rect 3056 6656 3108 6662
rect 3056 6598 3108 6604
rect 3068 5302 3096 6598
rect 3148 6248 3200 6254
rect 3148 6190 3200 6196
rect 3056 5296 3108 5302
rect 3056 5238 3108 5244
rect 2872 5228 2924 5234
rect 2872 5170 2924 5176
rect 3160 4865 3188 6190
rect 3146 4856 3202 4865
rect 3146 4791 3202 4800
rect 3148 4616 3200 4622
rect 3148 4558 3200 4564
rect 2778 4176 2834 4185
rect 2778 4111 2834 4120
rect 3160 3602 3188 4558
rect 3240 4004 3292 4010
rect 3240 3946 3292 3952
rect 3148 3596 3200 3602
rect 3148 3538 3200 3544
rect 2778 3496 2834 3505
rect 2504 3460 2556 3466
rect 2778 3431 2834 3440
rect 2504 3402 2556 3408
rect 2516 3194 2544 3402
rect 2504 3188 2556 3194
rect 2504 3130 2556 3136
rect 2596 2848 2648 2854
rect 2596 2790 2648 2796
rect 2320 2576 2372 2582
rect 2320 2518 2372 2524
rect 2608 800 2636 2790
rect 2792 2514 2820 3431
rect 2780 2508 2832 2514
rect 2780 2450 2832 2456
rect 3252 800 3280 3946
rect 3344 1465 3372 8366
rect 3896 7886 3924 35022
rect 4172 31822 4200 36502
rect 4423 36476 4731 36485
rect 4423 36474 4429 36476
rect 4485 36474 4509 36476
rect 4565 36474 4589 36476
rect 4645 36474 4669 36476
rect 4725 36474 4731 36476
rect 4485 36422 4487 36474
rect 4667 36422 4669 36474
rect 4423 36420 4429 36422
rect 4485 36420 4509 36422
rect 4565 36420 4589 36422
rect 4645 36420 4669 36422
rect 4725 36420 4731 36422
rect 4423 36411 4731 36420
rect 4816 36242 4844 44950
rect 6012 37262 6040 46854
rect 6000 37256 6052 37262
rect 6000 37198 6052 37204
rect 4252 36236 4304 36242
rect 4252 36178 4304 36184
rect 4804 36236 4856 36242
rect 4804 36178 4856 36184
rect 4160 31816 4212 31822
rect 4160 31758 4212 31764
rect 4264 25294 4292 36178
rect 5908 36100 5960 36106
rect 5908 36042 5960 36048
rect 5920 35766 5948 36042
rect 6748 36038 6776 46854
rect 7024 46578 7052 46990
rect 7896 46812 8204 46821
rect 7896 46810 7902 46812
rect 7958 46810 7982 46812
rect 8038 46810 8062 46812
rect 8118 46810 8142 46812
rect 8198 46810 8204 46812
rect 7958 46758 7960 46810
rect 8140 46758 8142 46810
rect 7896 46756 7902 46758
rect 7958 46756 7982 46758
rect 8038 46756 8062 46758
rect 8118 46756 8142 46758
rect 8198 46756 8204 46758
rect 7896 46747 8204 46756
rect 7012 46572 7064 46578
rect 7012 46514 7064 46520
rect 8404 46510 8432 49200
rect 10336 47122 10364 49200
rect 10324 47116 10376 47122
rect 10324 47058 10376 47064
rect 9312 47048 9364 47054
rect 9312 46990 9364 46996
rect 7840 46504 7892 46510
rect 7840 46446 7892 46452
rect 8392 46504 8444 46510
rect 8392 46446 8444 46452
rect 7852 46170 7880 46446
rect 7840 46164 7892 46170
rect 7840 46106 7892 46112
rect 7748 45960 7800 45966
rect 7748 45902 7800 45908
rect 6736 36032 6788 36038
rect 6736 35974 6788 35980
rect 5908 35760 5960 35766
rect 5908 35702 5960 35708
rect 4344 35624 4396 35630
rect 4344 35566 4396 35572
rect 4356 33998 4384 35566
rect 4423 35388 4731 35397
rect 4423 35386 4429 35388
rect 4485 35386 4509 35388
rect 4565 35386 4589 35388
rect 4645 35386 4669 35388
rect 4725 35386 4731 35388
rect 4485 35334 4487 35386
rect 4667 35334 4669 35386
rect 4423 35332 4429 35334
rect 4485 35332 4509 35334
rect 4565 35332 4589 35334
rect 4645 35332 4669 35334
rect 4725 35332 4731 35334
rect 4423 35323 4731 35332
rect 5920 35086 5948 35702
rect 7760 35698 7788 45902
rect 7896 45724 8204 45733
rect 7896 45722 7902 45724
rect 7958 45722 7982 45724
rect 8038 45722 8062 45724
rect 8118 45722 8142 45724
rect 8198 45722 8204 45724
rect 7958 45670 7960 45722
rect 8140 45670 8142 45722
rect 7896 45668 7902 45670
rect 7958 45668 7982 45670
rect 8038 45668 8062 45670
rect 8118 45668 8142 45670
rect 8198 45668 8204 45670
rect 7896 45659 8204 45668
rect 9324 45490 9352 46990
rect 9864 46980 9916 46986
rect 9864 46922 9916 46928
rect 9876 46170 9904 46922
rect 10980 46510 11008 49200
rect 11624 47546 11652 49200
rect 13556 47954 13584 49200
rect 13464 47926 13584 47954
rect 11624 47518 11836 47546
rect 11369 47356 11677 47365
rect 11369 47354 11375 47356
rect 11431 47354 11455 47356
rect 11511 47354 11535 47356
rect 11591 47354 11615 47356
rect 11671 47354 11677 47356
rect 11431 47302 11433 47354
rect 11613 47302 11615 47354
rect 11369 47300 11375 47302
rect 11431 47300 11455 47302
rect 11511 47300 11535 47302
rect 11591 47300 11615 47302
rect 11671 47300 11677 47302
rect 11369 47291 11677 47300
rect 11704 47048 11756 47054
rect 11704 46990 11756 46996
rect 10508 46504 10560 46510
rect 10508 46446 10560 46452
rect 10968 46504 11020 46510
rect 10968 46446 11020 46452
rect 10324 46436 10376 46442
rect 10324 46378 10376 46384
rect 9864 46164 9916 46170
rect 9864 46106 9916 46112
rect 9956 45960 10008 45966
rect 9956 45902 10008 45908
rect 9312 45484 9364 45490
rect 9312 45426 9364 45432
rect 9968 45422 9996 45902
rect 10336 45490 10364 46378
rect 10520 46170 10548 46446
rect 10600 46368 10652 46374
rect 10600 46310 10652 46316
rect 10508 46164 10560 46170
rect 10508 46106 10560 46112
rect 10612 45966 10640 46310
rect 11369 46268 11677 46277
rect 11369 46266 11375 46268
rect 11431 46266 11455 46268
rect 11511 46266 11535 46268
rect 11591 46266 11615 46268
rect 11671 46266 11677 46268
rect 11431 46214 11433 46266
rect 11613 46214 11615 46266
rect 11369 46212 11375 46214
rect 11431 46212 11455 46214
rect 11511 46212 11535 46214
rect 11591 46212 11615 46214
rect 11671 46212 11677 46214
rect 11369 46203 11677 46212
rect 11716 46034 11744 46990
rect 11808 46034 11836 47518
rect 13464 46510 13492 47926
rect 13912 47048 13964 47054
rect 13912 46990 13964 46996
rect 14372 47048 14424 47054
rect 14844 47002 14872 49200
rect 14372 46990 14424 46996
rect 13924 46578 13952 46990
rect 14384 46578 14412 46990
rect 14752 46974 14872 47002
rect 13912 46572 13964 46578
rect 13912 46514 13964 46520
rect 14372 46572 14424 46578
rect 14372 46514 14424 46520
rect 14752 46510 14780 46974
rect 14842 46812 15150 46821
rect 14842 46810 14848 46812
rect 14904 46810 14928 46812
rect 14984 46810 15008 46812
rect 15064 46810 15088 46812
rect 15144 46810 15150 46812
rect 14904 46758 14906 46810
rect 15086 46758 15088 46810
rect 14842 46756 14848 46758
rect 14904 46756 14928 46758
rect 14984 46756 15008 46758
rect 15064 46756 15088 46758
rect 15144 46756 15150 46758
rect 14842 46747 15150 46756
rect 13452 46504 13504 46510
rect 13452 46446 13504 46452
rect 13544 46504 13596 46510
rect 13544 46446 13596 46452
rect 14556 46504 14608 46510
rect 14556 46446 14608 46452
rect 14740 46504 14792 46510
rect 14740 46446 14792 46452
rect 16396 46504 16448 46510
rect 16396 46446 16448 46452
rect 13556 46170 13584 46446
rect 14568 46170 14596 46446
rect 16408 46170 16436 46446
rect 16776 46442 16804 49200
rect 18315 47356 18623 47365
rect 18315 47354 18321 47356
rect 18377 47354 18401 47356
rect 18457 47354 18481 47356
rect 18537 47354 18561 47356
rect 18617 47354 18623 47356
rect 18377 47302 18379 47354
rect 18559 47302 18561 47354
rect 18315 47300 18321 47302
rect 18377 47300 18401 47302
rect 18457 47300 18481 47302
rect 18537 47300 18561 47302
rect 18617 47300 18623 47302
rect 18315 47291 18623 47300
rect 16856 47048 16908 47054
rect 16856 46990 16908 46996
rect 18512 47048 18564 47054
rect 18512 46990 18564 46996
rect 16868 46578 16896 46990
rect 18524 46578 18552 46990
rect 16856 46572 16908 46578
rect 16856 46514 16908 46520
rect 18512 46572 18564 46578
rect 18512 46514 18564 46520
rect 18708 46442 18736 49200
rect 19340 46504 19392 46510
rect 19340 46446 19392 46452
rect 16764 46436 16816 46442
rect 16764 46378 16816 46384
rect 18696 46436 18748 46442
rect 18696 46378 18748 46384
rect 18144 46368 18196 46374
rect 18144 46310 18196 46316
rect 13544 46164 13596 46170
rect 13544 46106 13596 46112
rect 14556 46164 14608 46170
rect 14556 46106 14608 46112
rect 16396 46164 16448 46170
rect 16396 46106 16448 46112
rect 11704 46028 11756 46034
rect 11704 45970 11756 45976
rect 11796 46028 11848 46034
rect 11796 45970 11848 45976
rect 18156 45966 18184 46310
rect 18315 46268 18623 46277
rect 18315 46266 18321 46268
rect 18377 46266 18401 46268
rect 18457 46266 18481 46268
rect 18537 46266 18561 46268
rect 18617 46266 18623 46268
rect 18377 46214 18379 46266
rect 18559 46214 18561 46266
rect 18315 46212 18321 46214
rect 18377 46212 18401 46214
rect 18457 46212 18481 46214
rect 18537 46212 18561 46214
rect 18617 46212 18623 46214
rect 18315 46203 18623 46212
rect 19352 46170 19380 46446
rect 19340 46164 19392 46170
rect 19340 46106 19392 46112
rect 19996 46034 20024 49200
rect 20812 47048 20864 47054
rect 20812 46990 20864 46996
rect 20824 46578 20852 46990
rect 20812 46572 20864 46578
rect 20812 46514 20864 46520
rect 21284 46442 21312 49200
rect 22192 47184 22244 47190
rect 22192 47126 22244 47132
rect 21788 46812 22096 46821
rect 21788 46810 21794 46812
rect 21850 46810 21874 46812
rect 21930 46810 21954 46812
rect 22010 46810 22034 46812
rect 22090 46810 22096 46812
rect 21850 46758 21852 46810
rect 22032 46758 22034 46810
rect 21788 46756 21794 46758
rect 21850 46756 21874 46758
rect 21930 46756 21954 46758
rect 22010 46756 22034 46758
rect 22090 46756 22096 46758
rect 21788 46747 22096 46756
rect 21272 46436 21324 46442
rect 21272 46378 21324 46384
rect 22204 46102 22232 47126
rect 22468 47116 22520 47122
rect 22468 47058 22520 47064
rect 22376 46504 22428 46510
rect 22376 46446 22428 46452
rect 22192 46096 22244 46102
rect 22192 46038 22244 46044
rect 19984 46028 20036 46034
rect 19984 45970 20036 45976
rect 10600 45960 10652 45966
rect 10600 45902 10652 45908
rect 13636 45960 13688 45966
rect 13636 45902 13688 45908
rect 14464 45960 14516 45966
rect 14464 45902 14516 45908
rect 18144 45960 18196 45966
rect 18144 45902 18196 45908
rect 19432 45960 19484 45966
rect 19432 45902 19484 45908
rect 11796 45892 11848 45898
rect 11796 45834 11848 45840
rect 11808 45626 11836 45834
rect 11796 45620 11848 45626
rect 11796 45562 11848 45568
rect 13648 45558 13676 45902
rect 13636 45552 13688 45558
rect 13636 45494 13688 45500
rect 10324 45484 10376 45490
rect 10324 45426 10376 45432
rect 11888 45484 11940 45490
rect 11888 45426 11940 45432
rect 9956 45416 10008 45422
rect 9956 45358 10008 45364
rect 11369 45180 11677 45189
rect 11369 45178 11375 45180
rect 11431 45178 11455 45180
rect 11511 45178 11535 45180
rect 11591 45178 11615 45180
rect 11671 45178 11677 45180
rect 11431 45126 11433 45178
rect 11613 45126 11615 45178
rect 11369 45124 11375 45126
rect 11431 45124 11455 45126
rect 11511 45124 11535 45126
rect 11591 45124 11615 45126
rect 11671 45124 11677 45126
rect 11369 45115 11677 45124
rect 7896 44636 8204 44645
rect 7896 44634 7902 44636
rect 7958 44634 7982 44636
rect 8038 44634 8062 44636
rect 8118 44634 8142 44636
rect 8198 44634 8204 44636
rect 7958 44582 7960 44634
rect 8140 44582 8142 44634
rect 7896 44580 7902 44582
rect 7958 44580 7982 44582
rect 8038 44580 8062 44582
rect 8118 44580 8142 44582
rect 8198 44580 8204 44582
rect 7896 44571 8204 44580
rect 11369 44092 11677 44101
rect 11369 44090 11375 44092
rect 11431 44090 11455 44092
rect 11511 44090 11535 44092
rect 11591 44090 11615 44092
rect 11671 44090 11677 44092
rect 11431 44038 11433 44090
rect 11613 44038 11615 44090
rect 11369 44036 11375 44038
rect 11431 44036 11455 44038
rect 11511 44036 11535 44038
rect 11591 44036 11615 44038
rect 11671 44036 11677 44038
rect 11369 44027 11677 44036
rect 11900 43858 11928 45426
rect 11888 43852 11940 43858
rect 11888 43794 11940 43800
rect 7896 43548 8204 43557
rect 7896 43546 7902 43548
rect 7958 43546 7982 43548
rect 8038 43546 8062 43548
rect 8118 43546 8142 43548
rect 8198 43546 8204 43548
rect 7958 43494 7960 43546
rect 8140 43494 8142 43546
rect 7896 43492 7902 43494
rect 7958 43492 7982 43494
rect 8038 43492 8062 43494
rect 8118 43492 8142 43494
rect 8198 43492 8204 43494
rect 7896 43483 8204 43492
rect 11369 43004 11677 43013
rect 11369 43002 11375 43004
rect 11431 43002 11455 43004
rect 11511 43002 11535 43004
rect 11591 43002 11615 43004
rect 11671 43002 11677 43004
rect 11431 42950 11433 43002
rect 11613 42950 11615 43002
rect 11369 42948 11375 42950
rect 11431 42948 11455 42950
rect 11511 42948 11535 42950
rect 11591 42948 11615 42950
rect 11671 42948 11677 42950
rect 11369 42939 11677 42948
rect 7896 42460 8204 42469
rect 7896 42458 7902 42460
rect 7958 42458 7982 42460
rect 8038 42458 8062 42460
rect 8118 42458 8142 42460
rect 8198 42458 8204 42460
rect 7958 42406 7960 42458
rect 8140 42406 8142 42458
rect 7896 42404 7902 42406
rect 7958 42404 7982 42406
rect 8038 42404 8062 42406
rect 8118 42404 8142 42406
rect 8198 42404 8204 42406
rect 7896 42395 8204 42404
rect 11369 41916 11677 41925
rect 11369 41914 11375 41916
rect 11431 41914 11455 41916
rect 11511 41914 11535 41916
rect 11591 41914 11615 41916
rect 11671 41914 11677 41916
rect 11431 41862 11433 41914
rect 11613 41862 11615 41914
rect 11369 41860 11375 41862
rect 11431 41860 11455 41862
rect 11511 41860 11535 41862
rect 11591 41860 11615 41862
rect 11671 41860 11677 41862
rect 11369 41851 11677 41860
rect 7896 41372 8204 41381
rect 7896 41370 7902 41372
rect 7958 41370 7982 41372
rect 8038 41370 8062 41372
rect 8118 41370 8142 41372
rect 8198 41370 8204 41372
rect 7958 41318 7960 41370
rect 8140 41318 8142 41370
rect 7896 41316 7902 41318
rect 7958 41316 7982 41318
rect 8038 41316 8062 41318
rect 8118 41316 8142 41318
rect 8198 41316 8204 41318
rect 7896 41307 8204 41316
rect 11369 40828 11677 40837
rect 11369 40826 11375 40828
rect 11431 40826 11455 40828
rect 11511 40826 11535 40828
rect 11591 40826 11615 40828
rect 11671 40826 11677 40828
rect 11431 40774 11433 40826
rect 11613 40774 11615 40826
rect 11369 40772 11375 40774
rect 11431 40772 11455 40774
rect 11511 40772 11535 40774
rect 11591 40772 11615 40774
rect 11671 40772 11677 40774
rect 11369 40763 11677 40772
rect 7896 40284 8204 40293
rect 7896 40282 7902 40284
rect 7958 40282 7982 40284
rect 8038 40282 8062 40284
rect 8118 40282 8142 40284
rect 8198 40282 8204 40284
rect 7958 40230 7960 40282
rect 8140 40230 8142 40282
rect 7896 40228 7902 40230
rect 7958 40228 7982 40230
rect 8038 40228 8062 40230
rect 8118 40228 8142 40230
rect 8198 40228 8204 40230
rect 7896 40219 8204 40228
rect 11369 39740 11677 39749
rect 11369 39738 11375 39740
rect 11431 39738 11455 39740
rect 11511 39738 11535 39740
rect 11591 39738 11615 39740
rect 11671 39738 11677 39740
rect 11431 39686 11433 39738
rect 11613 39686 11615 39738
rect 11369 39684 11375 39686
rect 11431 39684 11455 39686
rect 11511 39684 11535 39686
rect 11591 39684 11615 39686
rect 11671 39684 11677 39686
rect 11369 39675 11677 39684
rect 7896 39196 8204 39205
rect 7896 39194 7902 39196
rect 7958 39194 7982 39196
rect 8038 39194 8062 39196
rect 8118 39194 8142 39196
rect 8198 39194 8204 39196
rect 7958 39142 7960 39194
rect 8140 39142 8142 39194
rect 7896 39140 7902 39142
rect 7958 39140 7982 39142
rect 8038 39140 8062 39142
rect 8118 39140 8142 39142
rect 8198 39140 8204 39142
rect 7896 39131 8204 39140
rect 11369 38652 11677 38661
rect 11369 38650 11375 38652
rect 11431 38650 11455 38652
rect 11511 38650 11535 38652
rect 11591 38650 11615 38652
rect 11671 38650 11677 38652
rect 11431 38598 11433 38650
rect 11613 38598 11615 38650
rect 11369 38596 11375 38598
rect 11431 38596 11455 38598
rect 11511 38596 11535 38598
rect 11591 38596 11615 38598
rect 11671 38596 11677 38598
rect 11369 38587 11677 38596
rect 7896 38108 8204 38117
rect 7896 38106 7902 38108
rect 7958 38106 7982 38108
rect 8038 38106 8062 38108
rect 8118 38106 8142 38108
rect 8198 38106 8204 38108
rect 7958 38054 7960 38106
rect 8140 38054 8142 38106
rect 7896 38052 7902 38054
rect 7958 38052 7982 38054
rect 8038 38052 8062 38054
rect 8118 38052 8142 38054
rect 8198 38052 8204 38054
rect 7896 38043 8204 38052
rect 11369 37564 11677 37573
rect 11369 37562 11375 37564
rect 11431 37562 11455 37564
rect 11511 37562 11535 37564
rect 11591 37562 11615 37564
rect 11671 37562 11677 37564
rect 11431 37510 11433 37562
rect 11613 37510 11615 37562
rect 11369 37508 11375 37510
rect 11431 37508 11455 37510
rect 11511 37508 11535 37510
rect 11591 37508 11615 37510
rect 11671 37508 11677 37510
rect 11369 37499 11677 37508
rect 7896 37020 8204 37029
rect 7896 37018 7902 37020
rect 7958 37018 7982 37020
rect 8038 37018 8062 37020
rect 8118 37018 8142 37020
rect 8198 37018 8204 37020
rect 7958 36966 7960 37018
rect 8140 36966 8142 37018
rect 7896 36964 7902 36966
rect 7958 36964 7982 36966
rect 8038 36964 8062 36966
rect 8118 36964 8142 36966
rect 8198 36964 8204 36966
rect 7896 36955 8204 36964
rect 9588 36712 9640 36718
rect 9588 36654 9640 36660
rect 9600 36106 9628 36654
rect 10692 36576 10744 36582
rect 10692 36518 10744 36524
rect 9588 36100 9640 36106
rect 9588 36042 9640 36048
rect 9772 36100 9824 36106
rect 9772 36042 9824 36048
rect 7896 35932 8204 35941
rect 7896 35930 7902 35932
rect 7958 35930 7982 35932
rect 8038 35930 8062 35932
rect 8118 35930 8142 35932
rect 8198 35930 8204 35932
rect 7958 35878 7960 35930
rect 8140 35878 8142 35930
rect 9784 35894 9812 36042
rect 7896 35876 7902 35878
rect 7958 35876 7982 35878
rect 8038 35876 8062 35878
rect 8118 35876 8142 35878
rect 8198 35876 8204 35878
rect 7896 35867 8204 35876
rect 9600 35866 9812 35894
rect 7748 35692 7800 35698
rect 7748 35634 7800 35640
rect 5908 35080 5960 35086
rect 5908 35022 5960 35028
rect 7896 34844 8204 34853
rect 7896 34842 7902 34844
rect 7958 34842 7982 34844
rect 8038 34842 8062 34844
rect 8118 34842 8142 34844
rect 8198 34842 8204 34844
rect 7958 34790 7960 34842
rect 8140 34790 8142 34842
rect 7896 34788 7902 34790
rect 7958 34788 7982 34790
rect 8038 34788 8062 34790
rect 8118 34788 8142 34790
rect 8198 34788 8204 34790
rect 7896 34779 8204 34788
rect 4423 34300 4731 34309
rect 4423 34298 4429 34300
rect 4485 34298 4509 34300
rect 4565 34298 4589 34300
rect 4645 34298 4669 34300
rect 4725 34298 4731 34300
rect 4485 34246 4487 34298
rect 4667 34246 4669 34298
rect 4423 34244 4429 34246
rect 4485 34244 4509 34246
rect 4565 34244 4589 34246
rect 4645 34244 4669 34246
rect 4725 34244 4731 34246
rect 4423 34235 4731 34244
rect 4344 33992 4396 33998
rect 4344 33934 4396 33940
rect 7896 33756 8204 33765
rect 7896 33754 7902 33756
rect 7958 33754 7982 33756
rect 8038 33754 8062 33756
rect 8118 33754 8142 33756
rect 8198 33754 8204 33756
rect 7958 33702 7960 33754
rect 8140 33702 8142 33754
rect 7896 33700 7902 33702
rect 7958 33700 7982 33702
rect 8038 33700 8062 33702
rect 8118 33700 8142 33702
rect 8198 33700 8204 33702
rect 7896 33691 8204 33700
rect 9128 33380 9180 33386
rect 9128 33322 9180 33328
rect 4423 33212 4731 33221
rect 4423 33210 4429 33212
rect 4485 33210 4509 33212
rect 4565 33210 4589 33212
rect 4645 33210 4669 33212
rect 4725 33210 4731 33212
rect 4485 33158 4487 33210
rect 4667 33158 4669 33210
rect 4423 33156 4429 33158
rect 4485 33156 4509 33158
rect 4565 33156 4589 33158
rect 4645 33156 4669 33158
rect 4725 33156 4731 33158
rect 4423 33147 4731 33156
rect 7896 32668 8204 32677
rect 7896 32666 7902 32668
rect 7958 32666 7982 32668
rect 8038 32666 8062 32668
rect 8118 32666 8142 32668
rect 8198 32666 8204 32668
rect 7958 32614 7960 32666
rect 8140 32614 8142 32666
rect 7896 32612 7902 32614
rect 7958 32612 7982 32614
rect 8038 32612 8062 32614
rect 8118 32612 8142 32614
rect 8198 32612 8204 32614
rect 7896 32603 8204 32612
rect 4423 32124 4731 32133
rect 4423 32122 4429 32124
rect 4485 32122 4509 32124
rect 4565 32122 4589 32124
rect 4645 32122 4669 32124
rect 4725 32122 4731 32124
rect 4485 32070 4487 32122
rect 4667 32070 4669 32122
rect 4423 32068 4429 32070
rect 4485 32068 4509 32070
rect 4565 32068 4589 32070
rect 4645 32068 4669 32070
rect 4725 32068 4731 32070
rect 4423 32059 4731 32068
rect 7896 31580 8204 31589
rect 7896 31578 7902 31580
rect 7958 31578 7982 31580
rect 8038 31578 8062 31580
rect 8118 31578 8142 31580
rect 8198 31578 8204 31580
rect 7958 31526 7960 31578
rect 8140 31526 8142 31578
rect 7896 31524 7902 31526
rect 7958 31524 7982 31526
rect 8038 31524 8062 31526
rect 8118 31524 8142 31526
rect 8198 31524 8204 31526
rect 7896 31515 8204 31524
rect 4423 31036 4731 31045
rect 4423 31034 4429 31036
rect 4485 31034 4509 31036
rect 4565 31034 4589 31036
rect 4645 31034 4669 31036
rect 4725 31034 4731 31036
rect 4485 30982 4487 31034
rect 4667 30982 4669 31034
rect 4423 30980 4429 30982
rect 4485 30980 4509 30982
rect 4565 30980 4589 30982
rect 4645 30980 4669 30982
rect 4725 30980 4731 30982
rect 4423 30971 4731 30980
rect 9140 30734 9168 33322
rect 9128 30728 9180 30734
rect 9128 30670 9180 30676
rect 9600 30666 9628 35866
rect 9588 30660 9640 30666
rect 9588 30602 9640 30608
rect 9956 30660 10008 30666
rect 9956 30602 10008 30608
rect 7896 30492 8204 30501
rect 7896 30490 7902 30492
rect 7958 30490 7982 30492
rect 8038 30490 8062 30492
rect 8118 30490 8142 30492
rect 8198 30490 8204 30492
rect 7958 30438 7960 30490
rect 8140 30438 8142 30490
rect 7896 30436 7902 30438
rect 7958 30436 7982 30438
rect 8038 30436 8062 30438
rect 8118 30436 8142 30438
rect 8198 30436 8204 30438
rect 7896 30427 8204 30436
rect 4423 29948 4731 29957
rect 4423 29946 4429 29948
rect 4485 29946 4509 29948
rect 4565 29946 4589 29948
rect 4645 29946 4669 29948
rect 4725 29946 4731 29948
rect 4485 29894 4487 29946
rect 4667 29894 4669 29946
rect 4423 29892 4429 29894
rect 4485 29892 4509 29894
rect 4565 29892 4589 29894
rect 4645 29892 4669 29894
rect 4725 29892 4731 29894
rect 4423 29883 4731 29892
rect 7896 29404 8204 29413
rect 7896 29402 7902 29404
rect 7958 29402 7982 29404
rect 8038 29402 8062 29404
rect 8118 29402 8142 29404
rect 8198 29402 8204 29404
rect 7958 29350 7960 29402
rect 8140 29350 8142 29402
rect 7896 29348 7902 29350
rect 7958 29348 7982 29350
rect 8038 29348 8062 29350
rect 8118 29348 8142 29350
rect 8198 29348 8204 29350
rect 7896 29339 8204 29348
rect 4423 28860 4731 28869
rect 4423 28858 4429 28860
rect 4485 28858 4509 28860
rect 4565 28858 4589 28860
rect 4645 28858 4669 28860
rect 4725 28858 4731 28860
rect 4485 28806 4487 28858
rect 4667 28806 4669 28858
rect 4423 28804 4429 28806
rect 4485 28804 4509 28806
rect 4565 28804 4589 28806
rect 4645 28804 4669 28806
rect 4725 28804 4731 28806
rect 4423 28795 4731 28804
rect 7896 28316 8204 28325
rect 7896 28314 7902 28316
rect 7958 28314 7982 28316
rect 8038 28314 8062 28316
rect 8118 28314 8142 28316
rect 8198 28314 8204 28316
rect 7958 28262 7960 28314
rect 8140 28262 8142 28314
rect 7896 28260 7902 28262
rect 7958 28260 7982 28262
rect 8038 28260 8062 28262
rect 8118 28260 8142 28262
rect 8198 28260 8204 28262
rect 7896 28251 8204 28260
rect 4423 27772 4731 27781
rect 4423 27770 4429 27772
rect 4485 27770 4509 27772
rect 4565 27770 4589 27772
rect 4645 27770 4669 27772
rect 4725 27770 4731 27772
rect 4485 27718 4487 27770
rect 4667 27718 4669 27770
rect 4423 27716 4429 27718
rect 4485 27716 4509 27718
rect 4565 27716 4589 27718
rect 4645 27716 4669 27718
rect 4725 27716 4731 27718
rect 4423 27707 4731 27716
rect 7896 27228 8204 27237
rect 7896 27226 7902 27228
rect 7958 27226 7982 27228
rect 8038 27226 8062 27228
rect 8118 27226 8142 27228
rect 8198 27226 8204 27228
rect 7958 27174 7960 27226
rect 8140 27174 8142 27226
rect 7896 27172 7902 27174
rect 7958 27172 7982 27174
rect 8038 27172 8062 27174
rect 8118 27172 8142 27174
rect 8198 27172 8204 27174
rect 7896 27163 8204 27172
rect 4423 26684 4731 26693
rect 4423 26682 4429 26684
rect 4485 26682 4509 26684
rect 4565 26682 4589 26684
rect 4645 26682 4669 26684
rect 4725 26682 4731 26684
rect 4485 26630 4487 26682
rect 4667 26630 4669 26682
rect 4423 26628 4429 26630
rect 4485 26628 4509 26630
rect 4565 26628 4589 26630
rect 4645 26628 4669 26630
rect 4725 26628 4731 26630
rect 4423 26619 4731 26628
rect 7896 26140 8204 26149
rect 7896 26138 7902 26140
rect 7958 26138 7982 26140
rect 8038 26138 8062 26140
rect 8118 26138 8142 26140
rect 8198 26138 8204 26140
rect 7958 26086 7960 26138
rect 8140 26086 8142 26138
rect 7896 26084 7902 26086
rect 7958 26084 7982 26086
rect 8038 26084 8062 26086
rect 8118 26084 8142 26086
rect 8198 26084 8204 26086
rect 7896 26075 8204 26084
rect 4423 25596 4731 25605
rect 4423 25594 4429 25596
rect 4485 25594 4509 25596
rect 4565 25594 4589 25596
rect 4645 25594 4669 25596
rect 4725 25594 4731 25596
rect 4485 25542 4487 25594
rect 4667 25542 4669 25594
rect 4423 25540 4429 25542
rect 4485 25540 4509 25542
rect 4565 25540 4589 25542
rect 4645 25540 4669 25542
rect 4725 25540 4731 25542
rect 4423 25531 4731 25540
rect 4252 25288 4304 25294
rect 4252 25230 4304 25236
rect 7896 25052 8204 25061
rect 7896 25050 7902 25052
rect 7958 25050 7982 25052
rect 8038 25050 8062 25052
rect 8118 25050 8142 25052
rect 8198 25050 8204 25052
rect 7958 24998 7960 25050
rect 8140 24998 8142 25050
rect 7896 24996 7902 24998
rect 7958 24996 7982 24998
rect 8038 24996 8062 24998
rect 8118 24996 8142 24998
rect 8198 24996 8204 24998
rect 7896 24987 8204 24996
rect 4423 24508 4731 24517
rect 4423 24506 4429 24508
rect 4485 24506 4509 24508
rect 4565 24506 4589 24508
rect 4645 24506 4669 24508
rect 4725 24506 4731 24508
rect 4485 24454 4487 24506
rect 4667 24454 4669 24506
rect 4423 24452 4429 24454
rect 4485 24452 4509 24454
rect 4565 24452 4589 24454
rect 4645 24452 4669 24454
rect 4725 24452 4731 24454
rect 4423 24443 4731 24452
rect 9404 24064 9456 24070
rect 9404 24006 9456 24012
rect 7896 23964 8204 23973
rect 7896 23962 7902 23964
rect 7958 23962 7982 23964
rect 8038 23962 8062 23964
rect 8118 23962 8142 23964
rect 8198 23962 8204 23964
rect 7958 23910 7960 23962
rect 8140 23910 8142 23962
rect 7896 23908 7902 23910
rect 7958 23908 7982 23910
rect 8038 23908 8062 23910
rect 8118 23908 8142 23910
rect 8198 23908 8204 23910
rect 7896 23899 8204 23908
rect 4423 23420 4731 23429
rect 4423 23418 4429 23420
rect 4485 23418 4509 23420
rect 4565 23418 4589 23420
rect 4645 23418 4669 23420
rect 4725 23418 4731 23420
rect 4485 23366 4487 23418
rect 4667 23366 4669 23418
rect 4423 23364 4429 23366
rect 4485 23364 4509 23366
rect 4565 23364 4589 23366
rect 4645 23364 4669 23366
rect 4725 23364 4731 23366
rect 4423 23355 4731 23364
rect 7896 22876 8204 22885
rect 7896 22874 7902 22876
rect 7958 22874 7982 22876
rect 8038 22874 8062 22876
rect 8118 22874 8142 22876
rect 8198 22874 8204 22876
rect 7958 22822 7960 22874
rect 8140 22822 8142 22874
rect 7896 22820 7902 22822
rect 7958 22820 7982 22822
rect 8038 22820 8062 22822
rect 8118 22820 8142 22822
rect 8198 22820 8204 22822
rect 7896 22811 8204 22820
rect 4423 22332 4731 22341
rect 4423 22330 4429 22332
rect 4485 22330 4509 22332
rect 4565 22330 4589 22332
rect 4645 22330 4669 22332
rect 4725 22330 4731 22332
rect 4485 22278 4487 22330
rect 4667 22278 4669 22330
rect 4423 22276 4429 22278
rect 4485 22276 4509 22278
rect 4565 22276 4589 22278
rect 4645 22276 4669 22278
rect 4725 22276 4731 22278
rect 4423 22267 4731 22276
rect 7896 21788 8204 21797
rect 7896 21786 7902 21788
rect 7958 21786 7982 21788
rect 8038 21786 8062 21788
rect 8118 21786 8142 21788
rect 8198 21786 8204 21788
rect 7958 21734 7960 21786
rect 8140 21734 8142 21786
rect 7896 21732 7902 21734
rect 7958 21732 7982 21734
rect 8038 21732 8062 21734
rect 8118 21732 8142 21734
rect 8198 21732 8204 21734
rect 7896 21723 8204 21732
rect 4423 21244 4731 21253
rect 4423 21242 4429 21244
rect 4485 21242 4509 21244
rect 4565 21242 4589 21244
rect 4645 21242 4669 21244
rect 4725 21242 4731 21244
rect 4485 21190 4487 21242
rect 4667 21190 4669 21242
rect 4423 21188 4429 21190
rect 4485 21188 4509 21190
rect 4565 21188 4589 21190
rect 4645 21188 4669 21190
rect 4725 21188 4731 21190
rect 4423 21179 4731 21188
rect 7896 20700 8204 20709
rect 7896 20698 7902 20700
rect 7958 20698 7982 20700
rect 8038 20698 8062 20700
rect 8118 20698 8142 20700
rect 8198 20698 8204 20700
rect 7958 20646 7960 20698
rect 8140 20646 8142 20698
rect 7896 20644 7902 20646
rect 7958 20644 7982 20646
rect 8038 20644 8062 20646
rect 8118 20644 8142 20646
rect 8198 20644 8204 20646
rect 7896 20635 8204 20644
rect 4423 20156 4731 20165
rect 4423 20154 4429 20156
rect 4485 20154 4509 20156
rect 4565 20154 4589 20156
rect 4645 20154 4669 20156
rect 4725 20154 4731 20156
rect 4485 20102 4487 20154
rect 4667 20102 4669 20154
rect 4423 20100 4429 20102
rect 4485 20100 4509 20102
rect 4565 20100 4589 20102
rect 4645 20100 4669 20102
rect 4725 20100 4731 20102
rect 4423 20091 4731 20100
rect 7896 19612 8204 19621
rect 7896 19610 7902 19612
rect 7958 19610 7982 19612
rect 8038 19610 8062 19612
rect 8118 19610 8142 19612
rect 8198 19610 8204 19612
rect 7958 19558 7960 19610
rect 8140 19558 8142 19610
rect 7896 19556 7902 19558
rect 7958 19556 7982 19558
rect 8038 19556 8062 19558
rect 8118 19556 8142 19558
rect 8198 19556 8204 19558
rect 7896 19547 8204 19556
rect 4423 19068 4731 19077
rect 4423 19066 4429 19068
rect 4485 19066 4509 19068
rect 4565 19066 4589 19068
rect 4645 19066 4669 19068
rect 4725 19066 4731 19068
rect 4485 19014 4487 19066
rect 4667 19014 4669 19066
rect 4423 19012 4429 19014
rect 4485 19012 4509 19014
rect 4565 19012 4589 19014
rect 4645 19012 4669 19014
rect 4725 19012 4731 19014
rect 4423 19003 4731 19012
rect 7896 18524 8204 18533
rect 7896 18522 7902 18524
rect 7958 18522 7982 18524
rect 8038 18522 8062 18524
rect 8118 18522 8142 18524
rect 8198 18522 8204 18524
rect 7958 18470 7960 18522
rect 8140 18470 8142 18522
rect 7896 18468 7902 18470
rect 7958 18468 7982 18470
rect 8038 18468 8062 18470
rect 8118 18468 8142 18470
rect 8198 18468 8204 18470
rect 7896 18459 8204 18468
rect 4423 17980 4731 17989
rect 4423 17978 4429 17980
rect 4485 17978 4509 17980
rect 4565 17978 4589 17980
rect 4645 17978 4669 17980
rect 4725 17978 4731 17980
rect 4485 17926 4487 17978
rect 4667 17926 4669 17978
rect 4423 17924 4429 17926
rect 4485 17924 4509 17926
rect 4565 17924 4589 17926
rect 4645 17924 4669 17926
rect 4725 17924 4731 17926
rect 4423 17915 4731 17924
rect 7748 17536 7800 17542
rect 7748 17478 7800 17484
rect 4344 17196 4396 17202
rect 4344 17138 4396 17144
rect 4356 11218 4384 17138
rect 4423 16892 4731 16901
rect 4423 16890 4429 16892
rect 4485 16890 4509 16892
rect 4565 16890 4589 16892
rect 4645 16890 4669 16892
rect 4725 16890 4731 16892
rect 4485 16838 4487 16890
rect 4667 16838 4669 16890
rect 4423 16836 4429 16838
rect 4485 16836 4509 16838
rect 4565 16836 4589 16838
rect 4645 16836 4669 16838
rect 4725 16836 4731 16838
rect 4423 16827 4731 16836
rect 4423 15804 4731 15813
rect 4423 15802 4429 15804
rect 4485 15802 4509 15804
rect 4565 15802 4589 15804
rect 4645 15802 4669 15804
rect 4725 15802 4731 15804
rect 4485 15750 4487 15802
rect 4667 15750 4669 15802
rect 4423 15748 4429 15750
rect 4485 15748 4509 15750
rect 4565 15748 4589 15750
rect 4645 15748 4669 15750
rect 4725 15748 4731 15750
rect 4423 15739 4731 15748
rect 4423 14716 4731 14725
rect 4423 14714 4429 14716
rect 4485 14714 4509 14716
rect 4565 14714 4589 14716
rect 4645 14714 4669 14716
rect 4725 14714 4731 14716
rect 4485 14662 4487 14714
rect 4667 14662 4669 14714
rect 4423 14660 4429 14662
rect 4485 14660 4509 14662
rect 4565 14660 4589 14662
rect 4645 14660 4669 14662
rect 4725 14660 4731 14662
rect 4423 14651 4731 14660
rect 4423 13628 4731 13637
rect 4423 13626 4429 13628
rect 4485 13626 4509 13628
rect 4565 13626 4589 13628
rect 4645 13626 4669 13628
rect 4725 13626 4731 13628
rect 4485 13574 4487 13626
rect 4667 13574 4669 13626
rect 4423 13572 4429 13574
rect 4485 13572 4509 13574
rect 4565 13572 4589 13574
rect 4645 13572 4669 13574
rect 4725 13572 4731 13574
rect 4423 13563 4731 13572
rect 4988 12844 5040 12850
rect 4988 12786 5040 12792
rect 4423 12540 4731 12549
rect 4423 12538 4429 12540
rect 4485 12538 4509 12540
rect 4565 12538 4589 12540
rect 4645 12538 4669 12540
rect 4725 12538 4731 12540
rect 4485 12486 4487 12538
rect 4667 12486 4669 12538
rect 4423 12484 4429 12486
rect 4485 12484 4509 12486
rect 4565 12484 4589 12486
rect 4645 12484 4669 12486
rect 4725 12484 4731 12486
rect 4423 12475 4731 12484
rect 4423 11452 4731 11461
rect 4423 11450 4429 11452
rect 4485 11450 4509 11452
rect 4565 11450 4589 11452
rect 4645 11450 4669 11452
rect 4725 11450 4731 11452
rect 4485 11398 4487 11450
rect 4667 11398 4669 11450
rect 4423 11396 4429 11398
rect 4485 11396 4509 11398
rect 4565 11396 4589 11398
rect 4645 11396 4669 11398
rect 4725 11396 4731 11398
rect 4423 11387 4731 11396
rect 4344 11212 4396 11218
rect 4344 11154 4396 11160
rect 4068 9920 4120 9926
rect 4068 9862 4120 9868
rect 4080 8566 4108 9862
rect 4252 9376 4304 9382
rect 4252 9318 4304 9324
rect 4068 8560 4120 8566
rect 4068 8502 4120 8508
rect 4264 8498 4292 9318
rect 4356 8634 4384 11154
rect 4423 10364 4731 10373
rect 4423 10362 4429 10364
rect 4485 10362 4509 10364
rect 4565 10362 4589 10364
rect 4645 10362 4669 10364
rect 4725 10362 4731 10364
rect 4485 10310 4487 10362
rect 4667 10310 4669 10362
rect 4423 10308 4429 10310
rect 4485 10308 4509 10310
rect 4565 10308 4589 10310
rect 4645 10308 4669 10310
rect 4725 10308 4731 10310
rect 4423 10299 4731 10308
rect 4423 9276 4731 9285
rect 4423 9274 4429 9276
rect 4485 9274 4509 9276
rect 4565 9274 4589 9276
rect 4645 9274 4669 9276
rect 4725 9274 4731 9276
rect 4485 9222 4487 9274
rect 4667 9222 4669 9274
rect 4423 9220 4429 9222
rect 4485 9220 4509 9222
rect 4565 9220 4589 9222
rect 4645 9220 4669 9222
rect 4725 9220 4731 9222
rect 4423 9211 4731 9220
rect 4344 8628 4396 8634
rect 4344 8570 4396 8576
rect 4252 8492 4304 8498
rect 4252 8434 4304 8440
rect 4423 8188 4731 8197
rect 4423 8186 4429 8188
rect 4485 8186 4509 8188
rect 4565 8186 4589 8188
rect 4645 8186 4669 8188
rect 4725 8186 4731 8188
rect 4485 8134 4487 8186
rect 4667 8134 4669 8186
rect 4423 8132 4429 8134
rect 4485 8132 4509 8134
rect 4565 8132 4589 8134
rect 4645 8132 4669 8134
rect 4725 8132 4731 8134
rect 4423 8123 4731 8132
rect 3884 7880 3936 7886
rect 3936 7828 4016 7834
rect 3884 7822 4016 7828
rect 3896 7806 4016 7822
rect 3988 7002 4016 7806
rect 4896 7812 4948 7818
rect 4896 7754 4948 7760
rect 4712 7744 4764 7750
rect 4712 7686 4764 7692
rect 4724 7478 4752 7686
rect 4712 7472 4764 7478
rect 4712 7414 4764 7420
rect 4908 7410 4936 7754
rect 4896 7404 4948 7410
rect 4896 7346 4948 7352
rect 4423 7100 4731 7109
rect 4423 7098 4429 7100
rect 4485 7098 4509 7100
rect 4565 7098 4589 7100
rect 4645 7098 4669 7100
rect 4725 7098 4731 7100
rect 4485 7046 4487 7098
rect 4667 7046 4669 7098
rect 4423 7044 4429 7046
rect 4485 7044 4509 7046
rect 4565 7044 4589 7046
rect 4645 7044 4669 7046
rect 4725 7044 4731 7046
rect 4423 7035 4731 7044
rect 3976 6996 4028 7002
rect 3976 6938 4028 6944
rect 3988 6866 4016 6938
rect 3976 6860 4028 6866
rect 3976 6802 4028 6808
rect 4068 6860 4120 6866
rect 4068 6802 4120 6808
rect 3976 6248 4028 6254
rect 4080 6225 4108 6802
rect 4160 6656 4212 6662
rect 4160 6598 4212 6604
rect 4172 6390 4200 6598
rect 4160 6384 4212 6390
rect 4160 6326 4212 6332
rect 4344 6248 4396 6254
rect 3976 6190 4028 6196
rect 4066 6216 4122 6225
rect 3988 5914 4016 6190
rect 4344 6190 4396 6196
rect 4066 6151 4122 6160
rect 3976 5908 4028 5914
rect 3976 5850 4028 5856
rect 4252 5024 4304 5030
rect 4252 4966 4304 4972
rect 3976 4616 4028 4622
rect 3976 4558 4028 4564
rect 3988 4146 4016 4558
rect 4160 4480 4212 4486
rect 4160 4422 4212 4428
rect 4172 4214 4200 4422
rect 4160 4208 4212 4214
rect 4160 4150 4212 4156
rect 3976 4140 4028 4146
rect 3976 4082 4028 4088
rect 4264 3074 4292 4966
rect 3804 3046 4292 3074
rect 3804 2514 3832 3046
rect 3884 2984 3936 2990
rect 3884 2926 3936 2932
rect 3976 2984 4028 2990
rect 3976 2926 4028 2932
rect 3896 2650 3924 2926
rect 3884 2644 3936 2650
rect 3884 2586 3936 2592
rect 3792 2508 3844 2514
rect 3792 2450 3844 2456
rect 3330 1456 3386 1465
rect 3330 1391 3386 1400
rect 3988 1170 4016 2926
rect 4160 2440 4212 2446
rect 4160 2382 4212 2388
rect 4068 2304 4120 2310
rect 4068 2246 4120 2252
rect 4080 2145 4108 2246
rect 4066 2136 4122 2145
rect 4172 2106 4200 2382
rect 4066 2071 4122 2080
rect 4160 2100 4212 2106
rect 4160 2042 4212 2048
rect 3896 1142 4016 1170
rect 3896 800 3924 1142
rect 4356 1034 4384 6190
rect 4423 6012 4731 6021
rect 4423 6010 4429 6012
rect 4485 6010 4509 6012
rect 4565 6010 4589 6012
rect 4645 6010 4669 6012
rect 4725 6010 4731 6012
rect 4485 5958 4487 6010
rect 4667 5958 4669 6010
rect 4423 5956 4429 5958
rect 4485 5956 4509 5958
rect 4565 5956 4589 5958
rect 4645 5956 4669 5958
rect 4725 5956 4731 5958
rect 4423 5947 4731 5956
rect 4804 5160 4856 5166
rect 4804 5102 4856 5108
rect 4423 4924 4731 4933
rect 4423 4922 4429 4924
rect 4485 4922 4509 4924
rect 4565 4922 4589 4924
rect 4645 4922 4669 4924
rect 4725 4922 4731 4924
rect 4485 4870 4487 4922
rect 4667 4870 4669 4922
rect 4423 4868 4429 4870
rect 4485 4868 4509 4870
rect 4565 4868 4589 4870
rect 4645 4868 4669 4870
rect 4725 4868 4731 4870
rect 4423 4859 4731 4868
rect 4423 3836 4731 3845
rect 4423 3834 4429 3836
rect 4485 3834 4509 3836
rect 4565 3834 4589 3836
rect 4645 3834 4669 3836
rect 4725 3834 4731 3836
rect 4485 3782 4487 3834
rect 4667 3782 4669 3834
rect 4423 3780 4429 3782
rect 4485 3780 4509 3782
rect 4565 3780 4589 3782
rect 4645 3780 4669 3782
rect 4725 3780 4731 3782
rect 4423 3771 4731 3780
rect 4816 2854 4844 5102
rect 5000 4690 5028 12786
rect 5356 6996 5408 7002
rect 5356 6938 5408 6944
rect 5368 6798 5396 6938
rect 7760 6934 7788 17478
rect 7896 17436 8204 17445
rect 7896 17434 7902 17436
rect 7958 17434 7982 17436
rect 8038 17434 8062 17436
rect 8118 17434 8142 17436
rect 8198 17434 8204 17436
rect 7958 17382 7960 17434
rect 8140 17382 8142 17434
rect 7896 17380 7902 17382
rect 7958 17380 7982 17382
rect 8038 17380 8062 17382
rect 8118 17380 8142 17382
rect 8198 17380 8204 17382
rect 7896 17371 8204 17380
rect 7896 16348 8204 16357
rect 7896 16346 7902 16348
rect 7958 16346 7982 16348
rect 8038 16346 8062 16348
rect 8118 16346 8142 16348
rect 8198 16346 8204 16348
rect 7958 16294 7960 16346
rect 8140 16294 8142 16346
rect 7896 16292 7902 16294
rect 7958 16292 7982 16294
rect 8038 16292 8062 16294
rect 8118 16292 8142 16294
rect 8198 16292 8204 16294
rect 7896 16283 8204 16292
rect 7896 15260 8204 15269
rect 7896 15258 7902 15260
rect 7958 15258 7982 15260
rect 8038 15258 8062 15260
rect 8118 15258 8142 15260
rect 8198 15258 8204 15260
rect 7958 15206 7960 15258
rect 8140 15206 8142 15258
rect 7896 15204 7902 15206
rect 7958 15204 7982 15206
rect 8038 15204 8062 15206
rect 8118 15204 8142 15206
rect 8198 15204 8204 15206
rect 7896 15195 8204 15204
rect 7896 14172 8204 14181
rect 7896 14170 7902 14172
rect 7958 14170 7982 14172
rect 8038 14170 8062 14172
rect 8118 14170 8142 14172
rect 8198 14170 8204 14172
rect 7958 14118 7960 14170
rect 8140 14118 8142 14170
rect 7896 14116 7902 14118
rect 7958 14116 7982 14118
rect 8038 14116 8062 14118
rect 8118 14116 8142 14118
rect 8198 14116 8204 14118
rect 7896 14107 8204 14116
rect 7896 13084 8204 13093
rect 7896 13082 7902 13084
rect 7958 13082 7982 13084
rect 8038 13082 8062 13084
rect 8118 13082 8142 13084
rect 8198 13082 8204 13084
rect 7958 13030 7960 13082
rect 8140 13030 8142 13082
rect 7896 13028 7902 13030
rect 7958 13028 7982 13030
rect 8038 13028 8062 13030
rect 8118 13028 8142 13030
rect 8198 13028 8204 13030
rect 7896 13019 8204 13028
rect 7896 11996 8204 12005
rect 7896 11994 7902 11996
rect 7958 11994 7982 11996
rect 8038 11994 8062 11996
rect 8118 11994 8142 11996
rect 8198 11994 8204 11996
rect 7958 11942 7960 11994
rect 8140 11942 8142 11994
rect 7896 11940 7902 11942
rect 7958 11940 7982 11942
rect 8038 11940 8062 11942
rect 8118 11940 8142 11942
rect 8198 11940 8204 11942
rect 7896 11931 8204 11940
rect 7896 10908 8204 10917
rect 7896 10906 7902 10908
rect 7958 10906 7982 10908
rect 8038 10906 8062 10908
rect 8118 10906 8142 10908
rect 8198 10906 8204 10908
rect 7958 10854 7960 10906
rect 8140 10854 8142 10906
rect 7896 10852 7902 10854
rect 7958 10852 7982 10854
rect 8038 10852 8062 10854
rect 8118 10852 8142 10854
rect 8198 10852 8204 10854
rect 7896 10843 8204 10852
rect 7896 9820 8204 9829
rect 7896 9818 7902 9820
rect 7958 9818 7982 9820
rect 8038 9818 8062 9820
rect 8118 9818 8142 9820
rect 8198 9818 8204 9820
rect 7958 9766 7960 9818
rect 8140 9766 8142 9818
rect 7896 9764 7902 9766
rect 7958 9764 7982 9766
rect 8038 9764 8062 9766
rect 8118 9764 8142 9766
rect 8198 9764 8204 9766
rect 7896 9755 8204 9764
rect 7896 8732 8204 8741
rect 7896 8730 7902 8732
rect 7958 8730 7982 8732
rect 8038 8730 8062 8732
rect 8118 8730 8142 8732
rect 8198 8730 8204 8732
rect 7958 8678 7960 8730
rect 8140 8678 8142 8730
rect 7896 8676 7902 8678
rect 7958 8676 7982 8678
rect 8038 8676 8062 8678
rect 8118 8676 8142 8678
rect 8198 8676 8204 8678
rect 7896 8667 8204 8676
rect 7896 7644 8204 7653
rect 7896 7642 7902 7644
rect 7958 7642 7982 7644
rect 8038 7642 8062 7644
rect 8118 7642 8142 7644
rect 8198 7642 8204 7644
rect 7958 7590 7960 7642
rect 8140 7590 8142 7642
rect 7896 7588 7902 7590
rect 7958 7588 7982 7590
rect 8038 7588 8062 7590
rect 8118 7588 8142 7590
rect 8198 7588 8204 7590
rect 7896 7579 8204 7588
rect 7748 6928 7800 6934
rect 7748 6870 7800 6876
rect 5356 6792 5408 6798
rect 5356 6734 5408 6740
rect 5540 6792 5592 6798
rect 5540 6734 5592 6740
rect 4988 4684 5040 4690
rect 4988 4626 5040 4632
rect 5552 4622 5580 6734
rect 7896 6556 8204 6565
rect 7896 6554 7902 6556
rect 7958 6554 7982 6556
rect 8038 6554 8062 6556
rect 8118 6554 8142 6556
rect 8198 6554 8204 6556
rect 7958 6502 7960 6554
rect 8140 6502 8142 6554
rect 7896 6500 7902 6502
rect 7958 6500 7982 6502
rect 8038 6500 8062 6502
rect 8118 6500 8142 6502
rect 8198 6500 8204 6502
rect 7896 6491 8204 6500
rect 7896 5468 8204 5477
rect 7896 5466 7902 5468
rect 7958 5466 7982 5468
rect 8038 5466 8062 5468
rect 8118 5466 8142 5468
rect 8198 5466 8204 5468
rect 7958 5414 7960 5466
rect 8140 5414 8142 5466
rect 7896 5412 7902 5414
rect 7958 5412 7982 5414
rect 8038 5412 8062 5414
rect 8118 5412 8142 5414
rect 8198 5412 8204 5414
rect 7896 5403 8204 5412
rect 5724 4684 5776 4690
rect 5724 4626 5776 4632
rect 4896 4616 4948 4622
rect 4896 4558 4948 4564
rect 5540 4616 5592 4622
rect 5540 4558 5592 4564
rect 4908 4078 4936 4558
rect 4896 4072 4948 4078
rect 4896 4014 4948 4020
rect 5264 3460 5316 3466
rect 5264 3402 5316 3408
rect 4804 2848 4856 2854
rect 4804 2790 4856 2796
rect 4423 2748 4731 2757
rect 4423 2746 4429 2748
rect 4485 2746 4509 2748
rect 4565 2746 4589 2748
rect 4645 2746 4669 2748
rect 4725 2746 4731 2748
rect 4485 2694 4487 2746
rect 4667 2694 4669 2746
rect 4423 2692 4429 2694
rect 4485 2692 4509 2694
rect 4565 2692 4589 2694
rect 4645 2692 4669 2694
rect 4725 2692 4731 2694
rect 4423 2683 4731 2692
rect 5276 2650 5304 3402
rect 5264 2644 5316 2650
rect 5264 2586 5316 2592
rect 5736 2446 5764 4626
rect 6736 4480 6788 4486
rect 6736 4422 6788 4428
rect 6552 3936 6604 3942
rect 6552 3878 6604 3884
rect 5816 3596 5868 3602
rect 5816 3538 5868 3544
rect 5724 2440 5776 2446
rect 5724 2382 5776 2388
rect 4356 1006 4568 1034
rect 4540 800 4568 1006
rect 5828 800 5856 3538
rect 6564 3058 6592 3878
rect 6552 3052 6604 3058
rect 6552 2994 6604 3000
rect 6748 2990 6776 4422
rect 7896 4380 8204 4389
rect 7896 4378 7902 4380
rect 7958 4378 7982 4380
rect 8038 4378 8062 4380
rect 8118 4378 8142 4380
rect 8198 4378 8204 4380
rect 7958 4326 7960 4378
rect 8140 4326 8142 4378
rect 7896 4324 7902 4326
rect 7958 4324 7982 4326
rect 8038 4324 8062 4326
rect 8118 4324 8142 4326
rect 8198 4324 8204 4326
rect 7896 4315 8204 4324
rect 7748 4072 7800 4078
rect 7748 4014 7800 4020
rect 8392 4072 8444 4078
rect 8392 4014 8444 4020
rect 7656 4004 7708 4010
rect 7656 3946 7708 3952
rect 6736 2984 6788 2990
rect 6736 2926 6788 2932
rect 6460 2916 6512 2922
rect 6460 2858 6512 2864
rect 6472 800 6500 2858
rect 7668 2650 7696 3946
rect 7760 3738 7788 4014
rect 7748 3732 7800 3738
rect 7748 3674 7800 3680
rect 7896 3292 8204 3301
rect 7896 3290 7902 3292
rect 7958 3290 7982 3292
rect 8038 3290 8062 3292
rect 8118 3290 8142 3292
rect 8198 3290 8204 3292
rect 7958 3238 7960 3290
rect 8140 3238 8142 3290
rect 7896 3236 7902 3238
rect 7958 3236 7982 3238
rect 8038 3236 8062 3238
rect 8118 3236 8142 3238
rect 8198 3236 8204 3238
rect 7896 3227 8204 3236
rect 7656 2644 7708 2650
rect 7656 2586 7708 2592
rect 7896 2204 8204 2213
rect 7896 2202 7902 2204
rect 7958 2202 7982 2204
rect 8038 2202 8062 2204
rect 8118 2202 8142 2204
rect 8198 2202 8204 2204
rect 7958 2150 7960 2202
rect 8140 2150 8142 2202
rect 7896 2148 7902 2150
rect 7958 2148 7982 2150
rect 8038 2148 8062 2150
rect 8118 2148 8142 2150
rect 8198 2148 8204 2150
rect 7896 2139 8204 2148
rect 8404 800 8432 4014
rect 8944 3528 8996 3534
rect 8944 3470 8996 3476
rect 8956 3058 8984 3470
rect 9128 3392 9180 3398
rect 9128 3334 9180 3340
rect 9140 3126 9168 3334
rect 9128 3120 9180 3126
rect 9128 3062 9180 3068
rect 8944 3052 8996 3058
rect 8944 2994 8996 3000
rect 9416 2514 9444 24006
rect 9968 3534 9996 30602
rect 10704 15502 10732 36518
rect 11369 36476 11677 36485
rect 11369 36474 11375 36476
rect 11431 36474 11455 36476
rect 11511 36474 11535 36476
rect 11591 36474 11615 36476
rect 11671 36474 11677 36476
rect 11431 36422 11433 36474
rect 11613 36422 11615 36474
rect 11369 36420 11375 36422
rect 11431 36420 11455 36422
rect 11511 36420 11535 36422
rect 11591 36420 11615 36422
rect 11671 36420 11677 36422
rect 11369 36411 11677 36420
rect 14476 36106 14504 45902
rect 14842 45724 15150 45733
rect 14842 45722 14848 45724
rect 14904 45722 14928 45724
rect 14984 45722 15008 45724
rect 15064 45722 15088 45724
rect 15144 45722 15150 45724
rect 14904 45670 14906 45722
rect 15086 45670 15088 45722
rect 14842 45668 14848 45670
rect 14904 45668 14928 45670
rect 14984 45668 15008 45670
rect 15064 45668 15088 45670
rect 15144 45668 15150 45670
rect 14842 45659 15150 45668
rect 19444 45490 19472 45902
rect 19616 45892 19668 45898
rect 19616 45834 19668 45840
rect 22284 45892 22336 45898
rect 22284 45834 22336 45840
rect 19628 45626 19656 45834
rect 21788 45724 22096 45733
rect 21788 45722 21794 45724
rect 21850 45722 21874 45724
rect 21930 45722 21954 45724
rect 22010 45722 22034 45724
rect 22090 45722 22096 45724
rect 21850 45670 21852 45722
rect 22032 45670 22034 45722
rect 21788 45668 21794 45670
rect 21850 45668 21874 45670
rect 21930 45668 21954 45670
rect 22010 45668 22034 45670
rect 22090 45668 22096 45670
rect 21788 45659 22096 45668
rect 22296 45626 22324 45834
rect 19616 45620 19668 45626
rect 19616 45562 19668 45568
rect 22284 45620 22336 45626
rect 22284 45562 22336 45568
rect 22388 45490 22416 46446
rect 19340 45484 19392 45490
rect 19340 45426 19392 45432
rect 19432 45484 19484 45490
rect 19432 45426 19484 45432
rect 20628 45484 20680 45490
rect 20628 45426 20680 45432
rect 22376 45484 22428 45490
rect 22376 45426 22428 45432
rect 18315 45180 18623 45189
rect 18315 45178 18321 45180
rect 18377 45178 18401 45180
rect 18457 45178 18481 45180
rect 18537 45178 18561 45180
rect 18617 45178 18623 45180
rect 18377 45126 18379 45178
rect 18559 45126 18561 45178
rect 18315 45124 18321 45126
rect 18377 45124 18401 45126
rect 18457 45124 18481 45126
rect 18537 45124 18561 45126
rect 18617 45124 18623 45126
rect 18315 45115 18623 45124
rect 14842 44636 15150 44645
rect 14842 44634 14848 44636
rect 14904 44634 14928 44636
rect 14984 44634 15008 44636
rect 15064 44634 15088 44636
rect 15144 44634 15150 44636
rect 14904 44582 14906 44634
rect 15086 44582 15088 44634
rect 14842 44580 14848 44582
rect 14904 44580 14928 44582
rect 14984 44580 15008 44582
rect 15064 44580 15088 44582
rect 15144 44580 15150 44582
rect 14842 44571 15150 44580
rect 18315 44092 18623 44101
rect 18315 44090 18321 44092
rect 18377 44090 18401 44092
rect 18457 44090 18481 44092
rect 18537 44090 18561 44092
rect 18617 44090 18623 44092
rect 18377 44038 18379 44090
rect 18559 44038 18561 44090
rect 18315 44036 18321 44038
rect 18377 44036 18401 44038
rect 18457 44036 18481 44038
rect 18537 44036 18561 44038
rect 18617 44036 18623 44038
rect 18315 44027 18623 44036
rect 14842 43548 15150 43557
rect 14842 43546 14848 43548
rect 14904 43546 14928 43548
rect 14984 43546 15008 43548
rect 15064 43546 15088 43548
rect 15144 43546 15150 43548
rect 14904 43494 14906 43546
rect 15086 43494 15088 43546
rect 14842 43492 14848 43494
rect 14904 43492 14928 43494
rect 14984 43492 15008 43494
rect 15064 43492 15088 43494
rect 15144 43492 15150 43494
rect 14842 43483 15150 43492
rect 18315 43004 18623 43013
rect 18315 43002 18321 43004
rect 18377 43002 18401 43004
rect 18457 43002 18481 43004
rect 18537 43002 18561 43004
rect 18617 43002 18623 43004
rect 18377 42950 18379 43002
rect 18559 42950 18561 43002
rect 18315 42948 18321 42950
rect 18377 42948 18401 42950
rect 18457 42948 18481 42950
rect 18537 42948 18561 42950
rect 18617 42948 18623 42950
rect 18315 42939 18623 42948
rect 14842 42460 15150 42469
rect 14842 42458 14848 42460
rect 14904 42458 14928 42460
rect 14984 42458 15008 42460
rect 15064 42458 15088 42460
rect 15144 42458 15150 42460
rect 14904 42406 14906 42458
rect 15086 42406 15088 42458
rect 14842 42404 14848 42406
rect 14904 42404 14928 42406
rect 14984 42404 15008 42406
rect 15064 42404 15088 42406
rect 15144 42404 15150 42406
rect 14842 42395 15150 42404
rect 18315 41916 18623 41925
rect 18315 41914 18321 41916
rect 18377 41914 18401 41916
rect 18457 41914 18481 41916
rect 18537 41914 18561 41916
rect 18617 41914 18623 41916
rect 18377 41862 18379 41914
rect 18559 41862 18561 41914
rect 18315 41860 18321 41862
rect 18377 41860 18401 41862
rect 18457 41860 18481 41862
rect 18537 41860 18561 41862
rect 18617 41860 18623 41862
rect 18315 41851 18623 41860
rect 19352 41414 19380 45426
rect 20640 45354 20668 45426
rect 20628 45348 20680 45354
rect 20628 45290 20680 45296
rect 19352 41386 19472 41414
rect 14842 41372 15150 41381
rect 14842 41370 14848 41372
rect 14904 41370 14928 41372
rect 14984 41370 15008 41372
rect 15064 41370 15088 41372
rect 15144 41370 15150 41372
rect 14904 41318 14906 41370
rect 15086 41318 15088 41370
rect 14842 41316 14848 41318
rect 14904 41316 14928 41318
rect 14984 41316 15008 41318
rect 15064 41316 15088 41318
rect 15144 41316 15150 41318
rect 14842 41307 15150 41316
rect 18315 40828 18623 40837
rect 18315 40826 18321 40828
rect 18377 40826 18401 40828
rect 18457 40826 18481 40828
rect 18537 40826 18561 40828
rect 18617 40826 18623 40828
rect 18377 40774 18379 40826
rect 18559 40774 18561 40826
rect 18315 40772 18321 40774
rect 18377 40772 18401 40774
rect 18457 40772 18481 40774
rect 18537 40772 18561 40774
rect 18617 40772 18623 40774
rect 18315 40763 18623 40772
rect 14842 40284 15150 40293
rect 14842 40282 14848 40284
rect 14904 40282 14928 40284
rect 14984 40282 15008 40284
rect 15064 40282 15088 40284
rect 15144 40282 15150 40284
rect 14904 40230 14906 40282
rect 15086 40230 15088 40282
rect 14842 40228 14848 40230
rect 14904 40228 14928 40230
rect 14984 40228 15008 40230
rect 15064 40228 15088 40230
rect 15144 40228 15150 40230
rect 14842 40219 15150 40228
rect 18315 39740 18623 39749
rect 18315 39738 18321 39740
rect 18377 39738 18401 39740
rect 18457 39738 18481 39740
rect 18537 39738 18561 39740
rect 18617 39738 18623 39740
rect 18377 39686 18379 39738
rect 18559 39686 18561 39738
rect 18315 39684 18321 39686
rect 18377 39684 18401 39686
rect 18457 39684 18481 39686
rect 18537 39684 18561 39686
rect 18617 39684 18623 39686
rect 18315 39675 18623 39684
rect 14842 39196 15150 39205
rect 14842 39194 14848 39196
rect 14904 39194 14928 39196
rect 14984 39194 15008 39196
rect 15064 39194 15088 39196
rect 15144 39194 15150 39196
rect 14904 39142 14906 39194
rect 15086 39142 15088 39194
rect 14842 39140 14848 39142
rect 14904 39140 14928 39142
rect 14984 39140 15008 39142
rect 15064 39140 15088 39142
rect 15144 39140 15150 39142
rect 14842 39131 15150 39140
rect 18972 38956 19024 38962
rect 18972 38898 19024 38904
rect 18315 38652 18623 38661
rect 18315 38650 18321 38652
rect 18377 38650 18401 38652
rect 18457 38650 18481 38652
rect 18537 38650 18561 38652
rect 18617 38650 18623 38652
rect 18377 38598 18379 38650
rect 18559 38598 18561 38650
rect 18315 38596 18321 38598
rect 18377 38596 18401 38598
rect 18457 38596 18481 38598
rect 18537 38596 18561 38598
rect 18617 38596 18623 38598
rect 18315 38587 18623 38596
rect 18984 38554 19012 38898
rect 18696 38548 18748 38554
rect 18696 38490 18748 38496
rect 18972 38548 19024 38554
rect 18972 38490 19024 38496
rect 18052 38276 18104 38282
rect 18052 38218 18104 38224
rect 14842 38108 15150 38117
rect 14842 38106 14848 38108
rect 14904 38106 14928 38108
rect 14984 38106 15008 38108
rect 15064 38106 15088 38108
rect 15144 38106 15150 38108
rect 14904 38054 14906 38106
rect 15086 38054 15088 38106
rect 14842 38052 14848 38054
rect 14904 38052 14928 38054
rect 14984 38052 15008 38054
rect 15064 38052 15088 38054
rect 15144 38052 15150 38054
rect 14842 38043 15150 38052
rect 16856 37324 16908 37330
rect 16856 37266 16908 37272
rect 15292 37188 15344 37194
rect 15292 37130 15344 37136
rect 14842 37020 15150 37029
rect 14842 37018 14848 37020
rect 14904 37018 14928 37020
rect 14984 37018 15008 37020
rect 15064 37018 15088 37020
rect 15144 37018 15150 37020
rect 14904 36966 14906 37018
rect 15086 36966 15088 37018
rect 14842 36964 14848 36966
rect 14904 36964 14928 36966
rect 14984 36964 15008 36966
rect 15064 36964 15088 36966
rect 15144 36964 15150 36966
rect 14842 36955 15150 36964
rect 14464 36100 14516 36106
rect 14464 36042 14516 36048
rect 14842 35932 15150 35941
rect 14842 35930 14848 35932
rect 14904 35930 14928 35932
rect 14984 35930 15008 35932
rect 15064 35930 15088 35932
rect 15144 35930 15150 35932
rect 14904 35878 14906 35930
rect 15086 35878 15088 35930
rect 14842 35876 14848 35878
rect 14904 35876 14928 35878
rect 14984 35876 15008 35878
rect 15064 35876 15088 35878
rect 15144 35876 15150 35878
rect 14842 35867 15150 35876
rect 11369 35388 11677 35397
rect 11369 35386 11375 35388
rect 11431 35386 11455 35388
rect 11511 35386 11535 35388
rect 11591 35386 11615 35388
rect 11671 35386 11677 35388
rect 11431 35334 11433 35386
rect 11613 35334 11615 35386
rect 11369 35332 11375 35334
rect 11431 35332 11455 35334
rect 11511 35332 11535 35334
rect 11591 35332 11615 35334
rect 11671 35332 11677 35334
rect 11369 35323 11677 35332
rect 14842 34844 15150 34853
rect 14842 34842 14848 34844
rect 14904 34842 14928 34844
rect 14984 34842 15008 34844
rect 15064 34842 15088 34844
rect 15144 34842 15150 34844
rect 14904 34790 14906 34842
rect 15086 34790 15088 34842
rect 14842 34788 14848 34790
rect 14904 34788 14928 34790
rect 14984 34788 15008 34790
rect 15064 34788 15088 34790
rect 15144 34788 15150 34790
rect 14842 34779 15150 34788
rect 14740 34672 14792 34678
rect 14740 34614 14792 34620
rect 11369 34300 11677 34309
rect 11369 34298 11375 34300
rect 11431 34298 11455 34300
rect 11511 34298 11535 34300
rect 11591 34298 11615 34300
rect 11671 34298 11677 34300
rect 11431 34246 11433 34298
rect 11613 34246 11615 34298
rect 11369 34244 11375 34246
rect 11431 34244 11455 34246
rect 11511 34244 11535 34246
rect 11591 34244 11615 34246
rect 11671 34244 11677 34246
rect 11369 34235 11677 34244
rect 11369 33212 11677 33221
rect 11369 33210 11375 33212
rect 11431 33210 11455 33212
rect 11511 33210 11535 33212
rect 11591 33210 11615 33212
rect 11671 33210 11677 33212
rect 11431 33158 11433 33210
rect 11613 33158 11615 33210
rect 11369 33156 11375 33158
rect 11431 33156 11455 33158
rect 11511 33156 11535 33158
rect 11591 33156 11615 33158
rect 11671 33156 11677 33158
rect 11369 33147 11677 33156
rect 11369 32124 11677 32133
rect 11369 32122 11375 32124
rect 11431 32122 11455 32124
rect 11511 32122 11535 32124
rect 11591 32122 11615 32124
rect 11671 32122 11677 32124
rect 11431 32070 11433 32122
rect 11613 32070 11615 32122
rect 11369 32068 11375 32070
rect 11431 32068 11455 32070
rect 11511 32068 11535 32070
rect 11591 32068 11615 32070
rect 11671 32068 11677 32070
rect 11369 32059 11677 32068
rect 11369 31036 11677 31045
rect 11369 31034 11375 31036
rect 11431 31034 11455 31036
rect 11511 31034 11535 31036
rect 11591 31034 11615 31036
rect 11671 31034 11677 31036
rect 11431 30982 11433 31034
rect 11613 30982 11615 31034
rect 11369 30980 11375 30982
rect 11431 30980 11455 30982
rect 11511 30980 11535 30982
rect 11591 30980 11615 30982
rect 11671 30980 11677 30982
rect 11369 30971 11677 30980
rect 12624 30728 12676 30734
rect 12624 30670 12676 30676
rect 11369 29948 11677 29957
rect 11369 29946 11375 29948
rect 11431 29946 11455 29948
rect 11511 29946 11535 29948
rect 11591 29946 11615 29948
rect 11671 29946 11677 29948
rect 11431 29894 11433 29946
rect 11613 29894 11615 29946
rect 11369 29892 11375 29894
rect 11431 29892 11455 29894
rect 11511 29892 11535 29894
rect 11591 29892 11615 29894
rect 11671 29892 11677 29894
rect 11369 29883 11677 29892
rect 11369 28860 11677 28869
rect 11369 28858 11375 28860
rect 11431 28858 11455 28860
rect 11511 28858 11535 28860
rect 11591 28858 11615 28860
rect 11671 28858 11677 28860
rect 11431 28806 11433 28858
rect 11613 28806 11615 28858
rect 11369 28804 11375 28806
rect 11431 28804 11455 28806
rect 11511 28804 11535 28806
rect 11591 28804 11615 28806
rect 11671 28804 11677 28806
rect 11369 28795 11677 28804
rect 11369 27772 11677 27781
rect 11369 27770 11375 27772
rect 11431 27770 11455 27772
rect 11511 27770 11535 27772
rect 11591 27770 11615 27772
rect 11671 27770 11677 27772
rect 11431 27718 11433 27770
rect 11613 27718 11615 27770
rect 11369 27716 11375 27718
rect 11431 27716 11455 27718
rect 11511 27716 11535 27718
rect 11591 27716 11615 27718
rect 11671 27716 11677 27718
rect 11369 27707 11677 27716
rect 11369 26684 11677 26693
rect 11369 26682 11375 26684
rect 11431 26682 11455 26684
rect 11511 26682 11535 26684
rect 11591 26682 11615 26684
rect 11671 26682 11677 26684
rect 11431 26630 11433 26682
rect 11613 26630 11615 26682
rect 11369 26628 11375 26630
rect 11431 26628 11455 26630
rect 11511 26628 11535 26630
rect 11591 26628 11615 26630
rect 11671 26628 11677 26630
rect 11369 26619 11677 26628
rect 11369 25596 11677 25605
rect 11369 25594 11375 25596
rect 11431 25594 11455 25596
rect 11511 25594 11535 25596
rect 11591 25594 11615 25596
rect 11671 25594 11677 25596
rect 11431 25542 11433 25594
rect 11613 25542 11615 25594
rect 11369 25540 11375 25542
rect 11431 25540 11455 25542
rect 11511 25540 11535 25542
rect 11591 25540 11615 25542
rect 11671 25540 11677 25542
rect 11369 25531 11677 25540
rect 11369 24508 11677 24517
rect 11369 24506 11375 24508
rect 11431 24506 11455 24508
rect 11511 24506 11535 24508
rect 11591 24506 11615 24508
rect 11671 24506 11677 24508
rect 11431 24454 11433 24506
rect 11613 24454 11615 24506
rect 11369 24452 11375 24454
rect 11431 24452 11455 24454
rect 11511 24452 11535 24454
rect 11591 24452 11615 24454
rect 11671 24452 11677 24454
rect 11369 24443 11677 24452
rect 11369 23420 11677 23429
rect 11369 23418 11375 23420
rect 11431 23418 11455 23420
rect 11511 23418 11535 23420
rect 11591 23418 11615 23420
rect 11671 23418 11677 23420
rect 11431 23366 11433 23418
rect 11613 23366 11615 23418
rect 11369 23364 11375 23366
rect 11431 23364 11455 23366
rect 11511 23364 11535 23366
rect 11591 23364 11615 23366
rect 11671 23364 11677 23366
rect 11369 23355 11677 23364
rect 11369 22332 11677 22341
rect 11369 22330 11375 22332
rect 11431 22330 11455 22332
rect 11511 22330 11535 22332
rect 11591 22330 11615 22332
rect 11671 22330 11677 22332
rect 11431 22278 11433 22330
rect 11613 22278 11615 22330
rect 11369 22276 11375 22278
rect 11431 22276 11455 22278
rect 11511 22276 11535 22278
rect 11591 22276 11615 22278
rect 11671 22276 11677 22278
rect 11369 22267 11677 22276
rect 11369 21244 11677 21253
rect 11369 21242 11375 21244
rect 11431 21242 11455 21244
rect 11511 21242 11535 21244
rect 11591 21242 11615 21244
rect 11671 21242 11677 21244
rect 11431 21190 11433 21242
rect 11613 21190 11615 21242
rect 11369 21188 11375 21190
rect 11431 21188 11455 21190
rect 11511 21188 11535 21190
rect 11591 21188 11615 21190
rect 11671 21188 11677 21190
rect 11369 21179 11677 21188
rect 12636 20602 12664 30670
rect 14752 21146 14780 34614
rect 14842 33756 15150 33765
rect 14842 33754 14848 33756
rect 14904 33754 14928 33756
rect 14984 33754 15008 33756
rect 15064 33754 15088 33756
rect 15144 33754 15150 33756
rect 14904 33702 14906 33754
rect 15086 33702 15088 33754
rect 14842 33700 14848 33702
rect 14904 33700 14928 33702
rect 14984 33700 15008 33702
rect 15064 33700 15088 33702
rect 15144 33700 15150 33702
rect 14842 33691 15150 33700
rect 15304 32910 15332 37130
rect 15752 36916 15804 36922
rect 15752 36858 15804 36864
rect 15660 36236 15712 36242
rect 15660 36178 15712 36184
rect 15292 32904 15344 32910
rect 15292 32846 15344 32852
rect 14842 32668 15150 32677
rect 14842 32666 14848 32668
rect 14904 32666 14928 32668
rect 14984 32666 15008 32668
rect 15064 32666 15088 32668
rect 15144 32666 15150 32668
rect 14904 32614 14906 32666
rect 15086 32614 15088 32666
rect 14842 32612 14848 32614
rect 14904 32612 14928 32614
rect 14984 32612 15008 32614
rect 15064 32612 15088 32614
rect 15144 32612 15150 32614
rect 14842 32603 15150 32612
rect 15304 32502 15332 32846
rect 15476 32768 15528 32774
rect 15476 32710 15528 32716
rect 15488 32570 15516 32710
rect 15476 32564 15528 32570
rect 15476 32506 15528 32512
rect 15292 32496 15344 32502
rect 15292 32438 15344 32444
rect 15304 31822 15332 32438
rect 15292 31816 15344 31822
rect 15292 31758 15344 31764
rect 15672 31754 15700 36178
rect 15764 32502 15792 36858
rect 16672 36712 16724 36718
rect 16672 36654 16724 36660
rect 16580 36168 16632 36174
rect 16580 36110 16632 36116
rect 16488 36032 16540 36038
rect 16488 35974 16540 35980
rect 16500 35698 16528 35974
rect 16592 35766 16620 36110
rect 16580 35760 16632 35766
rect 16580 35702 16632 35708
rect 16488 35692 16540 35698
rect 16488 35634 16540 35640
rect 16684 35630 16712 36654
rect 16868 36242 16896 37266
rect 18064 37194 18092 38218
rect 18708 37874 18736 38490
rect 18696 37868 18748 37874
rect 18696 37810 18748 37816
rect 19064 37868 19116 37874
rect 19064 37810 19116 37816
rect 18236 37664 18288 37670
rect 18236 37606 18288 37612
rect 18248 37466 18276 37606
rect 18315 37564 18623 37573
rect 18315 37562 18321 37564
rect 18377 37562 18401 37564
rect 18457 37562 18481 37564
rect 18537 37562 18561 37564
rect 18617 37562 18623 37564
rect 18377 37510 18379 37562
rect 18559 37510 18561 37562
rect 18315 37508 18321 37510
rect 18377 37508 18401 37510
rect 18457 37508 18481 37510
rect 18537 37508 18561 37510
rect 18617 37508 18623 37510
rect 18315 37499 18623 37508
rect 18236 37460 18288 37466
rect 18236 37402 18288 37408
rect 19076 37398 19104 37810
rect 19340 37460 19392 37466
rect 19340 37402 19392 37408
rect 19064 37392 19116 37398
rect 19064 37334 19116 37340
rect 17960 37188 18012 37194
rect 17960 37130 18012 37136
rect 18052 37188 18104 37194
rect 18052 37130 18104 37136
rect 17408 37120 17460 37126
rect 17408 37062 17460 37068
rect 17420 36786 17448 37062
rect 17408 36780 17460 36786
rect 17408 36722 17460 36728
rect 17776 36576 17828 36582
rect 17776 36518 17828 36524
rect 16856 36236 16908 36242
rect 16856 36178 16908 36184
rect 17788 36174 17816 36518
rect 17776 36168 17828 36174
rect 17776 36110 17828 36116
rect 17132 36032 17184 36038
rect 17132 35974 17184 35980
rect 17592 36032 17644 36038
rect 17592 35974 17644 35980
rect 17144 35766 17172 35974
rect 17132 35760 17184 35766
rect 17132 35702 17184 35708
rect 16672 35624 16724 35630
rect 16672 35566 16724 35572
rect 16856 35624 16908 35630
rect 16856 35566 16908 35572
rect 16684 34542 16712 35566
rect 16868 35086 16896 35566
rect 16856 35080 16908 35086
rect 16856 35022 16908 35028
rect 16672 34536 16724 34542
rect 16672 34478 16724 34484
rect 16764 33380 16816 33386
rect 16764 33322 16816 33328
rect 16776 33046 16804 33322
rect 16764 33040 16816 33046
rect 16764 32982 16816 32988
rect 16212 32972 16264 32978
rect 16212 32914 16264 32920
rect 15936 32836 15988 32842
rect 15936 32778 15988 32784
rect 15752 32496 15804 32502
rect 15752 32438 15804 32444
rect 15580 31726 15700 31754
rect 14842 31580 15150 31589
rect 14842 31578 14848 31580
rect 14904 31578 14928 31580
rect 14984 31578 15008 31580
rect 15064 31578 15088 31580
rect 15144 31578 15150 31580
rect 14904 31526 14906 31578
rect 15086 31526 15088 31578
rect 14842 31524 14848 31526
rect 14904 31524 14928 31526
rect 14984 31524 15008 31526
rect 15064 31524 15088 31526
rect 15144 31524 15150 31526
rect 14842 31515 15150 31524
rect 14842 30492 15150 30501
rect 14842 30490 14848 30492
rect 14904 30490 14928 30492
rect 14984 30490 15008 30492
rect 15064 30490 15088 30492
rect 15144 30490 15150 30492
rect 14904 30438 14906 30490
rect 15086 30438 15088 30490
rect 14842 30436 14848 30438
rect 14904 30436 14928 30438
rect 14984 30436 15008 30438
rect 15064 30436 15088 30438
rect 15144 30436 15150 30438
rect 14842 30427 15150 30436
rect 14842 29404 15150 29413
rect 14842 29402 14848 29404
rect 14904 29402 14928 29404
rect 14984 29402 15008 29404
rect 15064 29402 15088 29404
rect 15144 29402 15150 29404
rect 14904 29350 14906 29402
rect 15086 29350 15088 29402
rect 14842 29348 14848 29350
rect 14904 29348 14928 29350
rect 14984 29348 15008 29350
rect 15064 29348 15088 29350
rect 15144 29348 15150 29350
rect 14842 29339 15150 29348
rect 14842 28316 15150 28325
rect 14842 28314 14848 28316
rect 14904 28314 14928 28316
rect 14984 28314 15008 28316
rect 15064 28314 15088 28316
rect 15144 28314 15150 28316
rect 14904 28262 14906 28314
rect 15086 28262 15088 28314
rect 14842 28260 14848 28262
rect 14904 28260 14928 28262
rect 14984 28260 15008 28262
rect 15064 28260 15088 28262
rect 15144 28260 15150 28262
rect 14842 28251 15150 28260
rect 15384 27532 15436 27538
rect 15384 27474 15436 27480
rect 14842 27228 15150 27237
rect 14842 27226 14848 27228
rect 14904 27226 14928 27228
rect 14984 27226 15008 27228
rect 15064 27226 15088 27228
rect 15144 27226 15150 27228
rect 14904 27174 14906 27226
rect 15086 27174 15088 27226
rect 14842 27172 14848 27174
rect 14904 27172 14928 27174
rect 14984 27172 15008 27174
rect 15064 27172 15088 27174
rect 15144 27172 15150 27174
rect 14842 27163 15150 27172
rect 14842 26140 15150 26149
rect 14842 26138 14848 26140
rect 14904 26138 14928 26140
rect 14984 26138 15008 26140
rect 15064 26138 15088 26140
rect 15144 26138 15150 26140
rect 14904 26086 14906 26138
rect 15086 26086 15088 26138
rect 14842 26084 14848 26086
rect 14904 26084 14928 26086
rect 14984 26084 15008 26086
rect 15064 26084 15088 26086
rect 15144 26084 15150 26086
rect 14842 26075 15150 26084
rect 14842 25052 15150 25061
rect 14842 25050 14848 25052
rect 14904 25050 14928 25052
rect 14984 25050 15008 25052
rect 15064 25050 15088 25052
rect 15144 25050 15150 25052
rect 14904 24998 14906 25050
rect 15086 24998 15088 25050
rect 14842 24996 14848 24998
rect 14904 24996 14928 24998
rect 14984 24996 15008 24998
rect 15064 24996 15088 24998
rect 15144 24996 15150 24998
rect 14842 24987 15150 24996
rect 14842 23964 15150 23973
rect 14842 23962 14848 23964
rect 14904 23962 14928 23964
rect 14984 23962 15008 23964
rect 15064 23962 15088 23964
rect 15144 23962 15150 23964
rect 14904 23910 14906 23962
rect 15086 23910 15088 23962
rect 14842 23908 14848 23910
rect 14904 23908 14928 23910
rect 14984 23908 15008 23910
rect 15064 23908 15088 23910
rect 15144 23908 15150 23910
rect 14842 23899 15150 23908
rect 14842 22876 15150 22885
rect 14842 22874 14848 22876
rect 14904 22874 14928 22876
rect 14984 22874 15008 22876
rect 15064 22874 15088 22876
rect 15144 22874 15150 22876
rect 14904 22822 14906 22874
rect 15086 22822 15088 22874
rect 14842 22820 14848 22822
rect 14904 22820 14928 22822
rect 14984 22820 15008 22822
rect 15064 22820 15088 22822
rect 15144 22820 15150 22822
rect 14842 22811 15150 22820
rect 15396 22574 15424 27474
rect 15580 25838 15608 31726
rect 15764 30682 15792 32438
rect 15948 32366 15976 32778
rect 16224 32570 16252 32914
rect 16764 32904 16816 32910
rect 16764 32846 16816 32852
rect 16580 32768 16632 32774
rect 16580 32710 16632 32716
rect 16212 32564 16264 32570
rect 16212 32506 16264 32512
rect 15936 32360 15988 32366
rect 15936 32302 15988 32308
rect 15844 32224 15896 32230
rect 15844 32166 15896 32172
rect 15856 31346 15884 32166
rect 15948 32026 15976 32302
rect 15936 32020 15988 32026
rect 15936 31962 15988 31968
rect 16592 31890 16620 32710
rect 16580 31884 16632 31890
rect 16580 31826 16632 31832
rect 16028 31680 16080 31686
rect 16028 31622 16080 31628
rect 15844 31340 15896 31346
rect 15844 31282 15896 31288
rect 15936 31136 15988 31142
rect 15936 31078 15988 31084
rect 15764 30666 15884 30682
rect 15948 30666 15976 31078
rect 16040 30938 16068 31622
rect 16592 31346 16620 31826
rect 16580 31340 16632 31346
rect 16580 31282 16632 31288
rect 16028 30932 16080 30938
rect 16028 30874 16080 30880
rect 15764 30660 15896 30666
rect 15764 30654 15844 30660
rect 15844 30602 15896 30608
rect 15936 30660 15988 30666
rect 15936 30602 15988 30608
rect 15752 29504 15804 29510
rect 15752 29446 15804 29452
rect 15764 28558 15792 29446
rect 15856 28762 15884 30602
rect 16040 29730 16068 30874
rect 16212 30592 16264 30598
rect 16212 30534 16264 30540
rect 16224 30258 16252 30534
rect 16212 30252 16264 30258
rect 16212 30194 16264 30200
rect 16776 29850 16804 32846
rect 16868 31890 16896 35022
rect 17604 35018 17632 35974
rect 17592 35012 17644 35018
rect 17592 34954 17644 34960
rect 17972 34950 18000 37130
rect 18064 36922 18092 37130
rect 18420 37120 18472 37126
rect 18420 37062 18472 37068
rect 18052 36916 18104 36922
rect 18052 36858 18104 36864
rect 18432 36786 18460 37062
rect 18420 36780 18472 36786
rect 18420 36722 18472 36728
rect 18788 36576 18840 36582
rect 18788 36518 18840 36524
rect 18315 36476 18623 36485
rect 18315 36474 18321 36476
rect 18377 36474 18401 36476
rect 18457 36474 18481 36476
rect 18537 36474 18561 36476
rect 18617 36474 18623 36476
rect 18377 36422 18379 36474
rect 18559 36422 18561 36474
rect 18315 36420 18321 36422
rect 18377 36420 18401 36422
rect 18457 36420 18481 36422
rect 18537 36420 18561 36422
rect 18617 36420 18623 36422
rect 18315 36411 18623 36420
rect 18236 36100 18288 36106
rect 18236 36042 18288 36048
rect 18144 36032 18196 36038
rect 18144 35974 18196 35980
rect 17960 34944 18012 34950
rect 17960 34886 18012 34892
rect 18156 33522 18184 35974
rect 18248 35562 18276 36042
rect 18800 35698 18828 36518
rect 19352 36038 19380 37402
rect 19444 36854 19472 41386
rect 20076 38956 20128 38962
rect 20076 38898 20128 38904
rect 20088 38826 20116 38898
rect 20536 38888 20588 38894
rect 20536 38830 20588 38836
rect 19708 38820 19760 38826
rect 19708 38762 19760 38768
rect 20076 38820 20128 38826
rect 20076 38762 20128 38768
rect 19616 38752 19668 38758
rect 19616 38694 19668 38700
rect 19522 38448 19578 38457
rect 19522 38383 19578 38392
rect 19536 37330 19564 38383
rect 19628 38282 19656 38694
rect 19616 38276 19668 38282
rect 19616 38218 19668 38224
rect 19616 37936 19668 37942
rect 19616 37878 19668 37884
rect 19628 37466 19656 37878
rect 19616 37460 19668 37466
rect 19616 37402 19668 37408
rect 19524 37324 19576 37330
rect 19524 37266 19576 37272
rect 19432 36848 19484 36854
rect 19432 36790 19484 36796
rect 19340 36032 19392 36038
rect 19340 35974 19392 35980
rect 18788 35692 18840 35698
rect 18788 35634 18840 35640
rect 18236 35556 18288 35562
rect 18236 35498 18288 35504
rect 17960 33516 18012 33522
rect 17960 33458 18012 33464
rect 18144 33516 18196 33522
rect 18144 33458 18196 33464
rect 17972 33114 18000 33458
rect 18248 33402 18276 35498
rect 18315 35388 18623 35397
rect 18315 35386 18321 35388
rect 18377 35386 18401 35388
rect 18457 35386 18481 35388
rect 18537 35386 18561 35388
rect 18617 35386 18623 35388
rect 18377 35334 18379 35386
rect 18559 35334 18561 35386
rect 18315 35332 18321 35334
rect 18377 35332 18401 35334
rect 18457 35332 18481 35334
rect 18537 35332 18561 35334
rect 18617 35332 18623 35334
rect 18315 35323 18623 35332
rect 18880 34944 18932 34950
rect 18880 34886 18932 34892
rect 18315 34300 18623 34309
rect 18315 34298 18321 34300
rect 18377 34298 18401 34300
rect 18457 34298 18481 34300
rect 18537 34298 18561 34300
rect 18617 34298 18623 34300
rect 18377 34246 18379 34298
rect 18559 34246 18561 34298
rect 18315 34244 18321 34246
rect 18377 34244 18401 34246
rect 18457 34244 18481 34246
rect 18537 34244 18561 34246
rect 18617 34244 18623 34246
rect 18315 34235 18623 34244
rect 18696 33584 18748 33590
rect 18696 33526 18748 33532
rect 18064 33374 18276 33402
rect 17868 33108 17920 33114
rect 17868 33050 17920 33056
rect 17960 33108 18012 33114
rect 17960 33050 18012 33056
rect 17880 32994 17908 33050
rect 17880 32966 18000 32994
rect 17040 32224 17092 32230
rect 17040 32166 17092 32172
rect 16856 31884 16908 31890
rect 16856 31826 16908 31832
rect 16868 30258 16896 31826
rect 17052 31822 17080 32166
rect 17040 31816 17092 31822
rect 17040 31758 17092 31764
rect 17972 31754 18000 32966
rect 18064 32910 18092 33374
rect 18144 33312 18196 33318
rect 18144 33254 18196 33260
rect 18052 32904 18104 32910
rect 18052 32846 18104 32852
rect 18052 32768 18104 32774
rect 18052 32710 18104 32716
rect 18064 32434 18092 32710
rect 18156 32434 18184 33254
rect 18315 33212 18623 33221
rect 18315 33210 18321 33212
rect 18377 33210 18401 33212
rect 18457 33210 18481 33212
rect 18537 33210 18561 33212
rect 18617 33210 18623 33212
rect 18377 33158 18379 33210
rect 18559 33158 18561 33210
rect 18315 33156 18321 33158
rect 18377 33156 18401 33158
rect 18457 33156 18481 33158
rect 18537 33156 18561 33158
rect 18617 33156 18623 33158
rect 18315 33147 18623 33156
rect 18236 33108 18288 33114
rect 18236 33050 18288 33056
rect 18248 32892 18276 33050
rect 18708 32978 18736 33526
rect 18892 33522 18920 34886
rect 19352 34746 19380 35974
rect 19616 35488 19668 35494
rect 19616 35430 19668 35436
rect 19340 34740 19392 34746
rect 19340 34682 19392 34688
rect 19628 34610 19656 35430
rect 19720 35018 19748 38762
rect 20088 38486 20116 38762
rect 20352 38752 20404 38758
rect 20352 38694 20404 38700
rect 20076 38480 20128 38486
rect 20076 38422 20128 38428
rect 19984 37868 20036 37874
rect 19984 37810 20036 37816
rect 19996 37262 20024 37810
rect 20088 37670 20116 38422
rect 20076 37664 20128 37670
rect 20076 37606 20128 37612
rect 19984 37256 20036 37262
rect 19984 37198 20036 37204
rect 20364 36174 20392 38694
rect 20444 38208 20496 38214
rect 20444 38150 20496 38156
rect 20456 37466 20484 38150
rect 20548 37738 20576 38830
rect 20640 38457 20668 45290
rect 22480 45082 22508 47058
rect 22572 46034 22600 49200
rect 23216 47122 23244 49200
rect 23204 47116 23256 47122
rect 23204 47058 23256 47064
rect 23020 46980 23072 46986
rect 23020 46922 23072 46928
rect 22560 46028 22612 46034
rect 22560 45970 22612 45976
rect 23032 45558 23060 46922
rect 23860 45966 23888 49200
rect 26606 49056 26662 49065
rect 26606 48991 26662 49000
rect 25261 47356 25569 47365
rect 25261 47354 25267 47356
rect 25323 47354 25347 47356
rect 25403 47354 25427 47356
rect 25483 47354 25507 47356
rect 25563 47354 25569 47356
rect 25323 47302 25325 47354
rect 25505 47302 25507 47354
rect 25261 47300 25267 47302
rect 25323 47300 25347 47302
rect 25403 47300 25427 47302
rect 25483 47300 25507 47302
rect 25563 47300 25569 47302
rect 25261 47291 25569 47300
rect 26620 47122 26648 48991
rect 26608 47116 26660 47122
rect 26608 47058 26660 47064
rect 24768 47048 24820 47054
rect 24768 46990 24820 46996
rect 26146 47016 26202 47025
rect 24308 46504 24360 46510
rect 24308 46446 24360 46452
rect 23848 45960 23900 45966
rect 23848 45902 23900 45908
rect 23572 45824 23624 45830
rect 23572 45766 23624 45772
rect 23020 45552 23072 45558
rect 23020 45494 23072 45500
rect 23112 45484 23164 45490
rect 23112 45426 23164 45432
rect 22468 45076 22520 45082
rect 22468 45018 22520 45024
rect 23124 45014 23152 45426
rect 23112 45008 23164 45014
rect 23112 44950 23164 44956
rect 21788 44636 22096 44645
rect 21788 44634 21794 44636
rect 21850 44634 21874 44636
rect 21930 44634 21954 44636
rect 22010 44634 22034 44636
rect 22090 44634 22096 44636
rect 21850 44582 21852 44634
rect 22032 44582 22034 44634
rect 21788 44580 21794 44582
rect 21850 44580 21874 44582
rect 21930 44580 21954 44582
rect 22010 44580 22034 44582
rect 22090 44580 22096 44582
rect 21788 44571 22096 44580
rect 21788 43548 22096 43557
rect 21788 43546 21794 43548
rect 21850 43546 21874 43548
rect 21930 43546 21954 43548
rect 22010 43546 22034 43548
rect 22090 43546 22096 43548
rect 21850 43494 21852 43546
rect 22032 43494 22034 43546
rect 21788 43492 21794 43494
rect 21850 43492 21874 43494
rect 21930 43492 21954 43494
rect 22010 43492 22034 43494
rect 22090 43492 22096 43494
rect 21788 43483 22096 43492
rect 21788 42460 22096 42469
rect 21788 42458 21794 42460
rect 21850 42458 21874 42460
rect 21930 42458 21954 42460
rect 22010 42458 22034 42460
rect 22090 42458 22096 42460
rect 21850 42406 21852 42458
rect 22032 42406 22034 42458
rect 21788 42404 21794 42406
rect 21850 42404 21874 42406
rect 21930 42404 21954 42406
rect 22010 42404 22034 42406
rect 22090 42404 22096 42406
rect 21788 42395 22096 42404
rect 21788 41372 22096 41381
rect 21788 41370 21794 41372
rect 21850 41370 21874 41372
rect 21930 41370 21954 41372
rect 22010 41370 22034 41372
rect 22090 41370 22096 41372
rect 21850 41318 21852 41370
rect 22032 41318 22034 41370
rect 21788 41316 21794 41318
rect 21850 41316 21874 41318
rect 21930 41316 21954 41318
rect 22010 41316 22034 41318
rect 22090 41316 22096 41318
rect 21788 41307 22096 41316
rect 21788 40284 22096 40293
rect 21788 40282 21794 40284
rect 21850 40282 21874 40284
rect 21930 40282 21954 40284
rect 22010 40282 22034 40284
rect 22090 40282 22096 40284
rect 21850 40230 21852 40282
rect 22032 40230 22034 40282
rect 21788 40228 21794 40230
rect 21850 40228 21874 40230
rect 21930 40228 21954 40230
rect 22010 40228 22034 40230
rect 22090 40228 22096 40230
rect 21788 40219 22096 40228
rect 21788 39196 22096 39205
rect 21788 39194 21794 39196
rect 21850 39194 21874 39196
rect 21930 39194 21954 39196
rect 22010 39194 22034 39196
rect 22090 39194 22096 39196
rect 21850 39142 21852 39194
rect 22032 39142 22034 39194
rect 21788 39140 21794 39142
rect 21850 39140 21874 39142
rect 21930 39140 21954 39142
rect 22010 39140 22034 39142
rect 22090 39140 22096 39142
rect 21788 39131 22096 39140
rect 20720 38956 20772 38962
rect 20720 38898 20772 38904
rect 20732 38554 20760 38898
rect 21640 38888 21692 38894
rect 21640 38830 21692 38836
rect 21272 38752 21324 38758
rect 21272 38694 21324 38700
rect 20720 38548 20772 38554
rect 20720 38490 20772 38496
rect 20626 38448 20682 38457
rect 20626 38383 20682 38392
rect 21284 38282 21312 38694
rect 21652 38282 21680 38830
rect 21824 38820 21876 38826
rect 21824 38762 21876 38768
rect 21836 38350 21864 38762
rect 21824 38344 21876 38350
rect 21824 38286 21876 38292
rect 21272 38276 21324 38282
rect 21272 38218 21324 38224
rect 21640 38276 21692 38282
rect 21640 38218 21692 38224
rect 21364 38208 21416 38214
rect 21364 38150 21416 38156
rect 20720 38004 20772 38010
rect 20720 37946 20772 37952
rect 20812 38004 20864 38010
rect 20812 37946 20864 37952
rect 20732 37738 20760 37946
rect 20536 37732 20588 37738
rect 20536 37674 20588 37680
rect 20720 37732 20772 37738
rect 20720 37674 20772 37680
rect 20444 37460 20496 37466
rect 20444 37402 20496 37408
rect 20076 36168 20128 36174
rect 20076 36110 20128 36116
rect 20352 36168 20404 36174
rect 20352 36110 20404 36116
rect 20088 35766 20116 36110
rect 20076 35760 20128 35766
rect 20076 35702 20128 35708
rect 20088 35086 20116 35702
rect 20548 35290 20576 37674
rect 20732 37262 20760 37674
rect 20824 37398 20852 37946
rect 20996 37936 21048 37942
rect 20996 37878 21048 37884
rect 20812 37392 20864 37398
rect 20812 37334 20864 37340
rect 20720 37256 20772 37262
rect 20720 37198 20772 37204
rect 20732 36378 20760 37198
rect 20824 37126 20852 37334
rect 21008 37262 21036 37878
rect 21376 37874 21404 38150
rect 21364 37868 21416 37874
rect 21364 37810 21416 37816
rect 21652 37806 21680 38218
rect 21788 38108 22096 38117
rect 21788 38106 21794 38108
rect 21850 38106 21874 38108
rect 21930 38106 21954 38108
rect 22010 38106 22034 38108
rect 22090 38106 22096 38108
rect 21850 38054 21852 38106
rect 22032 38054 22034 38106
rect 21788 38052 21794 38054
rect 21850 38052 21874 38054
rect 21930 38052 21954 38054
rect 22010 38052 22034 38054
rect 22090 38052 22096 38054
rect 21788 38043 22096 38052
rect 21640 37800 21692 37806
rect 21640 37742 21692 37748
rect 21364 37324 21416 37330
rect 21364 37266 21416 37272
rect 20996 37256 21048 37262
rect 20996 37198 21048 37204
rect 20812 37120 20864 37126
rect 20812 37062 20864 37068
rect 20824 36582 20852 37062
rect 20812 36576 20864 36582
rect 20812 36518 20864 36524
rect 20720 36372 20772 36378
rect 20720 36314 20772 36320
rect 20732 35894 20760 36314
rect 20732 35866 20852 35894
rect 20536 35284 20588 35290
rect 20536 35226 20588 35232
rect 20076 35080 20128 35086
rect 20076 35022 20128 35028
rect 19708 35012 19760 35018
rect 19708 34954 19760 34960
rect 19616 34604 19668 34610
rect 19616 34546 19668 34552
rect 19432 33584 19484 33590
rect 19432 33526 19484 33532
rect 18880 33516 18932 33522
rect 18880 33458 18932 33464
rect 18788 33040 18840 33046
rect 18788 32982 18840 32988
rect 18696 32972 18748 32978
rect 18696 32914 18748 32920
rect 18328 32904 18380 32910
rect 18248 32864 18328 32892
rect 18052 32428 18104 32434
rect 18052 32370 18104 32376
rect 18144 32428 18196 32434
rect 18144 32370 18196 32376
rect 18248 32026 18276 32864
rect 18328 32846 18380 32852
rect 18708 32366 18736 32914
rect 18800 32366 18828 32982
rect 18696 32360 18748 32366
rect 18696 32302 18748 32308
rect 18788 32360 18840 32366
rect 18788 32302 18840 32308
rect 18315 32124 18623 32133
rect 18315 32122 18321 32124
rect 18377 32122 18401 32124
rect 18457 32122 18481 32124
rect 18537 32122 18561 32124
rect 18617 32122 18623 32124
rect 18377 32070 18379 32122
rect 18559 32070 18561 32122
rect 18315 32068 18321 32070
rect 18377 32068 18401 32070
rect 18457 32068 18481 32070
rect 18537 32068 18561 32070
rect 18617 32068 18623 32070
rect 18315 32059 18623 32068
rect 18236 32020 18288 32026
rect 18236 31962 18288 31968
rect 17972 31726 18092 31754
rect 17868 31340 17920 31346
rect 17868 31282 17920 31288
rect 17880 30938 17908 31282
rect 17868 30932 17920 30938
rect 17868 30874 17920 30880
rect 17960 30728 18012 30734
rect 17960 30670 18012 30676
rect 17972 30394 18000 30670
rect 17960 30388 18012 30394
rect 17960 30330 18012 30336
rect 16856 30252 16908 30258
rect 16856 30194 16908 30200
rect 16764 29844 16816 29850
rect 16764 29786 16816 29792
rect 15948 29702 16068 29730
rect 16672 29708 16724 29714
rect 15948 29646 15976 29702
rect 16672 29650 16724 29656
rect 15936 29640 15988 29646
rect 15936 29582 15988 29588
rect 16580 29640 16632 29646
rect 16580 29582 16632 29588
rect 15948 29170 15976 29582
rect 15936 29164 15988 29170
rect 15936 29106 15988 29112
rect 15936 28960 15988 28966
rect 15936 28902 15988 28908
rect 15844 28756 15896 28762
rect 15844 28698 15896 28704
rect 15752 28552 15804 28558
rect 15752 28494 15804 28500
rect 15660 27328 15712 27334
rect 15660 27270 15712 27276
rect 15672 27062 15700 27270
rect 15660 27056 15712 27062
rect 15660 26998 15712 27004
rect 15568 25832 15620 25838
rect 15568 25774 15620 25780
rect 15580 24274 15608 25774
rect 15568 24268 15620 24274
rect 15568 24210 15620 24216
rect 15384 22568 15436 22574
rect 15384 22510 15436 22516
rect 15580 22094 15608 24210
rect 15764 22094 15792 28494
rect 15948 28490 15976 28902
rect 16592 28762 16620 29582
rect 16684 29170 16712 29650
rect 16764 29504 16816 29510
rect 16764 29446 16816 29452
rect 16672 29164 16724 29170
rect 16672 29106 16724 29112
rect 16580 28756 16632 28762
rect 16580 28698 16632 28704
rect 16672 28688 16724 28694
rect 16672 28630 16724 28636
rect 15936 28484 15988 28490
rect 15936 28426 15988 28432
rect 16212 27056 16264 27062
rect 16212 26998 16264 27004
rect 15844 25832 15896 25838
rect 15844 25774 15896 25780
rect 15856 24954 15884 25774
rect 16120 25696 16172 25702
rect 16120 25638 16172 25644
rect 16132 25294 16160 25638
rect 16120 25288 16172 25294
rect 16120 25230 16172 25236
rect 15844 24948 15896 24954
rect 15844 24890 15896 24896
rect 16120 22432 16172 22438
rect 16120 22374 16172 22380
rect 15580 22066 15700 22094
rect 15764 22066 15884 22094
rect 14842 21788 15150 21797
rect 14842 21786 14848 21788
rect 14904 21786 14928 21788
rect 14984 21786 15008 21788
rect 15064 21786 15088 21788
rect 15144 21786 15150 21788
rect 14904 21734 14906 21786
rect 15086 21734 15088 21786
rect 14842 21732 14848 21734
rect 14904 21732 14928 21734
rect 14984 21732 15008 21734
rect 15064 21732 15088 21734
rect 15144 21732 15150 21734
rect 14842 21723 15150 21732
rect 15200 21548 15252 21554
rect 15200 21490 15252 21496
rect 14740 21140 14792 21146
rect 14740 21082 14792 21088
rect 14740 20868 14792 20874
rect 14740 20810 14792 20816
rect 12624 20596 12676 20602
rect 12624 20538 12676 20544
rect 14464 20528 14516 20534
rect 14464 20470 14516 20476
rect 14752 20482 14780 20810
rect 14842 20700 15150 20709
rect 14842 20698 14848 20700
rect 14904 20698 14928 20700
rect 14984 20698 15008 20700
rect 15064 20698 15088 20700
rect 15144 20698 15150 20700
rect 14904 20646 14906 20698
rect 15086 20646 15088 20698
rect 14842 20644 14848 20646
rect 14904 20644 14928 20646
rect 14984 20644 15008 20646
rect 15064 20644 15088 20646
rect 15144 20644 15150 20646
rect 14842 20635 15150 20644
rect 12992 20460 13044 20466
rect 12992 20402 13044 20408
rect 13084 20460 13136 20466
rect 13084 20402 13136 20408
rect 11369 20156 11677 20165
rect 11369 20154 11375 20156
rect 11431 20154 11455 20156
rect 11511 20154 11535 20156
rect 11591 20154 11615 20156
rect 11671 20154 11677 20156
rect 11431 20102 11433 20154
rect 11613 20102 11615 20154
rect 11369 20100 11375 20102
rect 11431 20100 11455 20102
rect 11511 20100 11535 20102
rect 11591 20100 11615 20102
rect 11671 20100 11677 20102
rect 11369 20091 11677 20100
rect 12808 19440 12860 19446
rect 12808 19382 12860 19388
rect 11369 19068 11677 19077
rect 11369 19066 11375 19068
rect 11431 19066 11455 19068
rect 11511 19066 11535 19068
rect 11591 19066 11615 19068
rect 11671 19066 11677 19068
rect 11431 19014 11433 19066
rect 11613 19014 11615 19066
rect 11369 19012 11375 19014
rect 11431 19012 11455 19014
rect 11511 19012 11535 19014
rect 11591 19012 11615 19014
rect 11671 19012 11677 19014
rect 11369 19003 11677 19012
rect 12820 18766 12848 19382
rect 13004 18970 13032 20402
rect 13096 20058 13124 20402
rect 13820 20392 13872 20398
rect 13820 20334 13872 20340
rect 13084 20052 13136 20058
rect 13084 19994 13136 20000
rect 13728 19848 13780 19854
rect 13728 19790 13780 19796
rect 13740 19378 13768 19790
rect 13832 19514 13860 20334
rect 14004 19780 14056 19786
rect 14004 19722 14056 19728
rect 13820 19508 13872 19514
rect 13820 19450 13872 19456
rect 14016 19378 14044 19722
rect 14280 19712 14332 19718
rect 14280 19654 14332 19660
rect 14096 19508 14148 19514
rect 14096 19450 14148 19456
rect 13728 19372 13780 19378
rect 13728 19314 13780 19320
rect 14004 19372 14056 19378
rect 14004 19314 14056 19320
rect 12992 18964 13044 18970
rect 12992 18906 13044 18912
rect 13740 18766 13768 19314
rect 14016 19242 14044 19314
rect 14004 19236 14056 19242
rect 14004 19178 14056 19184
rect 13820 18964 13872 18970
rect 13820 18906 13872 18912
rect 12256 18760 12308 18766
rect 12256 18702 12308 18708
rect 12808 18760 12860 18766
rect 12808 18702 12860 18708
rect 13728 18760 13780 18766
rect 13728 18702 13780 18708
rect 12268 18290 12296 18702
rect 12256 18284 12308 18290
rect 12820 18272 12848 18702
rect 13452 18624 13504 18630
rect 13452 18566 13504 18572
rect 13464 18290 13492 18566
rect 12900 18284 12952 18290
rect 12820 18244 12900 18272
rect 12256 18226 12308 18232
rect 12900 18226 12952 18232
rect 13452 18284 13504 18290
rect 13452 18226 13504 18232
rect 11888 18216 11940 18222
rect 11888 18158 11940 18164
rect 11369 17980 11677 17989
rect 11369 17978 11375 17980
rect 11431 17978 11455 17980
rect 11511 17978 11535 17980
rect 11591 17978 11615 17980
rect 11671 17978 11677 17980
rect 11431 17926 11433 17978
rect 11613 17926 11615 17978
rect 11369 17924 11375 17926
rect 11431 17924 11455 17926
rect 11511 17924 11535 17926
rect 11591 17924 11615 17926
rect 11671 17924 11677 17926
rect 11369 17915 11677 17924
rect 11369 16892 11677 16901
rect 11369 16890 11375 16892
rect 11431 16890 11455 16892
rect 11511 16890 11535 16892
rect 11591 16890 11615 16892
rect 11671 16890 11677 16892
rect 11431 16838 11433 16890
rect 11613 16838 11615 16890
rect 11369 16836 11375 16838
rect 11431 16836 11455 16838
rect 11511 16836 11535 16838
rect 11591 16836 11615 16838
rect 11671 16836 11677 16838
rect 11369 16827 11677 16836
rect 11369 15804 11677 15813
rect 11369 15802 11375 15804
rect 11431 15802 11455 15804
rect 11511 15802 11535 15804
rect 11591 15802 11615 15804
rect 11671 15802 11677 15804
rect 11431 15750 11433 15802
rect 11613 15750 11615 15802
rect 11369 15748 11375 15750
rect 11431 15748 11455 15750
rect 11511 15748 11535 15750
rect 11591 15748 11615 15750
rect 11671 15748 11677 15750
rect 11369 15739 11677 15748
rect 10692 15496 10744 15502
rect 10692 15438 10744 15444
rect 11060 15428 11112 15434
rect 11060 15370 11112 15376
rect 11072 12442 11100 15370
rect 11369 14716 11677 14725
rect 11369 14714 11375 14716
rect 11431 14714 11455 14716
rect 11511 14714 11535 14716
rect 11591 14714 11615 14716
rect 11671 14714 11677 14716
rect 11431 14662 11433 14714
rect 11613 14662 11615 14714
rect 11369 14660 11375 14662
rect 11431 14660 11455 14662
rect 11511 14660 11535 14662
rect 11591 14660 11615 14662
rect 11671 14660 11677 14662
rect 11369 14651 11677 14660
rect 11369 13628 11677 13637
rect 11369 13626 11375 13628
rect 11431 13626 11455 13628
rect 11511 13626 11535 13628
rect 11591 13626 11615 13628
rect 11671 13626 11677 13628
rect 11431 13574 11433 13626
rect 11613 13574 11615 13626
rect 11369 13572 11375 13574
rect 11431 13572 11455 13574
rect 11511 13572 11535 13574
rect 11591 13572 11615 13574
rect 11671 13572 11677 13574
rect 11369 13563 11677 13572
rect 11369 12540 11677 12549
rect 11369 12538 11375 12540
rect 11431 12538 11455 12540
rect 11511 12538 11535 12540
rect 11591 12538 11615 12540
rect 11671 12538 11677 12540
rect 11431 12486 11433 12538
rect 11613 12486 11615 12538
rect 11369 12484 11375 12486
rect 11431 12484 11455 12486
rect 11511 12484 11535 12486
rect 11591 12484 11615 12486
rect 11671 12484 11677 12486
rect 11369 12475 11677 12484
rect 11060 12436 11112 12442
rect 11060 12378 11112 12384
rect 11369 11452 11677 11461
rect 11369 11450 11375 11452
rect 11431 11450 11455 11452
rect 11511 11450 11535 11452
rect 11591 11450 11615 11452
rect 11671 11450 11677 11452
rect 11431 11398 11433 11450
rect 11613 11398 11615 11450
rect 11369 11396 11375 11398
rect 11431 11396 11455 11398
rect 11511 11396 11535 11398
rect 11591 11396 11615 11398
rect 11671 11396 11677 11398
rect 11369 11387 11677 11396
rect 11369 10364 11677 10373
rect 11369 10362 11375 10364
rect 11431 10362 11455 10364
rect 11511 10362 11535 10364
rect 11591 10362 11615 10364
rect 11671 10362 11677 10364
rect 11431 10310 11433 10362
rect 11613 10310 11615 10362
rect 11369 10308 11375 10310
rect 11431 10308 11455 10310
rect 11511 10308 11535 10310
rect 11591 10308 11615 10310
rect 11671 10308 11677 10310
rect 11369 10299 11677 10308
rect 11369 9276 11677 9285
rect 11369 9274 11375 9276
rect 11431 9274 11455 9276
rect 11511 9274 11535 9276
rect 11591 9274 11615 9276
rect 11671 9274 11677 9276
rect 11431 9222 11433 9274
rect 11613 9222 11615 9274
rect 11369 9220 11375 9222
rect 11431 9220 11455 9222
rect 11511 9220 11535 9222
rect 11591 9220 11615 9222
rect 11671 9220 11677 9222
rect 11369 9211 11677 9220
rect 11369 8188 11677 8197
rect 11369 8186 11375 8188
rect 11431 8186 11455 8188
rect 11511 8186 11535 8188
rect 11591 8186 11615 8188
rect 11671 8186 11677 8188
rect 11431 8134 11433 8186
rect 11613 8134 11615 8186
rect 11369 8132 11375 8134
rect 11431 8132 11455 8134
rect 11511 8132 11535 8134
rect 11591 8132 11615 8134
rect 11671 8132 11677 8134
rect 11369 8123 11677 8132
rect 11369 7100 11677 7109
rect 11369 7098 11375 7100
rect 11431 7098 11455 7100
rect 11511 7098 11535 7100
rect 11591 7098 11615 7100
rect 11671 7098 11677 7100
rect 11431 7046 11433 7098
rect 11613 7046 11615 7098
rect 11369 7044 11375 7046
rect 11431 7044 11455 7046
rect 11511 7044 11535 7046
rect 11591 7044 11615 7046
rect 11671 7044 11677 7046
rect 11369 7035 11677 7044
rect 11369 6012 11677 6021
rect 11369 6010 11375 6012
rect 11431 6010 11455 6012
rect 11511 6010 11535 6012
rect 11591 6010 11615 6012
rect 11671 6010 11677 6012
rect 11431 5958 11433 6010
rect 11613 5958 11615 6010
rect 11369 5956 11375 5958
rect 11431 5956 11455 5958
rect 11511 5956 11535 5958
rect 11591 5956 11615 5958
rect 11671 5956 11677 5958
rect 11369 5947 11677 5956
rect 11369 4924 11677 4933
rect 11369 4922 11375 4924
rect 11431 4922 11455 4924
rect 11511 4922 11535 4924
rect 11591 4922 11615 4924
rect 11671 4922 11677 4924
rect 11431 4870 11433 4922
rect 11613 4870 11615 4922
rect 11369 4868 11375 4870
rect 11431 4868 11455 4870
rect 11511 4868 11535 4870
rect 11591 4868 11615 4870
rect 11671 4868 11677 4870
rect 11369 4859 11677 4868
rect 11369 3836 11677 3845
rect 11369 3834 11375 3836
rect 11431 3834 11455 3836
rect 11511 3834 11535 3836
rect 11591 3834 11615 3836
rect 11671 3834 11677 3836
rect 11431 3782 11433 3834
rect 11613 3782 11615 3834
rect 11369 3780 11375 3782
rect 11431 3780 11455 3782
rect 11511 3780 11535 3782
rect 11591 3780 11615 3782
rect 11671 3780 11677 3782
rect 11369 3771 11677 3780
rect 11900 3602 11928 18158
rect 13452 18080 13504 18086
rect 13452 18022 13504 18028
rect 11980 16244 12032 16250
rect 11980 16186 12032 16192
rect 11992 15434 12020 16186
rect 13464 15570 13492 18022
rect 13740 17678 13768 18702
rect 13832 18290 13860 18906
rect 14004 18692 14056 18698
rect 14004 18634 14056 18640
rect 14016 18290 14044 18634
rect 14108 18290 14136 19450
rect 14292 19310 14320 19654
rect 14476 19514 14504 20470
rect 14752 20466 14872 20482
rect 14648 20460 14700 20466
rect 14752 20460 14884 20466
rect 14752 20454 14832 20460
rect 14648 20402 14700 20408
rect 14832 20402 14884 20408
rect 14660 20058 14688 20402
rect 14648 20052 14700 20058
rect 14648 19994 14700 20000
rect 14740 20052 14792 20058
rect 14740 19994 14792 20000
rect 14556 19848 14608 19854
rect 14556 19790 14608 19796
rect 14648 19848 14700 19854
rect 14648 19790 14700 19796
rect 14464 19508 14516 19514
rect 14464 19450 14516 19456
rect 14280 19304 14332 19310
rect 14280 19246 14332 19252
rect 14292 18698 14320 19246
rect 14280 18692 14332 18698
rect 14280 18634 14332 18640
rect 14476 18358 14504 19450
rect 14568 19446 14596 19790
rect 14556 19440 14608 19446
rect 14556 19382 14608 19388
rect 14556 19168 14608 19174
rect 14556 19110 14608 19116
rect 14568 18834 14596 19110
rect 14556 18828 14608 18834
rect 14556 18770 14608 18776
rect 14464 18352 14516 18358
rect 14464 18294 14516 18300
rect 14568 18290 14596 18770
rect 14660 18630 14688 19790
rect 14752 19718 14780 19994
rect 14740 19712 14792 19718
rect 14740 19654 14792 19660
rect 14752 19514 14780 19654
rect 14842 19612 15150 19621
rect 14842 19610 14848 19612
rect 14904 19610 14928 19612
rect 14984 19610 15008 19612
rect 15064 19610 15088 19612
rect 15144 19610 15150 19612
rect 14904 19558 14906 19610
rect 15086 19558 15088 19610
rect 14842 19556 14848 19558
rect 14904 19556 14928 19558
rect 14984 19556 15008 19558
rect 15064 19556 15088 19558
rect 15144 19556 15150 19558
rect 14842 19547 15150 19556
rect 14740 19508 14792 19514
rect 14740 19450 14792 19456
rect 14740 19236 14792 19242
rect 14740 19178 14792 19184
rect 14752 18698 14780 19178
rect 14740 18692 14792 18698
rect 14740 18634 14792 18640
rect 14648 18624 14700 18630
rect 14648 18566 14700 18572
rect 13820 18284 13872 18290
rect 13820 18226 13872 18232
rect 14004 18284 14056 18290
rect 14004 18226 14056 18232
rect 14096 18284 14148 18290
rect 14096 18226 14148 18232
rect 14556 18284 14608 18290
rect 14556 18226 14608 18232
rect 13832 17678 13860 18226
rect 13728 17672 13780 17678
rect 13728 17614 13780 17620
rect 13820 17672 13872 17678
rect 13820 17614 13872 17620
rect 14016 17270 14044 18226
rect 14556 18080 14608 18086
rect 14556 18022 14608 18028
rect 14004 17264 14056 17270
rect 14004 17206 14056 17212
rect 14568 17202 14596 18022
rect 14660 17814 14688 18566
rect 14752 18290 14780 18634
rect 14842 18524 15150 18533
rect 14842 18522 14848 18524
rect 14904 18522 14928 18524
rect 14984 18522 15008 18524
rect 15064 18522 15088 18524
rect 15144 18522 15150 18524
rect 14904 18470 14906 18522
rect 15086 18470 15088 18522
rect 14842 18468 14848 18470
rect 14904 18468 14928 18470
rect 14984 18468 15008 18470
rect 15064 18468 15088 18470
rect 15144 18468 15150 18470
rect 14842 18459 15150 18468
rect 14740 18284 14792 18290
rect 14740 18226 14792 18232
rect 14752 17814 14780 18226
rect 15212 18154 15240 21490
rect 15672 21486 15700 22066
rect 15660 21480 15712 21486
rect 15660 21422 15712 21428
rect 15384 20868 15436 20874
rect 15384 20810 15436 20816
rect 15396 20058 15424 20810
rect 15384 20052 15436 20058
rect 15384 19994 15436 20000
rect 15660 18760 15712 18766
rect 15660 18702 15712 18708
rect 15200 18148 15252 18154
rect 15200 18090 15252 18096
rect 14648 17808 14700 17814
rect 14648 17750 14700 17756
rect 14740 17808 14792 17814
rect 14740 17750 14792 17756
rect 14740 17672 14792 17678
rect 14740 17614 14792 17620
rect 14556 17196 14608 17202
rect 14556 17138 14608 17144
rect 14752 17066 14780 17614
rect 14842 17436 15150 17445
rect 14842 17434 14848 17436
rect 14904 17434 14928 17436
rect 14984 17434 15008 17436
rect 15064 17434 15088 17436
rect 15144 17434 15150 17436
rect 14904 17382 14906 17434
rect 15086 17382 15088 17434
rect 14842 17380 14848 17382
rect 14904 17380 14928 17382
rect 14984 17380 15008 17382
rect 15064 17380 15088 17382
rect 15144 17380 15150 17382
rect 14842 17371 15150 17380
rect 14556 17060 14608 17066
rect 14556 17002 14608 17008
rect 14740 17060 14792 17066
rect 14740 17002 14792 17008
rect 13452 15564 13504 15570
rect 13452 15506 13504 15512
rect 11980 15428 12032 15434
rect 11980 15370 12032 15376
rect 11992 4146 12020 15370
rect 12992 5024 13044 5030
rect 12992 4966 13044 4972
rect 12808 4616 12860 4622
rect 12808 4558 12860 4564
rect 12820 4146 12848 4558
rect 13004 4214 13032 4966
rect 12992 4208 13044 4214
rect 12992 4150 13044 4156
rect 11980 4140 12032 4146
rect 11980 4082 12032 4088
rect 12808 4140 12860 4146
rect 12808 4082 12860 4088
rect 13544 4072 13596 4078
rect 13544 4014 13596 4020
rect 12072 3936 12124 3942
rect 12072 3878 12124 3884
rect 12084 3602 12112 3878
rect 11888 3596 11940 3602
rect 11888 3538 11940 3544
rect 12072 3596 12124 3602
rect 12072 3538 12124 3544
rect 12440 3596 12492 3602
rect 12440 3538 12492 3544
rect 9956 3528 10008 3534
rect 9956 3470 10008 3476
rect 10600 3528 10652 3534
rect 10600 3470 10652 3476
rect 11704 3528 11756 3534
rect 11704 3470 11756 3476
rect 9968 3194 9996 3470
rect 9956 3188 10008 3194
rect 9956 3130 10008 3136
rect 9680 2984 9732 2990
rect 9680 2926 9732 2932
rect 9404 2508 9456 2514
rect 9404 2450 9456 2456
rect 9036 2440 9088 2446
rect 9036 2382 9088 2388
rect 9048 800 9076 2382
rect 9692 800 9720 2926
rect 10612 2106 10640 3470
rect 11716 3058 11744 3470
rect 11888 3392 11940 3398
rect 11888 3334 11940 3340
rect 11900 3126 11928 3334
rect 11888 3120 11940 3126
rect 11888 3062 11940 3068
rect 11704 3052 11756 3058
rect 11704 2994 11756 3000
rect 10968 2984 11020 2990
rect 10968 2926 11020 2932
rect 10600 2100 10652 2106
rect 10600 2042 10652 2048
rect 10980 800 11008 2926
rect 11369 2748 11677 2757
rect 11369 2746 11375 2748
rect 11431 2746 11455 2748
rect 11511 2746 11535 2748
rect 11591 2746 11615 2748
rect 11671 2746 11677 2748
rect 11431 2694 11433 2746
rect 11613 2694 11615 2746
rect 11369 2692 11375 2694
rect 11431 2692 11455 2694
rect 11511 2692 11535 2694
rect 11591 2692 11615 2694
rect 11671 2692 11677 2694
rect 11369 2683 11677 2692
rect 12452 2310 12480 3538
rect 12440 2304 12492 2310
rect 12440 2246 12492 2252
rect 13556 800 13584 4014
rect 14568 4010 14596 17002
rect 15672 16794 15700 18702
rect 15752 18284 15804 18290
rect 15752 18226 15804 18232
rect 15764 17338 15792 18226
rect 15856 17678 15884 22066
rect 16132 22030 16160 22374
rect 16120 22024 16172 22030
rect 16120 21966 16172 21972
rect 16224 21962 16252 26998
rect 16684 26518 16712 28630
rect 16776 28558 16804 29446
rect 16868 29102 16896 30194
rect 18064 29714 18092 31726
rect 18248 31482 18276 31962
rect 18328 31680 18380 31686
rect 18328 31622 18380 31628
rect 18236 31476 18288 31482
rect 18236 31418 18288 31424
rect 18340 31346 18368 31622
rect 18328 31340 18380 31346
rect 18328 31282 18380 31288
rect 18315 31036 18623 31045
rect 18315 31034 18321 31036
rect 18377 31034 18401 31036
rect 18457 31034 18481 31036
rect 18537 31034 18561 31036
rect 18617 31034 18623 31036
rect 18377 30982 18379 31034
rect 18559 30982 18561 31034
rect 18315 30980 18321 30982
rect 18377 30980 18401 30982
rect 18457 30980 18481 30982
rect 18537 30980 18561 30982
rect 18617 30980 18623 30982
rect 18315 30971 18623 30980
rect 18315 29948 18623 29957
rect 18315 29946 18321 29948
rect 18377 29946 18401 29948
rect 18457 29946 18481 29948
rect 18537 29946 18561 29948
rect 18617 29946 18623 29948
rect 18377 29894 18379 29946
rect 18559 29894 18561 29946
rect 18315 29892 18321 29894
rect 18377 29892 18401 29894
rect 18457 29892 18481 29894
rect 18537 29892 18561 29894
rect 18617 29892 18623 29894
rect 18315 29883 18623 29892
rect 18800 29850 18828 32302
rect 18892 31822 18920 33458
rect 18972 33380 19024 33386
rect 18972 33322 19024 33328
rect 18984 32842 19012 33322
rect 19340 33312 19392 33318
rect 19340 33254 19392 33260
rect 18972 32836 19024 32842
rect 18972 32778 19024 32784
rect 19156 32836 19208 32842
rect 19156 32778 19208 32784
rect 18880 31816 18932 31822
rect 18880 31758 18932 31764
rect 18236 29844 18288 29850
rect 18236 29786 18288 29792
rect 18788 29844 18840 29850
rect 18788 29786 18840 29792
rect 18052 29708 18104 29714
rect 18052 29650 18104 29656
rect 16856 29096 16908 29102
rect 16856 29038 16908 29044
rect 16868 28626 16896 29038
rect 16856 28620 16908 28626
rect 16856 28562 16908 28568
rect 16764 28552 16816 28558
rect 16764 28494 16816 28500
rect 16868 27554 16896 28562
rect 18064 27606 18092 29650
rect 18144 29640 18196 29646
rect 18248 29594 18276 29786
rect 18196 29588 18276 29594
rect 18144 29582 18276 29588
rect 18156 29566 18276 29582
rect 18248 28762 18276 29566
rect 18315 28860 18623 28869
rect 18315 28858 18321 28860
rect 18377 28858 18401 28860
rect 18457 28858 18481 28860
rect 18537 28858 18561 28860
rect 18617 28858 18623 28860
rect 18377 28806 18379 28858
rect 18559 28806 18561 28858
rect 18315 28804 18321 28806
rect 18377 28804 18401 28806
rect 18457 28804 18481 28806
rect 18537 28804 18561 28806
rect 18617 28804 18623 28806
rect 18315 28795 18623 28804
rect 18236 28756 18288 28762
rect 18236 28698 18288 28704
rect 18236 28416 18288 28422
rect 18236 28358 18288 28364
rect 18248 28150 18276 28358
rect 18236 28144 18288 28150
rect 18236 28086 18288 28092
rect 18880 28076 18932 28082
rect 18880 28018 18932 28024
rect 18892 27985 18920 28018
rect 18878 27976 18934 27985
rect 18878 27911 18880 27920
rect 18932 27911 18934 27920
rect 18880 27882 18932 27888
rect 18788 27872 18840 27878
rect 18892 27851 18920 27882
rect 18788 27814 18840 27820
rect 18315 27772 18623 27781
rect 18315 27770 18321 27772
rect 18377 27770 18401 27772
rect 18457 27770 18481 27772
rect 18537 27770 18561 27772
rect 18617 27770 18623 27772
rect 18377 27718 18379 27770
rect 18559 27718 18561 27770
rect 18315 27716 18321 27718
rect 18377 27716 18401 27718
rect 18457 27716 18481 27718
rect 18537 27716 18561 27718
rect 18617 27716 18623 27718
rect 18315 27707 18623 27716
rect 16776 27526 16896 27554
rect 18052 27600 18104 27606
rect 18052 27542 18104 27548
rect 16776 27470 16804 27526
rect 18800 27470 18828 27814
rect 16764 27464 16816 27470
rect 16764 27406 16816 27412
rect 18788 27464 18840 27470
rect 18788 27406 18840 27412
rect 16672 26512 16724 26518
rect 16672 26454 16724 26460
rect 16776 25906 16804 27406
rect 17040 27396 17092 27402
rect 17040 27338 17092 27344
rect 17052 27130 17080 27338
rect 17040 27124 17092 27130
rect 17040 27066 17092 27072
rect 18800 26994 18828 27406
rect 18788 26988 18840 26994
rect 18788 26930 18840 26936
rect 17040 26784 17092 26790
rect 17040 26726 17092 26732
rect 17052 26382 17080 26726
rect 18315 26684 18623 26693
rect 18315 26682 18321 26684
rect 18377 26682 18401 26684
rect 18457 26682 18481 26684
rect 18537 26682 18561 26684
rect 18617 26682 18623 26684
rect 18377 26630 18379 26682
rect 18559 26630 18561 26682
rect 18315 26628 18321 26630
rect 18377 26628 18401 26630
rect 18457 26628 18481 26630
rect 18537 26628 18561 26630
rect 18617 26628 18623 26630
rect 18315 26619 18623 26628
rect 17408 26512 17460 26518
rect 17408 26454 17460 26460
rect 17040 26376 17092 26382
rect 17040 26318 17092 26324
rect 16764 25900 16816 25906
rect 16764 25842 16816 25848
rect 16856 24608 16908 24614
rect 16856 24550 16908 24556
rect 16868 24206 16896 24550
rect 16764 24200 16816 24206
rect 16764 24142 16816 24148
rect 16856 24200 16908 24206
rect 16856 24142 16908 24148
rect 16776 23662 16804 24142
rect 16856 24064 16908 24070
rect 16856 24006 16908 24012
rect 16868 23798 16896 24006
rect 16856 23792 16908 23798
rect 16856 23734 16908 23740
rect 16764 23656 16816 23662
rect 16764 23598 16816 23604
rect 16396 23112 16448 23118
rect 16396 23054 16448 23060
rect 16408 22234 16436 23054
rect 16580 22976 16632 22982
rect 16580 22918 16632 22924
rect 16592 22710 16620 22918
rect 16580 22704 16632 22710
rect 16580 22646 16632 22652
rect 16776 22574 16804 23598
rect 16672 22568 16724 22574
rect 16672 22510 16724 22516
rect 16764 22568 16816 22574
rect 16764 22510 16816 22516
rect 16396 22228 16448 22234
rect 16396 22170 16448 22176
rect 16580 22024 16632 22030
rect 16580 21966 16632 21972
rect 16212 21956 16264 21962
rect 16212 21898 16264 21904
rect 16224 20874 16252 21898
rect 16304 21344 16356 21350
rect 16304 21286 16356 21292
rect 16316 20942 16344 21286
rect 16592 21146 16620 21966
rect 16580 21140 16632 21146
rect 16580 21082 16632 21088
rect 16304 20936 16356 20942
rect 16304 20878 16356 20884
rect 16212 20868 16264 20874
rect 16212 20810 16264 20816
rect 15936 19780 15988 19786
rect 15936 19722 15988 19728
rect 15948 19378 15976 19722
rect 15936 19372 15988 19378
rect 15936 19314 15988 19320
rect 15948 18698 15976 19314
rect 15936 18692 15988 18698
rect 15936 18634 15988 18640
rect 16120 18352 16172 18358
rect 16120 18294 16172 18300
rect 16132 17882 16160 18294
rect 16120 17876 16172 17882
rect 16120 17818 16172 17824
rect 16224 17746 16252 20810
rect 16580 19848 16632 19854
rect 16580 19790 16632 19796
rect 16304 19372 16356 19378
rect 16304 19314 16356 19320
rect 16316 18426 16344 19314
rect 16592 18970 16620 19790
rect 16580 18964 16632 18970
rect 16580 18906 16632 18912
rect 16304 18420 16356 18426
rect 16304 18362 16356 18368
rect 16212 17740 16264 17746
rect 16212 17682 16264 17688
rect 15844 17672 15896 17678
rect 15844 17614 15896 17620
rect 15752 17332 15804 17338
rect 15752 17274 15804 17280
rect 15856 17202 15884 17614
rect 16580 17604 16632 17610
rect 16580 17546 16632 17552
rect 15844 17196 15896 17202
rect 15844 17138 15896 17144
rect 15660 16788 15712 16794
rect 15660 16730 15712 16736
rect 14842 16348 15150 16357
rect 14842 16346 14848 16348
rect 14904 16346 14928 16348
rect 14984 16346 15008 16348
rect 15064 16346 15088 16348
rect 15144 16346 15150 16348
rect 14904 16294 14906 16346
rect 15086 16294 15088 16346
rect 14842 16292 14848 16294
rect 14904 16292 14928 16294
rect 14984 16292 15008 16294
rect 15064 16292 15088 16294
rect 15144 16292 15150 16294
rect 14842 16283 15150 16292
rect 14842 15260 15150 15269
rect 14842 15258 14848 15260
rect 14904 15258 14928 15260
rect 14984 15258 15008 15260
rect 15064 15258 15088 15260
rect 15144 15258 15150 15260
rect 14904 15206 14906 15258
rect 15086 15206 15088 15258
rect 14842 15204 14848 15206
rect 14904 15204 14928 15206
rect 14984 15204 15008 15206
rect 15064 15204 15088 15206
rect 15144 15204 15150 15206
rect 14842 15195 15150 15204
rect 15672 14414 15700 16730
rect 15856 16522 15884 17138
rect 16592 17134 16620 17546
rect 16580 17128 16632 17134
rect 16580 17070 16632 17076
rect 16592 16794 16620 17070
rect 16580 16788 16632 16794
rect 16580 16730 16632 16736
rect 15844 16516 15896 16522
rect 15844 16458 15896 16464
rect 16212 14816 16264 14822
rect 16212 14758 16264 14764
rect 15660 14408 15712 14414
rect 15660 14350 15712 14356
rect 16120 14408 16172 14414
rect 16120 14350 16172 14356
rect 14842 14172 15150 14181
rect 14842 14170 14848 14172
rect 14904 14170 14928 14172
rect 14984 14170 15008 14172
rect 15064 14170 15088 14172
rect 15144 14170 15150 14172
rect 14904 14118 14906 14170
rect 15086 14118 15088 14170
rect 14842 14116 14848 14118
rect 14904 14116 14928 14118
rect 14984 14116 15008 14118
rect 15064 14116 15088 14118
rect 15144 14116 15150 14118
rect 14842 14107 15150 14116
rect 16132 13938 16160 14350
rect 16224 14346 16252 14758
rect 16212 14340 16264 14346
rect 16212 14282 16264 14288
rect 16224 13938 16252 14282
rect 16304 14272 16356 14278
rect 16304 14214 16356 14220
rect 16316 14074 16344 14214
rect 16304 14068 16356 14074
rect 16304 14010 16356 14016
rect 16120 13932 16172 13938
rect 16120 13874 16172 13880
rect 16212 13932 16264 13938
rect 16212 13874 16264 13880
rect 14842 13084 15150 13093
rect 14842 13082 14848 13084
rect 14904 13082 14928 13084
rect 14984 13082 15008 13084
rect 15064 13082 15088 13084
rect 15144 13082 15150 13084
rect 14904 13030 14906 13082
rect 15086 13030 15088 13082
rect 14842 13028 14848 13030
rect 14904 13028 14928 13030
rect 14984 13028 15008 13030
rect 15064 13028 15088 13030
rect 15144 13028 15150 13030
rect 14842 13019 15150 13028
rect 16684 12850 16712 22510
rect 16776 21554 16804 22510
rect 16948 21888 17000 21894
rect 16948 21830 17000 21836
rect 16960 21554 16988 21830
rect 16764 21548 16816 21554
rect 16764 21490 16816 21496
rect 16948 21548 17000 21554
rect 16948 21490 17000 21496
rect 16776 19378 16804 21490
rect 16856 21412 16908 21418
rect 16856 21354 16908 21360
rect 16764 19372 16816 19378
rect 16764 19314 16816 19320
rect 16776 18766 16804 19314
rect 16764 18760 16816 18766
rect 16764 18702 16816 18708
rect 16776 18358 16804 18702
rect 16868 18612 16896 21354
rect 16948 19508 17000 19514
rect 16948 19450 17000 19456
rect 16960 18766 16988 19450
rect 17052 18970 17080 26318
rect 17132 25900 17184 25906
rect 17132 25842 17184 25848
rect 17144 25498 17172 25842
rect 17132 25492 17184 25498
rect 17132 25434 17184 25440
rect 17132 25220 17184 25226
rect 17132 25162 17184 25168
rect 17144 24886 17172 25162
rect 17132 24880 17184 24886
rect 17132 24822 17184 24828
rect 17144 23798 17172 24822
rect 17224 24812 17276 24818
rect 17224 24754 17276 24760
rect 17236 23866 17264 24754
rect 17224 23860 17276 23866
rect 17224 23802 17276 23808
rect 17132 23792 17184 23798
rect 17132 23734 17184 23740
rect 17224 19712 17276 19718
rect 17224 19654 17276 19660
rect 17236 19446 17264 19654
rect 17224 19440 17276 19446
rect 17224 19382 17276 19388
rect 17132 19168 17184 19174
rect 17132 19110 17184 19116
rect 17040 18964 17092 18970
rect 17040 18906 17092 18912
rect 16948 18760 17000 18766
rect 16948 18702 17000 18708
rect 16868 18584 16988 18612
rect 16764 18352 16816 18358
rect 16764 18294 16816 18300
rect 16856 18080 16908 18086
rect 16856 18022 16908 18028
rect 16868 14346 16896 18022
rect 16856 14340 16908 14346
rect 16856 14282 16908 14288
rect 16868 13870 16896 14282
rect 16856 13864 16908 13870
rect 16856 13806 16908 13812
rect 16672 12844 16724 12850
rect 16672 12786 16724 12792
rect 16684 12434 16712 12786
rect 16960 12782 16988 18584
rect 17040 18284 17092 18290
rect 17144 18272 17172 19110
rect 17224 18624 17276 18630
rect 17224 18566 17276 18572
rect 17236 18426 17264 18566
rect 17224 18420 17276 18426
rect 17224 18362 17276 18368
rect 17092 18244 17172 18272
rect 17040 18226 17092 18232
rect 17052 16522 17080 18226
rect 17420 18086 17448 26454
rect 18880 25900 18932 25906
rect 18880 25842 18932 25848
rect 18315 25596 18623 25605
rect 18315 25594 18321 25596
rect 18377 25594 18401 25596
rect 18457 25594 18481 25596
rect 18537 25594 18561 25596
rect 18617 25594 18623 25596
rect 18377 25542 18379 25594
rect 18559 25542 18561 25594
rect 18315 25540 18321 25542
rect 18377 25540 18401 25542
rect 18457 25540 18481 25542
rect 18537 25540 18561 25542
rect 18617 25540 18623 25542
rect 18315 25531 18623 25540
rect 18892 25498 18920 25842
rect 18880 25492 18932 25498
rect 18880 25434 18932 25440
rect 18315 24508 18623 24517
rect 18315 24506 18321 24508
rect 18377 24506 18401 24508
rect 18457 24506 18481 24508
rect 18537 24506 18561 24508
rect 18617 24506 18623 24508
rect 18377 24454 18379 24506
rect 18559 24454 18561 24506
rect 18315 24452 18321 24454
rect 18377 24452 18401 24454
rect 18457 24452 18481 24454
rect 18537 24452 18561 24454
rect 18617 24452 18623 24454
rect 18315 24443 18623 24452
rect 18788 24200 18840 24206
rect 18788 24142 18840 24148
rect 18604 24064 18656 24070
rect 18604 24006 18656 24012
rect 18616 23798 18644 24006
rect 18604 23792 18656 23798
rect 18604 23734 18656 23740
rect 18315 23420 18623 23429
rect 18315 23418 18321 23420
rect 18377 23418 18401 23420
rect 18457 23418 18481 23420
rect 18537 23418 18561 23420
rect 18617 23418 18623 23420
rect 18377 23366 18379 23418
rect 18559 23366 18561 23418
rect 18315 23364 18321 23366
rect 18377 23364 18401 23366
rect 18457 23364 18481 23366
rect 18537 23364 18561 23366
rect 18617 23364 18623 23366
rect 18315 23355 18623 23364
rect 18800 23322 18828 24142
rect 18788 23316 18840 23322
rect 18788 23258 18840 23264
rect 18788 23044 18840 23050
rect 18788 22986 18840 22992
rect 18144 22772 18196 22778
rect 18144 22714 18196 22720
rect 18052 18828 18104 18834
rect 18052 18770 18104 18776
rect 17960 18624 18012 18630
rect 17960 18566 18012 18572
rect 17408 18080 17460 18086
rect 17408 18022 17460 18028
rect 17972 16794 18000 18566
rect 18064 18358 18092 18770
rect 18052 18352 18104 18358
rect 18052 18294 18104 18300
rect 18064 17202 18092 18294
rect 18052 17196 18104 17202
rect 18052 17138 18104 17144
rect 17684 16788 17736 16794
rect 17684 16730 17736 16736
rect 17960 16788 18012 16794
rect 17960 16730 18012 16736
rect 17040 16516 17092 16522
rect 17040 16458 17092 16464
rect 17132 16108 17184 16114
rect 17132 16050 17184 16056
rect 17040 13932 17092 13938
rect 17040 13874 17092 13880
rect 17052 13326 17080 13874
rect 17040 13320 17092 13326
rect 17040 13262 17092 13268
rect 16948 12776 17000 12782
rect 16948 12718 17000 12724
rect 17144 12442 17172 16050
rect 17224 15904 17276 15910
rect 17224 15846 17276 15852
rect 17132 12436 17184 12442
rect 16684 12406 16896 12434
rect 16672 12232 16724 12238
rect 16672 12174 16724 12180
rect 14842 11996 15150 12005
rect 14842 11994 14848 11996
rect 14904 11994 14928 11996
rect 14984 11994 15008 11996
rect 15064 11994 15088 11996
rect 15144 11994 15150 11996
rect 14904 11942 14906 11994
rect 15086 11942 15088 11994
rect 14842 11940 14848 11942
rect 14904 11940 14928 11942
rect 14984 11940 15008 11942
rect 15064 11940 15088 11942
rect 15144 11940 15150 11942
rect 14842 11931 15150 11940
rect 16684 11898 16712 12174
rect 16672 11892 16724 11898
rect 16672 11834 16724 11840
rect 14842 10908 15150 10917
rect 14842 10906 14848 10908
rect 14904 10906 14928 10908
rect 14984 10906 15008 10908
rect 15064 10906 15088 10908
rect 15144 10906 15150 10908
rect 14904 10854 14906 10906
rect 15086 10854 15088 10906
rect 14842 10852 14848 10854
rect 14904 10852 14928 10854
rect 14984 10852 15008 10854
rect 15064 10852 15088 10854
rect 15144 10852 15150 10854
rect 14842 10843 15150 10852
rect 14842 9820 15150 9829
rect 14842 9818 14848 9820
rect 14904 9818 14928 9820
rect 14984 9818 15008 9820
rect 15064 9818 15088 9820
rect 15144 9818 15150 9820
rect 14904 9766 14906 9818
rect 15086 9766 15088 9818
rect 14842 9764 14848 9766
rect 14904 9764 14928 9766
rect 14984 9764 15008 9766
rect 15064 9764 15088 9766
rect 15144 9764 15150 9766
rect 14842 9755 15150 9764
rect 14842 8732 15150 8741
rect 14842 8730 14848 8732
rect 14904 8730 14928 8732
rect 14984 8730 15008 8732
rect 15064 8730 15088 8732
rect 15144 8730 15150 8732
rect 14904 8678 14906 8730
rect 15086 8678 15088 8730
rect 14842 8676 14848 8678
rect 14904 8676 14928 8678
rect 14984 8676 15008 8678
rect 15064 8676 15088 8678
rect 15144 8676 15150 8678
rect 14842 8667 15150 8676
rect 14842 7644 15150 7653
rect 14842 7642 14848 7644
rect 14904 7642 14928 7644
rect 14984 7642 15008 7644
rect 15064 7642 15088 7644
rect 15144 7642 15150 7644
rect 14904 7590 14906 7642
rect 15086 7590 15088 7642
rect 14842 7588 14848 7590
rect 14904 7588 14928 7590
rect 14984 7588 15008 7590
rect 15064 7588 15088 7590
rect 15144 7588 15150 7590
rect 14842 7579 15150 7588
rect 14842 6556 15150 6565
rect 14842 6554 14848 6556
rect 14904 6554 14928 6556
rect 14984 6554 15008 6556
rect 15064 6554 15088 6556
rect 15144 6554 15150 6556
rect 14904 6502 14906 6554
rect 15086 6502 15088 6554
rect 14842 6500 14848 6502
rect 14904 6500 14928 6502
rect 14984 6500 15008 6502
rect 15064 6500 15088 6502
rect 15144 6500 15150 6502
rect 14842 6491 15150 6500
rect 14842 5468 15150 5477
rect 14842 5466 14848 5468
rect 14904 5466 14928 5468
rect 14984 5466 15008 5468
rect 15064 5466 15088 5468
rect 15144 5466 15150 5468
rect 14904 5414 14906 5466
rect 15086 5414 15088 5466
rect 14842 5412 14848 5414
rect 14904 5412 14928 5414
rect 14984 5412 15008 5414
rect 15064 5412 15088 5414
rect 15144 5412 15150 5414
rect 14842 5403 15150 5412
rect 16764 4548 16816 4554
rect 16764 4490 16816 4496
rect 14842 4380 15150 4389
rect 14842 4378 14848 4380
rect 14904 4378 14928 4380
rect 14984 4378 15008 4380
rect 15064 4378 15088 4380
rect 15144 4378 15150 4380
rect 14904 4326 14906 4378
rect 15086 4326 15088 4378
rect 14842 4324 14848 4326
rect 14904 4324 14928 4326
rect 14984 4324 15008 4326
rect 15064 4324 15088 4326
rect 15144 4324 15150 4326
rect 14842 4315 15150 4324
rect 16776 4078 16804 4490
rect 16764 4072 16816 4078
rect 16764 4014 16816 4020
rect 14188 4004 14240 4010
rect 14188 3946 14240 3952
rect 14556 4004 14608 4010
rect 14556 3946 14608 3952
rect 14200 3194 14228 3946
rect 16776 3534 16804 4014
rect 14280 3528 14332 3534
rect 14280 3470 14332 3476
rect 16304 3528 16356 3534
rect 16304 3470 16356 3476
rect 16764 3528 16816 3534
rect 16764 3470 16816 3476
rect 14188 3188 14240 3194
rect 14188 3130 14240 3136
rect 14200 2446 14228 3130
rect 14292 3058 14320 3470
rect 14842 3292 15150 3301
rect 14842 3290 14848 3292
rect 14904 3290 14928 3292
rect 14984 3290 15008 3292
rect 15064 3290 15088 3292
rect 15144 3290 15150 3292
rect 14904 3238 14906 3290
rect 15086 3238 15088 3290
rect 14842 3236 14848 3238
rect 14904 3236 14928 3238
rect 14984 3236 15008 3238
rect 15064 3236 15088 3238
rect 15144 3236 15150 3238
rect 14842 3227 15150 3236
rect 16316 3058 16344 3470
rect 14280 3052 14332 3058
rect 14280 2994 14332 3000
rect 16304 3052 16356 3058
rect 16304 2994 16356 3000
rect 14464 2984 14516 2990
rect 14464 2926 14516 2932
rect 14740 2984 14792 2990
rect 14740 2926 14792 2932
rect 16764 2984 16816 2990
rect 16764 2926 16816 2932
rect 14476 2650 14504 2926
rect 14464 2644 14516 2650
rect 14464 2586 14516 2592
rect 14188 2440 14240 2446
rect 14188 2382 14240 2388
rect 14752 1714 14780 2926
rect 16120 2372 16172 2378
rect 16120 2314 16172 2320
rect 14842 2204 15150 2213
rect 14842 2202 14848 2204
rect 14904 2202 14928 2204
rect 14984 2202 15008 2204
rect 15064 2202 15088 2204
rect 15144 2202 15150 2204
rect 14904 2150 14906 2202
rect 15086 2150 15088 2202
rect 14842 2148 14848 2150
rect 14904 2148 14928 2150
rect 14984 2148 15008 2150
rect 15064 2148 15088 2150
rect 15144 2148 15150 2150
rect 14842 2139 15150 2148
rect 14752 1686 14872 1714
rect 14844 800 14872 1686
rect 16132 800 16160 2314
rect 16776 800 16804 2926
rect 16868 2650 16896 12406
rect 17132 12378 17184 12384
rect 17236 11762 17264 15846
rect 17316 15428 17368 15434
rect 17316 15370 17368 15376
rect 17328 14074 17356 15370
rect 17408 14476 17460 14482
rect 17408 14418 17460 14424
rect 17316 14068 17368 14074
rect 17316 14010 17368 14016
rect 17420 13938 17448 14418
rect 17408 13932 17460 13938
rect 17408 13874 17460 13880
rect 17500 12708 17552 12714
rect 17500 12650 17552 12656
rect 17224 11756 17276 11762
rect 17224 11698 17276 11704
rect 17236 10606 17264 11698
rect 17512 11694 17540 12650
rect 17500 11688 17552 11694
rect 17500 11630 17552 11636
rect 17696 11150 17724 16730
rect 18064 16182 18092 17138
rect 18052 16176 18104 16182
rect 18052 16118 18104 16124
rect 18064 15502 18092 16118
rect 18052 15496 18104 15502
rect 18052 15438 18104 15444
rect 18064 15042 18092 15438
rect 18156 15144 18184 22714
rect 18315 22332 18623 22341
rect 18315 22330 18321 22332
rect 18377 22330 18401 22332
rect 18457 22330 18481 22332
rect 18537 22330 18561 22332
rect 18617 22330 18623 22332
rect 18377 22278 18379 22330
rect 18559 22278 18561 22330
rect 18315 22276 18321 22278
rect 18377 22276 18401 22278
rect 18457 22276 18481 22278
rect 18537 22276 18561 22278
rect 18617 22276 18623 22278
rect 18315 22267 18623 22276
rect 18315 21244 18623 21253
rect 18315 21242 18321 21244
rect 18377 21242 18401 21244
rect 18457 21242 18481 21244
rect 18537 21242 18561 21244
rect 18617 21242 18623 21244
rect 18377 21190 18379 21242
rect 18559 21190 18561 21242
rect 18315 21188 18321 21190
rect 18377 21188 18401 21190
rect 18457 21188 18481 21190
rect 18537 21188 18561 21190
rect 18617 21188 18623 21190
rect 18315 21179 18623 21188
rect 18800 21010 18828 22986
rect 18984 22094 19012 32778
rect 19168 32502 19196 32778
rect 19156 32496 19208 32502
rect 19156 32438 19208 32444
rect 19352 32434 19380 33254
rect 19444 33114 19472 33526
rect 19432 33108 19484 33114
rect 19432 33050 19484 33056
rect 19628 32910 19656 34546
rect 19708 34536 19760 34542
rect 19708 34478 19760 34484
rect 19616 32904 19668 32910
rect 19616 32846 19668 32852
rect 19340 32428 19392 32434
rect 19340 32370 19392 32376
rect 19064 32224 19116 32230
rect 19064 32166 19116 32172
rect 19076 28422 19104 32166
rect 19616 30048 19668 30054
rect 19616 29990 19668 29996
rect 19524 29708 19576 29714
rect 19524 29650 19576 29656
rect 19536 29594 19564 29650
rect 19628 29646 19656 29990
rect 19444 29566 19564 29594
rect 19616 29640 19668 29646
rect 19616 29582 19668 29588
rect 19444 29102 19472 29566
rect 19524 29504 19576 29510
rect 19524 29446 19576 29452
rect 19432 29096 19484 29102
rect 19432 29038 19484 29044
rect 19444 28626 19472 29038
rect 19432 28620 19484 28626
rect 19432 28562 19484 28568
rect 19064 28416 19116 28422
rect 19064 28358 19116 28364
rect 19076 28082 19104 28358
rect 19064 28076 19116 28082
rect 19064 28018 19116 28024
rect 19156 28076 19208 28082
rect 19156 28018 19208 28024
rect 18984 22066 19104 22094
rect 19076 21690 19104 22066
rect 19064 21684 19116 21690
rect 19064 21626 19116 21632
rect 18972 21548 19024 21554
rect 18972 21490 19024 21496
rect 18788 21004 18840 21010
rect 18788 20946 18840 20952
rect 18696 20800 18748 20806
rect 18696 20742 18748 20748
rect 18708 20466 18736 20742
rect 18696 20460 18748 20466
rect 18696 20402 18748 20408
rect 18315 20156 18623 20165
rect 18315 20154 18321 20156
rect 18377 20154 18401 20156
rect 18457 20154 18481 20156
rect 18537 20154 18561 20156
rect 18617 20154 18623 20156
rect 18377 20102 18379 20154
rect 18559 20102 18561 20154
rect 18315 20100 18321 20102
rect 18377 20100 18401 20102
rect 18457 20100 18481 20102
rect 18537 20100 18561 20102
rect 18617 20100 18623 20102
rect 18315 20091 18623 20100
rect 18315 19068 18623 19077
rect 18315 19066 18321 19068
rect 18377 19066 18401 19068
rect 18457 19066 18481 19068
rect 18537 19066 18561 19068
rect 18617 19066 18623 19068
rect 18377 19014 18379 19066
rect 18559 19014 18561 19066
rect 18315 19012 18321 19014
rect 18377 19012 18401 19014
rect 18457 19012 18481 19014
rect 18537 19012 18561 19014
rect 18617 19012 18623 19014
rect 18315 19003 18623 19012
rect 18696 18760 18748 18766
rect 18696 18702 18748 18708
rect 18236 18624 18288 18630
rect 18236 18566 18288 18572
rect 18248 17252 18276 18566
rect 18315 17980 18623 17989
rect 18315 17978 18321 17980
rect 18377 17978 18401 17980
rect 18457 17978 18481 17980
rect 18537 17978 18561 17980
rect 18617 17978 18623 17980
rect 18377 17926 18379 17978
rect 18559 17926 18561 17978
rect 18315 17924 18321 17926
rect 18377 17924 18401 17926
rect 18457 17924 18481 17926
rect 18537 17924 18561 17926
rect 18617 17924 18623 17926
rect 18315 17915 18623 17924
rect 18708 17882 18736 18702
rect 18696 17876 18748 17882
rect 18696 17818 18748 17824
rect 18800 17678 18828 20946
rect 18984 20602 19012 21490
rect 18972 20596 19024 20602
rect 18972 20538 19024 20544
rect 18788 17672 18840 17678
rect 18788 17614 18840 17620
rect 18328 17264 18380 17270
rect 18248 17224 18328 17252
rect 18328 17206 18380 17212
rect 18315 16892 18623 16901
rect 18315 16890 18321 16892
rect 18377 16890 18401 16892
rect 18457 16890 18481 16892
rect 18537 16890 18561 16892
rect 18617 16890 18623 16892
rect 18377 16838 18379 16890
rect 18559 16838 18561 16890
rect 18315 16836 18321 16838
rect 18377 16836 18401 16838
rect 18457 16836 18481 16838
rect 18537 16836 18561 16838
rect 18617 16836 18623 16838
rect 18315 16827 18623 16836
rect 18880 16516 18932 16522
rect 18880 16458 18932 16464
rect 18315 15804 18623 15813
rect 18315 15802 18321 15804
rect 18377 15802 18401 15804
rect 18457 15802 18481 15804
rect 18537 15802 18561 15804
rect 18617 15802 18623 15804
rect 18377 15750 18379 15802
rect 18559 15750 18561 15802
rect 18315 15748 18321 15750
rect 18377 15748 18401 15750
rect 18457 15748 18481 15750
rect 18537 15748 18561 15750
rect 18617 15748 18623 15750
rect 18315 15739 18623 15748
rect 18696 15360 18748 15366
rect 18696 15302 18748 15308
rect 18156 15116 18276 15144
rect 18064 15026 18184 15042
rect 17960 15020 18012 15026
rect 18064 15020 18196 15026
rect 18064 15014 18144 15020
rect 17960 14962 18012 14968
rect 18144 14962 18196 14968
rect 17972 14618 18000 14962
rect 17960 14612 18012 14618
rect 17960 14554 18012 14560
rect 18144 13796 18196 13802
rect 18144 13738 18196 13744
rect 17960 13728 18012 13734
rect 17960 13670 18012 13676
rect 18052 13728 18104 13734
rect 18052 13670 18104 13676
rect 17972 13190 18000 13670
rect 18064 13530 18092 13670
rect 18052 13524 18104 13530
rect 18052 13466 18104 13472
rect 17960 13184 18012 13190
rect 17960 13126 18012 13132
rect 17684 11144 17736 11150
rect 17684 11086 17736 11092
rect 17776 11008 17828 11014
rect 17776 10950 17828 10956
rect 17788 10742 17816 10950
rect 17776 10736 17828 10742
rect 17776 10678 17828 10684
rect 17972 10606 18000 13126
rect 18064 12850 18092 13466
rect 18156 13326 18184 13738
rect 18248 13512 18276 15116
rect 18315 14716 18623 14725
rect 18315 14714 18321 14716
rect 18377 14714 18401 14716
rect 18457 14714 18481 14716
rect 18537 14714 18561 14716
rect 18617 14714 18623 14716
rect 18377 14662 18379 14714
rect 18559 14662 18561 14714
rect 18315 14660 18321 14662
rect 18377 14660 18401 14662
rect 18457 14660 18481 14662
rect 18537 14660 18561 14662
rect 18617 14660 18623 14662
rect 18315 14651 18623 14660
rect 18708 13938 18736 15302
rect 18696 13932 18748 13938
rect 18696 13874 18748 13880
rect 18315 13628 18623 13637
rect 18315 13626 18321 13628
rect 18377 13626 18401 13628
rect 18457 13626 18481 13628
rect 18537 13626 18561 13628
rect 18617 13626 18623 13628
rect 18377 13574 18379 13626
rect 18559 13574 18561 13626
rect 18315 13572 18321 13574
rect 18377 13572 18401 13574
rect 18457 13572 18481 13574
rect 18537 13572 18561 13574
rect 18617 13572 18623 13574
rect 18315 13563 18623 13572
rect 18248 13484 18368 13512
rect 18340 13326 18368 13484
rect 18144 13320 18196 13326
rect 18144 13262 18196 13268
rect 18328 13320 18380 13326
rect 18328 13262 18380 13268
rect 18052 12844 18104 12850
rect 18052 12786 18104 12792
rect 18708 12646 18736 13874
rect 18788 13184 18840 13190
rect 18788 13126 18840 13132
rect 18236 12640 18288 12646
rect 18236 12582 18288 12588
rect 18696 12640 18748 12646
rect 18696 12582 18748 12588
rect 18248 11830 18276 12582
rect 18315 12540 18623 12549
rect 18315 12538 18321 12540
rect 18377 12538 18401 12540
rect 18457 12538 18481 12540
rect 18537 12538 18561 12540
rect 18617 12538 18623 12540
rect 18377 12486 18379 12538
rect 18559 12486 18561 12538
rect 18315 12484 18321 12486
rect 18377 12484 18401 12486
rect 18457 12484 18481 12486
rect 18537 12484 18561 12486
rect 18617 12484 18623 12486
rect 18315 12475 18623 12484
rect 18236 11824 18288 11830
rect 18236 11766 18288 11772
rect 18052 11756 18104 11762
rect 18052 11698 18104 11704
rect 17224 10600 17276 10606
rect 17224 10542 17276 10548
rect 17960 10600 18012 10606
rect 17960 10542 18012 10548
rect 17972 10062 18000 10542
rect 17960 10056 18012 10062
rect 17960 9998 18012 10004
rect 17132 4140 17184 4146
rect 17132 4082 17184 4088
rect 17144 3398 17172 4082
rect 17224 3936 17276 3942
rect 17224 3878 17276 3884
rect 17040 3392 17092 3398
rect 17040 3334 17092 3340
rect 17132 3392 17184 3398
rect 17132 3334 17184 3340
rect 17052 3126 17080 3334
rect 17144 3194 17172 3334
rect 17132 3188 17184 3194
rect 17132 3130 17184 3136
rect 17040 3120 17092 3126
rect 17040 3062 17092 3068
rect 16856 2644 16908 2650
rect 16856 2586 16908 2592
rect 17236 2514 17264 3878
rect 18064 3738 18092 11698
rect 18248 10810 18276 11766
rect 18800 11762 18828 13126
rect 18892 12850 18920 16458
rect 18972 13320 19024 13326
rect 18972 13262 19024 13268
rect 18880 12844 18932 12850
rect 18880 12786 18932 12792
rect 18878 11928 18934 11937
rect 18878 11863 18880 11872
rect 18932 11863 18934 11872
rect 18880 11834 18932 11840
rect 18788 11756 18840 11762
rect 18788 11698 18840 11704
rect 18315 11452 18623 11461
rect 18315 11450 18321 11452
rect 18377 11450 18401 11452
rect 18457 11450 18481 11452
rect 18537 11450 18561 11452
rect 18617 11450 18623 11452
rect 18377 11398 18379 11450
rect 18559 11398 18561 11450
rect 18315 11396 18321 11398
rect 18377 11396 18401 11398
rect 18457 11396 18481 11398
rect 18537 11396 18561 11398
rect 18617 11396 18623 11398
rect 18315 11387 18623 11396
rect 18800 11354 18828 11698
rect 18880 11688 18932 11694
rect 18880 11630 18932 11636
rect 18788 11348 18840 11354
rect 18788 11290 18840 11296
rect 18328 11076 18380 11082
rect 18328 11018 18380 11024
rect 18236 10804 18288 10810
rect 18236 10746 18288 10752
rect 18340 10554 18368 11018
rect 18892 10810 18920 11630
rect 18880 10804 18932 10810
rect 18880 10746 18932 10752
rect 18984 10690 19012 13262
rect 19168 11354 19196 28018
rect 19444 27538 19472 28562
rect 19536 28558 19564 29446
rect 19524 28552 19576 28558
rect 19524 28494 19576 28500
rect 19432 27532 19484 27538
rect 19432 27474 19484 27480
rect 19432 26376 19484 26382
rect 19432 26318 19484 26324
rect 19444 24410 19472 26318
rect 19720 25294 19748 34478
rect 20548 33538 20576 35226
rect 20720 33856 20772 33862
rect 20720 33798 20772 33804
rect 20732 33590 20760 33798
rect 20456 33522 20576 33538
rect 20720 33584 20772 33590
rect 20720 33526 20772 33532
rect 20444 33516 20576 33522
rect 20496 33510 20576 33516
rect 20444 33458 20496 33464
rect 19984 33448 20036 33454
rect 19984 33390 20036 33396
rect 19892 33108 19944 33114
rect 19892 33050 19944 33056
rect 19904 32978 19932 33050
rect 19892 32972 19944 32978
rect 19892 32914 19944 32920
rect 19996 32910 20024 33390
rect 20456 33114 20484 33458
rect 20732 33114 20760 33526
rect 20444 33108 20496 33114
rect 20444 33050 20496 33056
rect 20720 33108 20772 33114
rect 20720 33050 20772 33056
rect 20352 33040 20404 33046
rect 20352 32982 20404 32988
rect 19800 32904 19852 32910
rect 19800 32846 19852 32852
rect 19984 32904 20036 32910
rect 19984 32846 20036 32852
rect 19812 32026 19840 32846
rect 20364 32434 20392 32982
rect 20824 32910 20852 35866
rect 20904 33652 20956 33658
rect 20904 33594 20956 33600
rect 20916 33046 20944 33594
rect 20904 33040 20956 33046
rect 20904 32982 20956 32988
rect 20812 32904 20864 32910
rect 20812 32846 20864 32852
rect 20536 32768 20588 32774
rect 20536 32710 20588 32716
rect 20548 32570 20576 32710
rect 20536 32564 20588 32570
rect 20536 32506 20588 32512
rect 20824 32502 20852 32846
rect 20812 32496 20864 32502
rect 20812 32438 20864 32444
rect 20076 32428 20128 32434
rect 20076 32370 20128 32376
rect 20352 32428 20404 32434
rect 20352 32370 20404 32376
rect 19800 32020 19852 32026
rect 19800 31962 19852 31968
rect 19892 28076 19944 28082
rect 19892 28018 19944 28024
rect 19904 26042 19932 28018
rect 20088 26586 20116 32370
rect 20168 32360 20220 32366
rect 20168 32302 20220 32308
rect 20180 30190 20208 32302
rect 20168 30184 20220 30190
rect 20168 30126 20220 30132
rect 20180 28762 20208 30126
rect 20168 28756 20220 28762
rect 20168 28698 20220 28704
rect 20364 28218 20392 32370
rect 21008 32366 21036 37198
rect 21376 36922 21404 37266
rect 21364 36916 21416 36922
rect 21364 36858 21416 36864
rect 21376 35894 21404 36858
rect 21456 36780 21508 36786
rect 21456 36722 21508 36728
rect 21100 35866 21404 35894
rect 20996 32360 21048 32366
rect 20996 32302 21048 32308
rect 20904 32020 20956 32026
rect 20904 31962 20956 31968
rect 20916 31822 20944 31962
rect 20904 31816 20956 31822
rect 20904 31758 20956 31764
rect 20536 30320 20588 30326
rect 20536 30262 20588 30268
rect 20548 28558 20576 30262
rect 20812 30048 20864 30054
rect 20812 29990 20864 29996
rect 20824 29714 20852 29990
rect 20812 29708 20864 29714
rect 20812 29650 20864 29656
rect 20916 29594 20944 31758
rect 20996 30252 21048 30258
rect 20996 30194 21048 30200
rect 20732 29566 20944 29594
rect 20536 28552 20588 28558
rect 20536 28494 20588 28500
rect 20352 28212 20404 28218
rect 20352 28154 20404 28160
rect 20548 27878 20576 28494
rect 20536 27872 20588 27878
rect 20536 27814 20588 27820
rect 20076 26580 20128 26586
rect 20076 26522 20128 26528
rect 19892 26036 19944 26042
rect 19892 25978 19944 25984
rect 20168 25900 20220 25906
rect 20168 25842 20220 25848
rect 19984 25832 20036 25838
rect 19984 25774 20036 25780
rect 19708 25288 19760 25294
rect 19708 25230 19760 25236
rect 19432 24404 19484 24410
rect 19432 24346 19484 24352
rect 19616 23520 19668 23526
rect 19616 23462 19668 23468
rect 19628 23118 19656 23462
rect 19616 23112 19668 23118
rect 19616 23054 19668 23060
rect 19524 20936 19576 20942
rect 19524 20878 19576 20884
rect 19536 20602 19564 20878
rect 19524 20596 19576 20602
rect 19524 20538 19576 20544
rect 19628 19514 19656 23054
rect 19720 23050 19748 25230
rect 19996 23186 20024 25774
rect 20180 25702 20208 25842
rect 20168 25696 20220 25702
rect 20168 25638 20220 25644
rect 20076 24200 20128 24206
rect 20076 24142 20128 24148
rect 20088 23866 20116 24142
rect 20076 23860 20128 23866
rect 20076 23802 20128 23808
rect 19984 23180 20036 23186
rect 19984 23122 20036 23128
rect 19708 23044 19760 23050
rect 19708 22986 19760 22992
rect 19708 22024 19760 22030
rect 19708 21966 19760 21972
rect 19720 21146 19748 21966
rect 19708 21140 19760 21146
rect 19708 21082 19760 21088
rect 19720 20534 19748 21082
rect 19800 20596 19852 20602
rect 19800 20538 19852 20544
rect 19708 20528 19760 20534
rect 19708 20470 19760 20476
rect 19616 19508 19668 19514
rect 19616 19450 19668 19456
rect 19340 19372 19392 19378
rect 19340 19314 19392 19320
rect 19248 16584 19300 16590
rect 19248 16526 19300 16532
rect 19260 15502 19288 16526
rect 19248 15496 19300 15502
rect 19248 15438 19300 15444
rect 19260 15094 19288 15438
rect 19248 15088 19300 15094
rect 19248 15030 19300 15036
rect 19352 14890 19380 19314
rect 19812 18766 19840 20538
rect 19996 20398 20024 23122
rect 20088 23118 20116 23802
rect 20076 23112 20128 23118
rect 20076 23054 20128 23060
rect 20076 21344 20128 21350
rect 20076 21286 20128 21292
rect 20088 20602 20116 21286
rect 20076 20596 20128 20602
rect 20076 20538 20128 20544
rect 19984 20392 20036 20398
rect 19984 20334 20036 20340
rect 19800 18760 19852 18766
rect 19800 18702 19852 18708
rect 19996 18086 20024 20334
rect 19984 18080 20036 18086
rect 19984 18022 20036 18028
rect 19892 17672 19944 17678
rect 19892 17614 19944 17620
rect 19800 17604 19852 17610
rect 19800 17546 19852 17552
rect 19812 17066 19840 17546
rect 19800 17060 19852 17066
rect 19800 17002 19852 17008
rect 19708 15428 19760 15434
rect 19708 15370 19760 15376
rect 19340 14884 19392 14890
rect 19340 14826 19392 14832
rect 19720 14618 19748 15370
rect 19708 14612 19760 14618
rect 19708 14554 19760 14560
rect 19432 14408 19484 14414
rect 19432 14350 19484 14356
rect 19444 14074 19472 14350
rect 19432 14068 19484 14074
rect 19432 14010 19484 14016
rect 19904 13938 19932 17614
rect 19996 17134 20024 18022
rect 20180 17746 20208 25638
rect 20548 22778 20576 27814
rect 20732 27130 20760 29566
rect 20904 29504 20956 29510
rect 20904 29446 20956 29452
rect 20916 29170 20944 29446
rect 21008 29306 21036 30194
rect 20996 29300 21048 29306
rect 20996 29242 21048 29248
rect 21100 29170 21128 35866
rect 21468 34202 21496 36722
rect 21652 35290 21680 37742
rect 22376 37664 22428 37670
rect 22376 37606 22428 37612
rect 21788 37020 22096 37029
rect 21788 37018 21794 37020
rect 21850 37018 21874 37020
rect 21930 37018 21954 37020
rect 22010 37018 22034 37020
rect 22090 37018 22096 37020
rect 21850 36966 21852 37018
rect 22032 36966 22034 37018
rect 21788 36964 21794 36966
rect 21850 36964 21874 36966
rect 21930 36964 21954 36966
rect 22010 36964 22034 36966
rect 22090 36964 22096 36966
rect 21788 36955 22096 36964
rect 21788 35932 22096 35941
rect 21788 35930 21794 35932
rect 21850 35930 21874 35932
rect 21930 35930 21954 35932
rect 22010 35930 22034 35932
rect 22090 35930 22096 35932
rect 21850 35878 21852 35930
rect 22032 35878 22034 35930
rect 21788 35876 21794 35878
rect 21850 35876 21874 35878
rect 21930 35876 21954 35878
rect 22010 35876 22034 35878
rect 22090 35876 22096 35878
rect 21788 35867 22096 35876
rect 21640 35284 21692 35290
rect 21640 35226 21692 35232
rect 21456 34196 21508 34202
rect 21456 34138 21508 34144
rect 21652 33658 21680 35226
rect 22388 35086 22416 37606
rect 23584 36242 23612 45766
rect 24320 45490 24348 46446
rect 24308 45484 24360 45490
rect 24308 45426 24360 45432
rect 24780 45082 24808 46990
rect 24952 46980 25004 46986
rect 26146 46951 26202 46960
rect 26700 46980 26752 46986
rect 24952 46922 25004 46928
rect 24964 45082 24992 46922
rect 26054 46336 26110 46345
rect 25261 46268 25569 46277
rect 26054 46271 26110 46280
rect 25261 46266 25267 46268
rect 25323 46266 25347 46268
rect 25403 46266 25427 46268
rect 25483 46266 25507 46268
rect 25563 46266 25569 46268
rect 25323 46214 25325 46266
rect 25505 46214 25507 46266
rect 25261 46212 25267 46214
rect 25323 46212 25347 46214
rect 25403 46212 25427 46214
rect 25483 46212 25507 46214
rect 25563 46212 25569 46214
rect 25261 46203 25569 46212
rect 25136 45892 25188 45898
rect 25136 45834 25188 45840
rect 24768 45076 24820 45082
rect 24768 45018 24820 45024
rect 24952 45076 25004 45082
rect 24952 45018 25004 45024
rect 25148 44946 25176 45834
rect 25780 45416 25832 45422
rect 25780 45358 25832 45364
rect 25261 45180 25569 45189
rect 25261 45178 25267 45180
rect 25323 45178 25347 45180
rect 25403 45178 25427 45180
rect 25483 45178 25507 45180
rect 25563 45178 25569 45180
rect 25323 45126 25325 45178
rect 25505 45126 25507 45178
rect 25261 45124 25267 45126
rect 25323 45124 25347 45126
rect 25403 45124 25427 45126
rect 25483 45124 25507 45126
rect 25563 45124 25569 45126
rect 25261 45115 25569 45124
rect 25136 44940 25188 44946
rect 25136 44882 25188 44888
rect 25261 44092 25569 44101
rect 25261 44090 25267 44092
rect 25323 44090 25347 44092
rect 25403 44090 25427 44092
rect 25483 44090 25507 44092
rect 25563 44090 25569 44092
rect 25323 44038 25325 44090
rect 25505 44038 25507 44090
rect 25261 44036 25267 44038
rect 25323 44036 25347 44038
rect 25403 44036 25427 44038
rect 25483 44036 25507 44038
rect 25563 44036 25569 44038
rect 25261 44027 25569 44036
rect 25792 43314 25820 45358
rect 25964 44940 26016 44946
rect 25964 44882 26016 44888
rect 25872 44872 25924 44878
rect 25872 44814 25924 44820
rect 25884 43858 25912 44814
rect 25872 43852 25924 43858
rect 25872 43794 25924 43800
rect 25780 43308 25832 43314
rect 25780 43250 25832 43256
rect 25261 43004 25569 43013
rect 25261 43002 25267 43004
rect 25323 43002 25347 43004
rect 25403 43002 25427 43004
rect 25483 43002 25507 43004
rect 25563 43002 25569 43004
rect 25323 42950 25325 43002
rect 25505 42950 25507 43002
rect 25261 42948 25267 42950
rect 25323 42948 25347 42950
rect 25403 42948 25427 42950
rect 25483 42948 25507 42950
rect 25563 42948 25569 42950
rect 25261 42939 25569 42948
rect 25261 41916 25569 41925
rect 25261 41914 25267 41916
rect 25323 41914 25347 41916
rect 25403 41914 25427 41916
rect 25483 41914 25507 41916
rect 25563 41914 25569 41916
rect 25323 41862 25325 41914
rect 25505 41862 25507 41914
rect 25261 41860 25267 41862
rect 25323 41860 25347 41862
rect 25403 41860 25427 41862
rect 25483 41860 25507 41862
rect 25563 41860 25569 41862
rect 25261 41851 25569 41860
rect 25261 40828 25569 40837
rect 25261 40826 25267 40828
rect 25323 40826 25347 40828
rect 25403 40826 25427 40828
rect 25483 40826 25507 40828
rect 25563 40826 25569 40828
rect 25323 40774 25325 40826
rect 25505 40774 25507 40826
rect 25261 40772 25267 40774
rect 25323 40772 25347 40774
rect 25403 40772 25427 40774
rect 25483 40772 25507 40774
rect 25563 40772 25569 40774
rect 25261 40763 25569 40772
rect 25261 39740 25569 39749
rect 25261 39738 25267 39740
rect 25323 39738 25347 39740
rect 25403 39738 25427 39740
rect 25483 39738 25507 39740
rect 25563 39738 25569 39740
rect 25323 39686 25325 39738
rect 25505 39686 25507 39738
rect 25261 39684 25267 39686
rect 25323 39684 25347 39686
rect 25403 39684 25427 39686
rect 25483 39684 25507 39686
rect 25563 39684 25569 39686
rect 25261 39675 25569 39684
rect 25261 38652 25569 38661
rect 25261 38650 25267 38652
rect 25323 38650 25347 38652
rect 25403 38650 25427 38652
rect 25483 38650 25507 38652
rect 25563 38650 25569 38652
rect 25323 38598 25325 38650
rect 25505 38598 25507 38650
rect 25261 38596 25267 38598
rect 25323 38596 25347 38598
rect 25403 38596 25427 38598
rect 25483 38596 25507 38598
rect 25563 38596 25569 38598
rect 25261 38587 25569 38596
rect 25261 37564 25569 37573
rect 25261 37562 25267 37564
rect 25323 37562 25347 37564
rect 25403 37562 25427 37564
rect 25483 37562 25507 37564
rect 25563 37562 25569 37564
rect 25323 37510 25325 37562
rect 25505 37510 25507 37562
rect 25261 37508 25267 37510
rect 25323 37508 25347 37510
rect 25403 37508 25427 37510
rect 25483 37508 25507 37510
rect 25563 37508 25569 37510
rect 25261 37499 25569 37508
rect 24860 36780 24912 36786
rect 24860 36722 24912 36728
rect 24676 36576 24728 36582
rect 24676 36518 24728 36524
rect 24768 36576 24820 36582
rect 24768 36518 24820 36524
rect 23572 36236 23624 36242
rect 23572 36178 23624 36184
rect 24492 36236 24544 36242
rect 24492 36178 24544 36184
rect 23480 36168 23532 36174
rect 23480 36110 23532 36116
rect 22652 36032 22704 36038
rect 22652 35974 22704 35980
rect 23112 36032 23164 36038
rect 23112 35974 23164 35980
rect 22664 35698 22692 35974
rect 22468 35692 22520 35698
rect 22652 35692 22704 35698
rect 22520 35652 22600 35680
rect 22468 35634 22520 35640
rect 22572 35086 22600 35652
rect 22652 35634 22704 35640
rect 23124 35086 23152 35974
rect 23492 35290 23520 36110
rect 23756 36032 23808 36038
rect 23756 35974 23808 35980
rect 23768 35494 23796 35974
rect 23756 35488 23808 35494
rect 23756 35430 23808 35436
rect 24124 35488 24176 35494
rect 24124 35430 24176 35436
rect 23480 35284 23532 35290
rect 23480 35226 23532 35232
rect 22376 35080 22428 35086
rect 22376 35022 22428 35028
rect 22560 35080 22612 35086
rect 22560 35022 22612 35028
rect 23112 35080 23164 35086
rect 23112 35022 23164 35028
rect 21788 34844 22096 34853
rect 21788 34842 21794 34844
rect 21850 34842 21874 34844
rect 21930 34842 21954 34844
rect 22010 34842 22034 34844
rect 22090 34842 22096 34844
rect 21850 34790 21852 34842
rect 22032 34790 22034 34842
rect 21788 34788 21794 34790
rect 21850 34788 21874 34790
rect 21930 34788 21954 34790
rect 22010 34788 22034 34790
rect 22090 34788 22096 34790
rect 21788 34779 22096 34788
rect 22468 33992 22520 33998
rect 22572 33980 22600 35022
rect 22744 35012 22796 35018
rect 22744 34954 22796 34960
rect 22520 33952 22600 33980
rect 22468 33934 22520 33940
rect 22192 33924 22244 33930
rect 22192 33866 22244 33872
rect 21788 33756 22096 33765
rect 21788 33754 21794 33756
rect 21850 33754 21874 33756
rect 21930 33754 21954 33756
rect 22010 33754 22034 33756
rect 22090 33754 22096 33756
rect 21850 33702 21852 33754
rect 22032 33702 22034 33754
rect 21788 33700 21794 33702
rect 21850 33700 21874 33702
rect 21930 33700 21954 33702
rect 22010 33700 22034 33702
rect 22090 33700 22096 33702
rect 21788 33691 22096 33700
rect 22204 33658 22232 33866
rect 21640 33652 21692 33658
rect 21640 33594 21692 33600
rect 22192 33652 22244 33658
rect 22192 33594 22244 33600
rect 22284 33516 22336 33522
rect 22284 33458 22336 33464
rect 21916 33312 21968 33318
rect 21916 33254 21968 33260
rect 21928 32910 21956 33254
rect 21916 32904 21968 32910
rect 21916 32846 21968 32852
rect 22192 32904 22244 32910
rect 22192 32846 22244 32852
rect 21788 32668 22096 32677
rect 21788 32666 21794 32668
rect 21850 32666 21874 32668
rect 21930 32666 21954 32668
rect 22010 32666 22034 32668
rect 22090 32666 22096 32668
rect 21850 32614 21852 32666
rect 22032 32614 22034 32666
rect 21788 32612 21794 32614
rect 21850 32612 21874 32614
rect 21930 32612 21954 32614
rect 22010 32612 22034 32614
rect 22090 32612 22096 32614
rect 21788 32603 22096 32612
rect 22100 32428 22152 32434
rect 22204 32416 22232 32846
rect 22152 32388 22232 32416
rect 22100 32370 22152 32376
rect 21640 32224 21692 32230
rect 21640 32166 21692 32172
rect 21652 31822 21680 32166
rect 21548 31816 21600 31822
rect 21548 31758 21600 31764
rect 21640 31816 21692 31822
rect 21640 31758 21692 31764
rect 21180 30320 21232 30326
rect 21180 30262 21232 30268
rect 21192 29646 21220 30262
rect 21180 29640 21232 29646
rect 21180 29582 21232 29588
rect 20904 29164 20956 29170
rect 20904 29106 20956 29112
rect 21088 29164 21140 29170
rect 21088 29106 21140 29112
rect 20812 27396 20864 27402
rect 20812 27338 20864 27344
rect 20720 27124 20772 27130
rect 20720 27066 20772 27072
rect 20628 25696 20680 25702
rect 20628 25638 20680 25644
rect 20640 25362 20668 25638
rect 20824 25498 20852 27338
rect 20916 25838 20944 29106
rect 21100 28150 21128 29106
rect 21088 28144 21140 28150
rect 21088 28086 21140 28092
rect 21192 26994 21220 29582
rect 21560 28762 21588 31758
rect 21652 29102 21680 31758
rect 21788 31580 22096 31589
rect 21788 31578 21794 31580
rect 21850 31578 21874 31580
rect 21930 31578 21954 31580
rect 22010 31578 22034 31580
rect 22090 31578 22096 31580
rect 21850 31526 21852 31578
rect 22032 31526 22034 31578
rect 21788 31524 21794 31526
rect 21850 31524 21874 31526
rect 21930 31524 21954 31526
rect 22010 31524 22034 31526
rect 22090 31524 22096 31526
rect 21788 31515 22096 31524
rect 22204 30598 22232 32388
rect 22296 32026 22324 33458
rect 22480 32910 22508 33934
rect 22468 32904 22520 32910
rect 22468 32846 22520 32852
rect 22652 32428 22704 32434
rect 22652 32370 22704 32376
rect 22284 32020 22336 32026
rect 22284 31962 22336 31968
rect 22664 31482 22692 32370
rect 22756 31890 22784 34954
rect 23768 33998 23796 35430
rect 24136 35018 24164 35430
rect 24124 35012 24176 35018
rect 24124 34954 24176 34960
rect 23756 33992 23808 33998
rect 23756 33934 23808 33940
rect 23388 33516 23440 33522
rect 23388 33458 23440 33464
rect 24032 33516 24084 33522
rect 24032 33458 24084 33464
rect 23204 33312 23256 33318
rect 23204 33254 23256 33260
rect 23216 32910 23244 33254
rect 23204 32904 23256 32910
rect 23204 32846 23256 32852
rect 23400 32026 23428 33458
rect 24044 33114 24072 33458
rect 24032 33108 24084 33114
rect 24032 33050 24084 33056
rect 24044 32570 24072 33050
rect 24032 32564 24084 32570
rect 24032 32506 24084 32512
rect 23480 32224 23532 32230
rect 23480 32166 23532 32172
rect 23664 32224 23716 32230
rect 23664 32166 23716 32172
rect 23388 32020 23440 32026
rect 23388 31962 23440 31968
rect 22744 31884 22796 31890
rect 22744 31826 22796 31832
rect 22652 31476 22704 31482
rect 22652 31418 22704 31424
rect 22756 31362 22784 31826
rect 22664 31346 22784 31362
rect 23492 31346 23520 32166
rect 23676 31822 23704 32166
rect 23664 31816 23716 31822
rect 23664 31758 23716 31764
rect 22652 31340 22784 31346
rect 22704 31334 22784 31340
rect 23480 31340 23532 31346
rect 22652 31282 22704 31288
rect 23480 31282 23532 31288
rect 22560 30660 22612 30666
rect 22560 30602 22612 30608
rect 22192 30592 22244 30598
rect 22192 30534 22244 30540
rect 21788 30492 22096 30501
rect 21788 30490 21794 30492
rect 21850 30490 21874 30492
rect 21930 30490 21954 30492
rect 22010 30490 22034 30492
rect 22090 30490 22096 30492
rect 21850 30438 21852 30490
rect 22032 30438 22034 30490
rect 21788 30436 21794 30438
rect 21850 30436 21874 30438
rect 21930 30436 21954 30438
rect 22010 30436 22034 30438
rect 22090 30436 22096 30438
rect 21788 30427 22096 30436
rect 21788 29404 22096 29413
rect 21788 29402 21794 29404
rect 21850 29402 21874 29404
rect 21930 29402 21954 29404
rect 22010 29402 22034 29404
rect 22090 29402 22096 29404
rect 21850 29350 21852 29402
rect 22032 29350 22034 29402
rect 21788 29348 21794 29350
rect 21850 29348 21874 29350
rect 21930 29348 21954 29350
rect 22010 29348 22034 29350
rect 22090 29348 22096 29350
rect 21788 29339 22096 29348
rect 22204 29186 22232 30534
rect 22376 30184 22428 30190
rect 22376 30126 22428 30132
rect 22112 29170 22232 29186
rect 22100 29164 22232 29170
rect 22152 29158 22232 29164
rect 22100 29106 22152 29112
rect 21640 29096 21692 29102
rect 21640 29038 21692 29044
rect 21548 28756 21600 28762
rect 21548 28698 21600 28704
rect 21456 27600 21508 27606
rect 21456 27542 21508 27548
rect 21364 27328 21416 27334
rect 21364 27270 21416 27276
rect 20996 26988 21048 26994
rect 20996 26930 21048 26936
rect 21180 26988 21232 26994
rect 21180 26930 21232 26936
rect 20904 25832 20956 25838
rect 20904 25774 20956 25780
rect 21008 25650 21036 26930
rect 21376 26450 21404 27270
rect 21468 26994 21496 27542
rect 21456 26988 21508 26994
rect 21560 26976 21588 28698
rect 22112 28626 22140 29106
rect 22284 28960 22336 28966
rect 22284 28902 22336 28908
rect 22100 28620 22152 28626
rect 22100 28562 22152 28568
rect 22112 28506 22140 28562
rect 22112 28478 22232 28506
rect 21788 28316 22096 28325
rect 21788 28314 21794 28316
rect 21850 28314 21874 28316
rect 21930 28314 21954 28316
rect 22010 28314 22034 28316
rect 22090 28314 22096 28316
rect 21850 28262 21852 28314
rect 22032 28262 22034 28314
rect 21788 28260 21794 28262
rect 21850 28260 21874 28262
rect 21930 28260 21954 28262
rect 22010 28260 22034 28262
rect 22090 28260 22096 28262
rect 21788 28251 22096 28260
rect 21788 27228 22096 27237
rect 21788 27226 21794 27228
rect 21850 27226 21874 27228
rect 21930 27226 21954 27228
rect 22010 27226 22034 27228
rect 22090 27226 22096 27228
rect 21850 27174 21852 27226
rect 22032 27174 22034 27226
rect 21788 27172 21794 27174
rect 21850 27172 21874 27174
rect 21930 27172 21954 27174
rect 22010 27172 22034 27174
rect 22090 27172 22096 27174
rect 21788 27163 22096 27172
rect 21560 26948 21680 26976
rect 21456 26930 21508 26936
rect 21548 26852 21600 26858
rect 21548 26794 21600 26800
rect 21364 26444 21416 26450
rect 21364 26386 21416 26392
rect 21272 26240 21324 26246
rect 21272 26182 21324 26188
rect 20916 25622 21036 25650
rect 20812 25492 20864 25498
rect 20812 25434 20864 25440
rect 20628 25356 20680 25362
rect 20628 25298 20680 25304
rect 20916 24886 20944 25622
rect 21284 25362 21312 26182
rect 21376 26042 21404 26386
rect 21560 26382 21588 26794
rect 21548 26376 21600 26382
rect 21548 26318 21600 26324
rect 21364 26036 21416 26042
rect 21364 25978 21416 25984
rect 21272 25356 21324 25362
rect 21272 25298 21324 25304
rect 20996 25288 21048 25294
rect 20996 25230 21048 25236
rect 20904 24880 20956 24886
rect 20904 24822 20956 24828
rect 20536 22772 20588 22778
rect 20536 22714 20588 22720
rect 20812 21344 20864 21350
rect 20812 21286 20864 21292
rect 20824 20942 20852 21286
rect 20812 20936 20864 20942
rect 20812 20878 20864 20884
rect 20260 19304 20312 19310
rect 20260 19246 20312 19252
rect 20272 18698 20300 19246
rect 20916 18698 20944 24822
rect 21008 23118 21036 25230
rect 21560 24206 21588 26318
rect 21652 26314 21680 26948
rect 21732 26784 21784 26790
rect 21732 26726 21784 26732
rect 21744 26382 21772 26726
rect 22204 26586 22232 28478
rect 22296 27062 22324 28902
rect 22388 27402 22416 30126
rect 22572 29238 22600 30602
rect 22664 30326 22692 31282
rect 22652 30320 22704 30326
rect 22652 30262 22704 30268
rect 22664 29714 22692 30262
rect 22652 29708 22704 29714
rect 22652 29650 22704 29656
rect 22836 29640 22888 29646
rect 22836 29582 22888 29588
rect 23940 29640 23992 29646
rect 23940 29582 23992 29588
rect 22848 29306 22876 29582
rect 23480 29572 23532 29578
rect 23480 29514 23532 29520
rect 22928 29504 22980 29510
rect 22928 29446 22980 29452
rect 22836 29300 22888 29306
rect 22836 29242 22888 29248
rect 22560 29232 22612 29238
rect 22560 29174 22612 29180
rect 22376 27396 22428 27402
rect 22376 27338 22428 27344
rect 22388 27146 22416 27338
rect 22388 27130 22508 27146
rect 22388 27124 22520 27130
rect 22388 27118 22468 27124
rect 22468 27066 22520 27072
rect 22284 27056 22336 27062
rect 22284 26998 22336 27004
rect 22192 26580 22244 26586
rect 22192 26522 22244 26528
rect 21732 26376 21784 26382
rect 21732 26318 21784 26324
rect 21640 26308 21692 26314
rect 21640 26250 21692 26256
rect 21652 24818 21680 26250
rect 21788 26140 22096 26149
rect 21788 26138 21794 26140
rect 21850 26138 21874 26140
rect 21930 26138 21954 26140
rect 22010 26138 22034 26140
rect 22090 26138 22096 26140
rect 21850 26086 21852 26138
rect 22032 26086 22034 26138
rect 21788 26084 21794 26086
rect 21850 26084 21874 26086
rect 21930 26084 21954 26086
rect 22010 26084 22034 26086
rect 22090 26084 22096 26086
rect 21788 26075 22096 26084
rect 22480 25362 22508 27066
rect 22572 25702 22600 29174
rect 22940 29170 22968 29446
rect 23492 29170 23520 29514
rect 22928 29164 22980 29170
rect 22928 29106 22980 29112
rect 23480 29164 23532 29170
rect 23480 29106 23532 29112
rect 23492 29034 23520 29106
rect 23480 29028 23532 29034
rect 23480 28970 23532 28976
rect 23388 28484 23440 28490
rect 23388 28426 23440 28432
rect 23400 28082 23428 28426
rect 23492 28082 23520 28970
rect 23664 28552 23716 28558
rect 23664 28494 23716 28500
rect 23848 28552 23900 28558
rect 23848 28494 23900 28500
rect 23388 28076 23440 28082
rect 23388 28018 23440 28024
rect 23480 28076 23532 28082
rect 23480 28018 23532 28024
rect 23020 27872 23072 27878
rect 23020 27814 23072 27820
rect 23032 27470 23060 27814
rect 23020 27464 23072 27470
rect 23020 27406 23072 27412
rect 22744 27056 22796 27062
rect 22744 26998 22796 27004
rect 22560 25696 22612 25702
rect 22560 25638 22612 25644
rect 22468 25356 22520 25362
rect 22468 25298 22520 25304
rect 22376 25288 22428 25294
rect 22376 25230 22428 25236
rect 21788 25052 22096 25061
rect 21788 25050 21794 25052
rect 21850 25050 21874 25052
rect 21930 25050 21954 25052
rect 22010 25050 22034 25052
rect 22090 25050 22096 25052
rect 21850 24998 21852 25050
rect 22032 24998 22034 25050
rect 21788 24996 21794 24998
rect 21850 24996 21874 24998
rect 21930 24996 21954 24998
rect 22010 24996 22034 24998
rect 22090 24996 22096 24998
rect 21788 24987 22096 24996
rect 22388 24954 22416 25230
rect 22376 24948 22428 24954
rect 22376 24890 22428 24896
rect 21640 24812 21692 24818
rect 21640 24754 21692 24760
rect 21824 24812 21876 24818
rect 21824 24754 21876 24760
rect 21548 24200 21600 24206
rect 21732 24200 21784 24206
rect 21548 24142 21600 24148
rect 21652 24148 21732 24154
rect 21652 24142 21784 24148
rect 21364 24132 21416 24138
rect 21364 24074 21416 24080
rect 21376 23798 21404 24074
rect 21456 24064 21508 24070
rect 21456 24006 21508 24012
rect 21364 23792 21416 23798
rect 21364 23734 21416 23740
rect 21180 23724 21232 23730
rect 21180 23666 21232 23672
rect 21192 23322 21220 23666
rect 21180 23316 21232 23322
rect 21180 23258 21232 23264
rect 20996 23112 21048 23118
rect 20996 23054 21048 23060
rect 21008 21554 21036 23054
rect 21272 22432 21324 22438
rect 21272 22374 21324 22380
rect 21180 21888 21232 21894
rect 21180 21830 21232 21836
rect 21088 21616 21140 21622
rect 21088 21558 21140 21564
rect 20996 21548 21048 21554
rect 20996 21490 21048 21496
rect 21100 21010 21128 21558
rect 21192 21554 21220 21830
rect 21180 21548 21232 21554
rect 21180 21490 21232 21496
rect 21284 21418 21312 22374
rect 21376 21894 21404 23734
rect 21468 23186 21496 24006
rect 21456 23180 21508 23186
rect 21456 23122 21508 23128
rect 21560 22094 21588 24142
rect 21652 24126 21772 24142
rect 21652 23662 21680 24126
rect 21836 24070 21864 24754
rect 21824 24064 21876 24070
rect 21824 24006 21876 24012
rect 21788 23964 22096 23973
rect 21788 23962 21794 23964
rect 21850 23962 21874 23964
rect 21930 23962 21954 23964
rect 22010 23962 22034 23964
rect 22090 23962 22096 23964
rect 21850 23910 21852 23962
rect 22032 23910 22034 23962
rect 21788 23908 21794 23910
rect 21850 23908 21874 23910
rect 21930 23908 21954 23910
rect 22010 23908 22034 23910
rect 22090 23908 22096 23910
rect 21788 23899 22096 23908
rect 22376 23792 22428 23798
rect 22376 23734 22428 23740
rect 21640 23656 21692 23662
rect 21640 23598 21692 23604
rect 21468 22066 21588 22094
rect 21468 22030 21496 22066
rect 21456 22024 21508 22030
rect 21456 21966 21508 21972
rect 21364 21888 21416 21894
rect 21364 21830 21416 21836
rect 21272 21412 21324 21418
rect 21272 21354 21324 21360
rect 21088 21004 21140 21010
rect 21088 20946 21140 20952
rect 21468 20466 21496 21966
rect 21652 21010 21680 23598
rect 22008 23520 22060 23526
rect 22008 23462 22060 23468
rect 22020 23322 22048 23462
rect 22008 23316 22060 23322
rect 22008 23258 22060 23264
rect 21788 22876 22096 22885
rect 21788 22874 21794 22876
rect 21850 22874 21874 22876
rect 21930 22874 21954 22876
rect 22010 22874 22034 22876
rect 22090 22874 22096 22876
rect 21850 22822 21852 22874
rect 22032 22822 22034 22874
rect 21788 22820 21794 22822
rect 21850 22820 21874 22822
rect 21930 22820 21954 22822
rect 22010 22820 22034 22822
rect 22090 22820 22096 22822
rect 21788 22811 22096 22820
rect 22388 22710 22416 23734
rect 22376 22704 22428 22710
rect 22376 22646 22428 22652
rect 22388 22234 22416 22646
rect 22376 22228 22428 22234
rect 22376 22170 22428 22176
rect 22284 21888 22336 21894
rect 22284 21830 22336 21836
rect 21788 21788 22096 21797
rect 21788 21786 21794 21788
rect 21850 21786 21874 21788
rect 21930 21786 21954 21788
rect 22010 21786 22034 21788
rect 22090 21786 22096 21788
rect 21850 21734 21852 21786
rect 22032 21734 22034 21786
rect 21788 21732 21794 21734
rect 21850 21732 21874 21734
rect 21930 21732 21954 21734
rect 22010 21732 22034 21734
rect 22090 21732 22096 21734
rect 21788 21723 22096 21732
rect 21640 21004 21692 21010
rect 21640 20946 21692 20952
rect 21456 20460 21508 20466
rect 21456 20402 21508 20408
rect 21180 19372 21232 19378
rect 21180 19314 21232 19320
rect 21088 19168 21140 19174
rect 21088 19110 21140 19116
rect 21100 18766 21128 19110
rect 21088 18760 21140 18766
rect 21088 18702 21140 18708
rect 20260 18692 20312 18698
rect 20260 18634 20312 18640
rect 20904 18692 20956 18698
rect 20904 18634 20956 18640
rect 20168 17740 20220 17746
rect 20168 17682 20220 17688
rect 20272 17542 20300 18634
rect 20812 18624 20864 18630
rect 20812 18566 20864 18572
rect 20076 17536 20128 17542
rect 20076 17478 20128 17484
rect 20260 17536 20312 17542
rect 20260 17478 20312 17484
rect 20088 17338 20116 17478
rect 20076 17332 20128 17338
rect 20076 17274 20128 17280
rect 19984 17128 20036 17134
rect 19984 17070 20036 17076
rect 20444 17128 20496 17134
rect 20444 17070 20496 17076
rect 20456 15162 20484 17070
rect 20536 16992 20588 16998
rect 20536 16934 20588 16940
rect 20444 15156 20496 15162
rect 20444 15098 20496 15104
rect 20352 15020 20404 15026
rect 20352 14962 20404 14968
rect 20364 14074 20392 14962
rect 20352 14068 20404 14074
rect 20352 14010 20404 14016
rect 19616 13932 19668 13938
rect 19616 13874 19668 13880
rect 19892 13932 19944 13938
rect 19892 13874 19944 13880
rect 20444 13932 20496 13938
rect 20444 13874 20496 13880
rect 19628 13530 19656 13874
rect 19616 13524 19668 13530
rect 19616 13466 19668 13472
rect 19904 12850 19932 13874
rect 20456 12986 20484 13874
rect 20444 12980 20496 12986
rect 20444 12922 20496 12928
rect 19892 12844 19944 12850
rect 19892 12786 19944 12792
rect 20168 12844 20220 12850
rect 20168 12786 20220 12792
rect 20180 12306 20208 12786
rect 20260 12640 20312 12646
rect 20260 12582 20312 12588
rect 20168 12300 20220 12306
rect 20168 12242 20220 12248
rect 19156 11348 19208 11354
rect 19156 11290 19208 11296
rect 19248 11008 19300 11014
rect 19248 10950 19300 10956
rect 18892 10674 19012 10690
rect 19260 10674 19288 10950
rect 20272 10674 20300 12582
rect 18880 10668 19012 10674
rect 18932 10662 19012 10668
rect 19156 10668 19208 10674
rect 18880 10610 18932 10616
rect 19156 10610 19208 10616
rect 19248 10668 19300 10674
rect 19248 10610 19300 10616
rect 20260 10668 20312 10674
rect 20260 10610 20312 10616
rect 18248 10526 18368 10554
rect 18144 10464 18196 10470
rect 18144 10406 18196 10412
rect 18156 10130 18184 10406
rect 18248 10266 18276 10526
rect 18315 10364 18623 10373
rect 18315 10362 18321 10364
rect 18377 10362 18401 10364
rect 18457 10362 18481 10364
rect 18537 10362 18561 10364
rect 18617 10362 18623 10364
rect 18377 10310 18379 10362
rect 18559 10310 18561 10362
rect 18315 10308 18321 10310
rect 18377 10308 18401 10310
rect 18457 10308 18481 10310
rect 18537 10308 18561 10310
rect 18617 10308 18623 10310
rect 18315 10299 18623 10308
rect 18236 10260 18288 10266
rect 18236 10202 18288 10208
rect 18144 10124 18196 10130
rect 18144 10066 18196 10072
rect 18892 9994 18920 10610
rect 19168 10198 19196 10610
rect 20168 10600 20220 10606
rect 20168 10542 20220 10548
rect 19156 10192 19208 10198
rect 19156 10134 19208 10140
rect 20180 10062 20208 10542
rect 20272 10130 20300 10610
rect 20260 10124 20312 10130
rect 20260 10066 20312 10072
rect 20168 10056 20220 10062
rect 20168 9998 20220 10004
rect 18880 9988 18932 9994
rect 18880 9930 18932 9936
rect 20548 9586 20576 16934
rect 20720 16516 20772 16522
rect 20720 16458 20772 16464
rect 20732 16250 20760 16458
rect 20720 16244 20772 16250
rect 20720 16186 20772 16192
rect 20824 15706 20852 18566
rect 21192 18426 21220 19314
rect 21180 18420 21232 18426
rect 21180 18362 21232 18368
rect 20904 18216 20956 18222
rect 20904 18158 20956 18164
rect 20916 17678 20944 18158
rect 21652 17882 21680 20946
rect 22296 20754 22324 21830
rect 22376 21344 22428 21350
rect 22376 21286 22428 21292
rect 22388 20942 22416 21286
rect 22376 20936 22428 20942
rect 22376 20878 22428 20884
rect 22468 20800 22520 20806
rect 22296 20726 22416 20754
rect 22468 20742 22520 20748
rect 21788 20700 22096 20709
rect 21788 20698 21794 20700
rect 21850 20698 21874 20700
rect 21930 20698 21954 20700
rect 22010 20698 22034 20700
rect 22090 20698 22096 20700
rect 21850 20646 21852 20698
rect 22032 20646 22034 20698
rect 21788 20644 21794 20646
rect 21850 20644 21874 20646
rect 21930 20644 21954 20646
rect 22010 20644 22034 20646
rect 22090 20644 22096 20646
rect 21788 20635 22096 20644
rect 22388 20466 22416 20726
rect 22376 20460 22428 20466
rect 22376 20402 22428 20408
rect 21788 19612 22096 19621
rect 21788 19610 21794 19612
rect 21850 19610 21874 19612
rect 21930 19610 21954 19612
rect 22010 19610 22034 19612
rect 22090 19610 22096 19612
rect 21850 19558 21852 19610
rect 22032 19558 22034 19610
rect 21788 19556 21794 19558
rect 21850 19556 21874 19558
rect 21930 19556 21954 19558
rect 22010 19556 22034 19558
rect 22090 19556 22096 19558
rect 21788 19547 22096 19556
rect 22388 18766 22416 20402
rect 22480 20398 22508 20742
rect 22468 20392 22520 20398
rect 22468 20334 22520 20340
rect 22376 18760 22428 18766
rect 22376 18702 22428 18708
rect 22192 18624 22244 18630
rect 22192 18566 22244 18572
rect 21788 18524 22096 18533
rect 21788 18522 21794 18524
rect 21850 18522 21874 18524
rect 21930 18522 21954 18524
rect 22010 18522 22034 18524
rect 22090 18522 22096 18524
rect 21850 18470 21852 18522
rect 22032 18470 22034 18522
rect 21788 18468 21794 18470
rect 21850 18468 21874 18470
rect 21930 18468 21954 18470
rect 22010 18468 22034 18470
rect 22090 18468 22096 18470
rect 21788 18459 22096 18468
rect 22204 18426 22232 18566
rect 22480 18426 22508 20334
rect 22192 18420 22244 18426
rect 22192 18362 22244 18368
rect 22468 18420 22520 18426
rect 22468 18362 22520 18368
rect 21640 17876 21692 17882
rect 21640 17818 21692 17824
rect 20904 17672 20956 17678
rect 20904 17614 20956 17620
rect 21652 17202 21680 17818
rect 21788 17436 22096 17445
rect 21788 17434 21794 17436
rect 21850 17434 21874 17436
rect 21930 17434 21954 17436
rect 22010 17434 22034 17436
rect 22090 17434 22096 17436
rect 21850 17382 21852 17434
rect 22032 17382 22034 17434
rect 21788 17380 21794 17382
rect 21850 17380 21874 17382
rect 21930 17380 21954 17382
rect 22010 17380 22034 17382
rect 22090 17380 22096 17382
rect 21788 17371 22096 17380
rect 22204 17270 22232 18362
rect 22572 18358 22600 25638
rect 22756 24886 22784 26998
rect 22744 24880 22796 24886
rect 22744 24822 22796 24828
rect 22756 24410 22784 24822
rect 22744 24404 22796 24410
rect 22744 24346 22796 24352
rect 22756 23798 22784 24346
rect 22836 24132 22888 24138
rect 22836 24074 22888 24080
rect 22848 23866 22876 24074
rect 22836 23860 22888 23866
rect 22836 23802 22888 23808
rect 22744 23792 22796 23798
rect 22744 23734 22796 23740
rect 22744 21888 22796 21894
rect 22744 21830 22796 21836
rect 22756 21554 22784 21830
rect 22744 21548 22796 21554
rect 22744 21490 22796 21496
rect 22836 21480 22888 21486
rect 22836 21422 22888 21428
rect 22848 20602 22876 21422
rect 22836 20596 22888 20602
rect 22836 20538 22888 20544
rect 23032 18630 23060 27406
rect 23400 26586 23428 28018
rect 23676 27946 23704 28494
rect 23664 27940 23716 27946
rect 23664 27882 23716 27888
rect 23860 27470 23888 28494
rect 23848 27464 23900 27470
rect 23848 27406 23900 27412
rect 23388 26580 23440 26586
rect 23388 26522 23440 26528
rect 23400 25838 23428 26522
rect 23860 26042 23888 27406
rect 23952 27334 23980 29582
rect 24032 29096 24084 29102
rect 24032 29038 24084 29044
rect 24044 27470 24072 29038
rect 24032 27464 24084 27470
rect 24032 27406 24084 27412
rect 23940 27328 23992 27334
rect 23940 27270 23992 27276
rect 23848 26036 23900 26042
rect 23848 25978 23900 25984
rect 23388 25832 23440 25838
rect 23388 25774 23440 25780
rect 23400 25498 23428 25774
rect 23388 25492 23440 25498
rect 23388 25434 23440 25440
rect 23400 24886 23428 25434
rect 23848 25152 23900 25158
rect 23848 25094 23900 25100
rect 23388 24880 23440 24886
rect 23388 24822 23440 24828
rect 23756 24812 23808 24818
rect 23756 24754 23808 24760
rect 23572 24676 23624 24682
rect 23572 24618 23624 24624
rect 23296 24608 23348 24614
rect 23296 24550 23348 24556
rect 23584 24562 23612 24618
rect 23308 23730 23336 24550
rect 23584 24534 23704 24562
rect 23296 23724 23348 23730
rect 23296 23666 23348 23672
rect 23676 23594 23704 24534
rect 23768 24070 23796 24754
rect 23756 24064 23808 24070
rect 23756 24006 23808 24012
rect 23664 23588 23716 23594
rect 23664 23530 23716 23536
rect 23676 22642 23704 23530
rect 23664 22636 23716 22642
rect 23664 22578 23716 22584
rect 23676 22030 23704 22578
rect 23664 22024 23716 22030
rect 23664 21966 23716 21972
rect 23676 20534 23704 21966
rect 23756 21888 23808 21894
rect 23756 21830 23808 21836
rect 23664 20528 23716 20534
rect 23664 20470 23716 20476
rect 23768 18766 23796 21830
rect 23388 18760 23440 18766
rect 23388 18702 23440 18708
rect 23756 18760 23808 18766
rect 23756 18702 23808 18708
rect 23112 18692 23164 18698
rect 23112 18634 23164 18640
rect 23296 18692 23348 18698
rect 23296 18634 23348 18640
rect 23020 18624 23072 18630
rect 23020 18566 23072 18572
rect 23020 18420 23072 18426
rect 23020 18362 23072 18368
rect 22560 18352 22612 18358
rect 22560 18294 22612 18300
rect 22572 17678 22600 18294
rect 22560 17672 22612 17678
rect 22560 17614 22612 17620
rect 22652 17536 22704 17542
rect 22652 17478 22704 17484
rect 22664 17270 22692 17478
rect 23032 17338 23060 18362
rect 23124 18358 23152 18634
rect 23112 18352 23164 18358
rect 23112 18294 23164 18300
rect 23308 18222 23336 18634
rect 23296 18216 23348 18222
rect 23296 18158 23348 18164
rect 23204 18080 23256 18086
rect 23204 18022 23256 18028
rect 23112 17876 23164 17882
rect 23112 17818 23164 17824
rect 23124 17678 23152 17818
rect 23216 17746 23244 18022
rect 23204 17740 23256 17746
rect 23204 17682 23256 17688
rect 23112 17672 23164 17678
rect 23112 17614 23164 17620
rect 23308 17626 23336 18158
rect 23400 17746 23428 18702
rect 23572 18624 23624 18630
rect 23572 18566 23624 18572
rect 23388 17740 23440 17746
rect 23388 17682 23440 17688
rect 23308 17610 23428 17626
rect 23308 17604 23440 17610
rect 23308 17598 23388 17604
rect 23020 17332 23072 17338
rect 23020 17274 23072 17280
rect 22192 17264 22244 17270
rect 22192 17206 22244 17212
rect 22560 17264 22612 17270
rect 22560 17206 22612 17212
rect 22652 17264 22704 17270
rect 22652 17206 22704 17212
rect 21640 17196 21692 17202
rect 21640 17138 21692 17144
rect 21456 16584 21508 16590
rect 21456 16526 21508 16532
rect 21468 16114 21496 16526
rect 21272 16108 21324 16114
rect 21272 16050 21324 16056
rect 21456 16108 21508 16114
rect 21456 16050 21508 16056
rect 20812 15700 20864 15706
rect 20812 15642 20864 15648
rect 20628 15156 20680 15162
rect 20628 15098 20680 15104
rect 20640 13394 20668 15098
rect 20628 13388 20680 13394
rect 20628 13330 20680 13336
rect 20824 13326 20852 15642
rect 21284 15162 21312 16050
rect 21652 15570 21680 17138
rect 22572 16454 22600 17206
rect 23032 16590 23060 17274
rect 23020 16584 23072 16590
rect 23020 16526 23072 16532
rect 22560 16448 22612 16454
rect 22560 16390 22612 16396
rect 21788 16348 22096 16357
rect 21788 16346 21794 16348
rect 21850 16346 21874 16348
rect 21930 16346 21954 16348
rect 22010 16346 22034 16348
rect 22090 16346 22096 16348
rect 21850 16294 21852 16346
rect 22032 16294 22034 16346
rect 21788 16292 21794 16294
rect 21850 16292 21874 16294
rect 21930 16292 21954 16294
rect 22010 16292 22034 16294
rect 22090 16292 22096 16294
rect 21788 16283 22096 16292
rect 21640 15564 21692 15570
rect 21640 15506 21692 15512
rect 21548 15428 21600 15434
rect 21548 15370 21600 15376
rect 21272 15156 21324 15162
rect 21272 15098 21324 15104
rect 21456 14816 21508 14822
rect 21456 14758 21508 14764
rect 21468 13326 21496 14758
rect 20812 13320 20864 13326
rect 20812 13262 20864 13268
rect 21456 13320 21508 13326
rect 21456 13262 21508 13268
rect 21088 13184 21140 13190
rect 21088 13126 21140 13132
rect 21100 12850 21128 13126
rect 21088 12844 21140 12850
rect 21088 12786 21140 12792
rect 21560 12442 21588 15370
rect 21788 15260 22096 15269
rect 21788 15258 21794 15260
rect 21850 15258 21874 15260
rect 21930 15258 21954 15260
rect 22010 15258 22034 15260
rect 22090 15258 22096 15260
rect 21850 15206 21852 15258
rect 22032 15206 22034 15258
rect 21788 15204 21794 15206
rect 21850 15204 21874 15206
rect 21930 15204 21954 15206
rect 22010 15204 22034 15206
rect 22090 15204 22096 15206
rect 21788 15195 22096 15204
rect 22572 15162 22600 16390
rect 23032 15450 23060 16526
rect 23032 15422 23152 15450
rect 23020 15360 23072 15366
rect 23020 15302 23072 15308
rect 22560 15156 22612 15162
rect 22560 15098 22612 15104
rect 22744 14884 22796 14890
rect 22744 14826 22796 14832
rect 21788 14172 22096 14181
rect 21788 14170 21794 14172
rect 21850 14170 21874 14172
rect 21930 14170 21954 14172
rect 22010 14170 22034 14172
rect 22090 14170 22096 14172
rect 21850 14118 21852 14170
rect 22032 14118 22034 14170
rect 21788 14116 21794 14118
rect 21850 14116 21874 14118
rect 21930 14116 21954 14118
rect 22010 14116 22034 14118
rect 22090 14116 22096 14118
rect 21788 14107 22096 14116
rect 22756 14074 22784 14826
rect 22744 14068 22796 14074
rect 22744 14010 22796 14016
rect 21640 13864 21692 13870
rect 21640 13806 21692 13812
rect 22468 13864 22520 13870
rect 22468 13806 22520 13812
rect 21548 12436 21600 12442
rect 21548 12378 21600 12384
rect 21652 12238 21680 13806
rect 22284 13796 22336 13802
rect 22284 13738 22336 13744
rect 22296 13530 22324 13738
rect 22284 13524 22336 13530
rect 22284 13466 22336 13472
rect 21788 13084 22096 13093
rect 21788 13082 21794 13084
rect 21850 13082 21874 13084
rect 21930 13082 21954 13084
rect 22010 13082 22034 13084
rect 22090 13082 22096 13084
rect 21850 13030 21852 13082
rect 22032 13030 22034 13082
rect 21788 13028 21794 13030
rect 21850 13028 21874 13030
rect 21930 13028 21954 13030
rect 22010 13028 22034 13030
rect 22090 13028 22096 13030
rect 21788 13019 22096 13028
rect 22480 12986 22508 13806
rect 22756 13190 22784 14010
rect 23032 14006 23060 15302
rect 23124 15162 23152 15422
rect 23112 15156 23164 15162
rect 23112 15098 23164 15104
rect 23020 14000 23072 14006
rect 23020 13942 23072 13948
rect 23032 13394 23060 13942
rect 23124 13734 23152 15098
rect 23308 14890 23336 17598
rect 23388 17546 23440 17552
rect 23480 17536 23532 17542
rect 23480 17478 23532 17484
rect 23492 16590 23520 17478
rect 23480 16584 23532 16590
rect 23480 16526 23532 16532
rect 23296 14884 23348 14890
rect 23296 14826 23348 14832
rect 23480 14068 23532 14074
rect 23480 14010 23532 14016
rect 23112 13728 23164 13734
rect 23112 13670 23164 13676
rect 23296 13728 23348 13734
rect 23296 13670 23348 13676
rect 23020 13388 23072 13394
rect 23020 13330 23072 13336
rect 23124 13258 23152 13670
rect 23308 13530 23336 13670
rect 23296 13524 23348 13530
rect 23296 13466 23348 13472
rect 23112 13252 23164 13258
rect 23112 13194 23164 13200
rect 22744 13184 22796 13190
rect 22744 13126 22796 13132
rect 22836 13184 22888 13190
rect 22836 13126 22888 13132
rect 22468 12980 22520 12986
rect 22468 12922 22520 12928
rect 22848 12866 22876 13126
rect 23308 12918 23336 13466
rect 23492 13258 23520 14010
rect 23584 13326 23612 18566
rect 23860 17882 23888 25094
rect 23952 23662 23980 27270
rect 24044 25702 24072 27406
rect 24032 25696 24084 25702
rect 24032 25638 24084 25644
rect 23940 23656 23992 23662
rect 23940 23598 23992 23604
rect 24032 22772 24084 22778
rect 24032 22714 24084 22720
rect 23940 22500 23992 22506
rect 23940 22442 23992 22448
rect 23952 21962 23980 22442
rect 23940 21956 23992 21962
rect 23940 21898 23992 21904
rect 23952 20466 23980 21898
rect 23940 20460 23992 20466
rect 23940 20402 23992 20408
rect 23940 19916 23992 19922
rect 23940 19858 23992 19864
rect 23952 18154 23980 19858
rect 23940 18148 23992 18154
rect 23940 18090 23992 18096
rect 23848 17876 23900 17882
rect 23768 17836 23848 17864
rect 23664 16448 23716 16454
rect 23664 16390 23716 16396
rect 23676 15094 23704 16390
rect 23664 15088 23716 15094
rect 23664 15030 23716 15036
rect 23768 14074 23796 17836
rect 23848 17818 23900 17824
rect 23848 17672 23900 17678
rect 23848 17614 23900 17620
rect 23860 16658 23888 17614
rect 23848 16652 23900 16658
rect 23848 16594 23900 16600
rect 23756 14068 23808 14074
rect 23756 14010 23808 14016
rect 23756 13932 23808 13938
rect 23756 13874 23808 13880
rect 23664 13864 23716 13870
rect 23664 13806 23716 13812
rect 23676 13462 23704 13806
rect 23664 13456 23716 13462
rect 23664 13398 23716 13404
rect 23572 13320 23624 13326
rect 23572 13262 23624 13268
rect 23480 13252 23532 13258
rect 23480 13194 23532 13200
rect 22756 12838 22876 12866
rect 23296 12912 23348 12918
rect 23296 12854 23348 12860
rect 23492 12850 23520 13194
rect 23768 12986 23796 13874
rect 23756 12980 23808 12986
rect 23756 12922 23808 12928
rect 23480 12844 23532 12850
rect 22756 12782 22784 12838
rect 23480 12786 23532 12792
rect 23860 12782 23888 16594
rect 23952 12918 23980 18090
rect 24044 17882 24072 22714
rect 24032 17876 24084 17882
rect 24032 17818 24084 17824
rect 24044 14074 24072 17818
rect 24136 17338 24164 34954
rect 24504 32366 24532 36178
rect 24688 33998 24716 36518
rect 24780 36242 24808 36518
rect 24768 36236 24820 36242
rect 24768 36178 24820 36184
rect 24872 35766 24900 36722
rect 25261 36476 25569 36485
rect 25261 36474 25267 36476
rect 25323 36474 25347 36476
rect 25403 36474 25427 36476
rect 25483 36474 25507 36476
rect 25563 36474 25569 36476
rect 25323 36422 25325 36474
rect 25505 36422 25507 36474
rect 25261 36420 25267 36422
rect 25323 36420 25347 36422
rect 25403 36420 25427 36422
rect 25483 36420 25507 36422
rect 25563 36420 25569 36422
rect 25261 36411 25569 36420
rect 25780 36168 25832 36174
rect 25780 36110 25832 36116
rect 25688 36032 25740 36038
rect 25688 35974 25740 35980
rect 24860 35760 24912 35766
rect 24860 35702 24912 35708
rect 24768 35692 24820 35698
rect 24768 35634 24820 35640
rect 24780 35290 24808 35634
rect 24768 35284 24820 35290
rect 24768 35226 24820 35232
rect 24872 34610 24900 35702
rect 25261 35388 25569 35397
rect 25261 35386 25267 35388
rect 25323 35386 25347 35388
rect 25403 35386 25427 35388
rect 25483 35386 25507 35388
rect 25563 35386 25569 35388
rect 25323 35334 25325 35386
rect 25505 35334 25507 35386
rect 25261 35332 25267 35334
rect 25323 35332 25347 35334
rect 25403 35332 25427 35334
rect 25483 35332 25507 35334
rect 25563 35332 25569 35334
rect 25261 35323 25569 35332
rect 24952 35080 25004 35086
rect 24952 35022 25004 35028
rect 24964 34678 24992 35022
rect 25700 34678 25728 35974
rect 25792 35290 25820 36110
rect 25780 35284 25832 35290
rect 25780 35226 25832 35232
rect 25976 35154 26004 44882
rect 26068 44334 26096 46271
rect 26056 44328 26108 44334
rect 26056 44270 26108 44276
rect 26160 43858 26188 46951
rect 26700 46922 26752 46928
rect 26712 46646 26740 46922
rect 26700 46640 26752 46646
rect 26700 46582 26752 46588
rect 26700 46436 26752 46442
rect 26700 46378 26752 46384
rect 26424 46368 26476 46374
rect 26424 46310 26476 46316
rect 26436 45558 26464 46310
rect 26240 45552 26292 45558
rect 26240 45494 26292 45500
rect 26424 45552 26476 45558
rect 26424 45494 26476 45500
rect 26252 45082 26280 45494
rect 26712 45490 26740 46378
rect 27080 46034 27108 49200
rect 27436 47048 27488 47054
rect 27436 46990 27488 46996
rect 27160 46572 27212 46578
rect 27160 46514 27212 46520
rect 27068 46028 27120 46034
rect 27068 45970 27120 45976
rect 26700 45484 26752 45490
rect 26700 45426 26752 45432
rect 27172 45354 27200 46514
rect 27344 46164 27396 46170
rect 27344 46106 27396 46112
rect 27252 45892 27304 45898
rect 27252 45834 27304 45840
rect 27264 45626 27292 45834
rect 27252 45620 27304 45626
rect 27252 45562 27304 45568
rect 27356 45490 27384 46106
rect 27448 46034 27476 46990
rect 27620 46640 27672 46646
rect 27620 46582 27672 46588
rect 27436 46028 27488 46034
rect 27436 45970 27488 45976
rect 27528 45960 27580 45966
rect 27528 45902 27580 45908
rect 27344 45484 27396 45490
rect 27344 45426 27396 45432
rect 27160 45348 27212 45354
rect 27160 45290 27212 45296
rect 26424 45280 26476 45286
rect 26424 45222 26476 45228
rect 26240 45076 26292 45082
rect 26240 45018 26292 45024
rect 26436 44470 26464 45222
rect 27252 44804 27304 44810
rect 27252 44746 27304 44752
rect 27264 44538 27292 44746
rect 27252 44532 27304 44538
rect 27252 44474 27304 44480
rect 26424 44464 26476 44470
rect 26424 44406 26476 44412
rect 27356 44402 27384 45426
rect 26884 44396 26936 44402
rect 26884 44338 26936 44344
rect 27344 44396 27396 44402
rect 27344 44338 27396 44344
rect 26148 43852 26200 43858
rect 26148 43794 26200 43800
rect 26056 43716 26108 43722
rect 26056 43658 26108 43664
rect 26068 43450 26096 43658
rect 26056 43444 26108 43450
rect 26056 43386 26108 43392
rect 26424 43104 26476 43110
rect 26424 43046 26476 43052
rect 26054 42936 26110 42945
rect 26054 42871 26110 42880
rect 26068 42158 26096 42871
rect 26148 42628 26200 42634
rect 26148 42570 26200 42576
rect 26056 42152 26108 42158
rect 26056 42094 26108 42100
rect 26160 41585 26188 42570
rect 26436 42294 26464 43046
rect 26424 42288 26476 42294
rect 26424 42230 26476 42236
rect 26146 41576 26202 41585
rect 26146 41511 26202 41520
rect 26516 40928 26568 40934
rect 26516 40870 26568 40876
rect 26528 40594 26556 40870
rect 26516 40588 26568 40594
rect 26516 40530 26568 40536
rect 26700 40452 26752 40458
rect 26700 40394 26752 40400
rect 26424 39364 26476 39370
rect 26424 39306 26476 39312
rect 26332 39296 26384 39302
rect 26332 39238 26384 39244
rect 26344 38962 26372 39238
rect 26332 38956 26384 38962
rect 26332 38898 26384 38904
rect 26436 38554 26464 39306
rect 26712 39098 26740 40394
rect 26700 39092 26752 39098
rect 26700 39034 26752 39040
rect 26516 38820 26568 38826
rect 26516 38762 26568 38768
rect 26424 38548 26476 38554
rect 26424 38490 26476 38496
rect 26528 38418 26556 38762
rect 26700 38752 26752 38758
rect 26700 38694 26752 38700
rect 26606 38448 26662 38457
rect 26516 38412 26568 38418
rect 26712 38418 26740 38694
rect 26606 38383 26662 38392
rect 26700 38412 26752 38418
rect 26516 38354 26568 38360
rect 26148 37188 26200 37194
rect 26148 37130 26200 37136
rect 26160 36145 26188 37130
rect 26146 36136 26202 36145
rect 26146 36071 26202 36080
rect 26240 36100 26292 36106
rect 26240 36042 26292 36048
rect 26252 35834 26280 36042
rect 26620 35894 26648 38383
rect 26700 38354 26752 38360
rect 26896 38282 26924 44338
rect 27540 44334 27568 45902
rect 27528 44328 27580 44334
rect 27528 44270 27580 44276
rect 27252 43784 27304 43790
rect 27252 43726 27304 43732
rect 27068 43308 27120 43314
rect 27068 43250 27120 43256
rect 26976 43240 27028 43246
rect 26976 43182 27028 43188
rect 26988 39982 27016 43182
rect 26976 39976 27028 39982
rect 26976 39918 27028 39924
rect 26884 38276 26936 38282
rect 26884 38218 26936 38224
rect 26620 35866 26832 35894
rect 26240 35828 26292 35834
rect 26240 35770 26292 35776
rect 26700 35692 26752 35698
rect 26700 35634 26752 35640
rect 26240 35488 26292 35494
rect 26240 35430 26292 35436
rect 26516 35488 26568 35494
rect 26516 35430 26568 35436
rect 25964 35148 26016 35154
rect 25964 35090 26016 35096
rect 24952 34672 25004 34678
rect 24952 34614 25004 34620
rect 25688 34672 25740 34678
rect 25688 34614 25740 34620
rect 24860 34604 24912 34610
rect 24860 34546 24912 34552
rect 24676 33992 24728 33998
rect 24676 33934 24728 33940
rect 24688 33046 24716 33934
rect 24872 33590 24900 34546
rect 25261 34300 25569 34309
rect 25261 34298 25267 34300
rect 25323 34298 25347 34300
rect 25403 34298 25427 34300
rect 25483 34298 25507 34300
rect 25563 34298 25569 34300
rect 25323 34246 25325 34298
rect 25505 34246 25507 34298
rect 25261 34244 25267 34246
rect 25323 34244 25347 34246
rect 25403 34244 25427 34246
rect 25483 34244 25507 34246
rect 25563 34244 25569 34246
rect 25261 34235 25569 34244
rect 26148 34128 26200 34134
rect 26148 34070 26200 34076
rect 24952 33856 25004 33862
rect 24952 33798 25004 33804
rect 24860 33584 24912 33590
rect 24860 33526 24912 33532
rect 24676 33040 24728 33046
rect 24676 32982 24728 32988
rect 24688 32858 24716 32982
rect 24596 32830 24716 32858
rect 24860 32904 24912 32910
rect 24964 32892 24992 33798
rect 25044 33312 25096 33318
rect 25044 33254 25096 33260
rect 25056 32910 25084 33254
rect 25261 33212 25569 33221
rect 25261 33210 25267 33212
rect 25323 33210 25347 33212
rect 25403 33210 25427 33212
rect 25483 33210 25507 33212
rect 25563 33210 25569 33212
rect 25323 33158 25325 33210
rect 25505 33158 25507 33210
rect 25261 33156 25267 33158
rect 25323 33156 25347 33158
rect 25403 33156 25427 33158
rect 25483 33156 25507 33158
rect 25563 33156 25569 33158
rect 25261 33147 25569 33156
rect 25136 32972 25188 32978
rect 25136 32914 25188 32920
rect 24912 32864 24992 32892
rect 25044 32904 25096 32910
rect 24860 32846 24912 32852
rect 25044 32846 25096 32852
rect 24492 32360 24544 32366
rect 24492 32302 24544 32308
rect 24400 31340 24452 31346
rect 24400 31282 24452 31288
rect 24412 30666 24440 31282
rect 24492 31272 24544 31278
rect 24492 31214 24544 31220
rect 24400 30660 24452 30666
rect 24400 30602 24452 30608
rect 24412 28490 24440 30602
rect 24400 28484 24452 28490
rect 24400 28426 24452 28432
rect 24504 28218 24532 31214
rect 24596 30190 24624 32830
rect 24676 32768 24728 32774
rect 24676 32710 24728 32716
rect 24584 30184 24636 30190
rect 24584 30126 24636 30132
rect 24584 29164 24636 29170
rect 24584 29106 24636 29112
rect 24596 28762 24624 29106
rect 24584 28756 24636 28762
rect 24584 28698 24636 28704
rect 24688 28558 24716 32710
rect 25148 31906 25176 32914
rect 25261 32124 25569 32133
rect 25261 32122 25267 32124
rect 25323 32122 25347 32124
rect 25403 32122 25427 32124
rect 25483 32122 25507 32124
rect 25563 32122 25569 32124
rect 25323 32070 25325 32122
rect 25505 32070 25507 32122
rect 25261 32068 25267 32070
rect 25323 32068 25347 32070
rect 25403 32068 25427 32070
rect 25483 32068 25507 32070
rect 25563 32068 25569 32070
rect 25261 32059 25569 32068
rect 25056 31878 25176 31906
rect 25872 31952 25924 31958
rect 25872 31894 25924 31900
rect 25056 31482 25084 31878
rect 25136 31816 25188 31822
rect 25136 31758 25188 31764
rect 25044 31476 25096 31482
rect 25044 31418 25096 31424
rect 25056 30734 25084 31418
rect 25148 30938 25176 31758
rect 25596 31748 25648 31754
rect 25596 31690 25648 31696
rect 25608 31414 25636 31690
rect 25596 31408 25648 31414
rect 25596 31350 25648 31356
rect 25608 31142 25636 31350
rect 25596 31136 25648 31142
rect 25596 31078 25648 31084
rect 25261 31036 25569 31045
rect 25261 31034 25267 31036
rect 25323 31034 25347 31036
rect 25403 31034 25427 31036
rect 25483 31034 25507 31036
rect 25563 31034 25569 31036
rect 25323 30982 25325 31034
rect 25505 30982 25507 31034
rect 25261 30980 25267 30982
rect 25323 30980 25347 30982
rect 25403 30980 25427 30982
rect 25483 30980 25507 30982
rect 25563 30980 25569 30982
rect 25261 30971 25569 30980
rect 25136 30932 25188 30938
rect 25136 30874 25188 30880
rect 24860 30728 24912 30734
rect 24860 30670 24912 30676
rect 25044 30728 25096 30734
rect 25044 30670 25096 30676
rect 24872 29578 24900 30670
rect 25261 29948 25569 29957
rect 25261 29946 25267 29948
rect 25323 29946 25347 29948
rect 25403 29946 25427 29948
rect 25483 29946 25507 29948
rect 25563 29946 25569 29948
rect 25323 29894 25325 29946
rect 25505 29894 25507 29946
rect 25261 29892 25267 29894
rect 25323 29892 25347 29894
rect 25403 29892 25427 29894
rect 25483 29892 25507 29894
rect 25563 29892 25569 29894
rect 25261 29883 25569 29892
rect 25608 29850 25636 31078
rect 25884 30734 25912 31894
rect 26160 31385 26188 34070
rect 26252 33862 26280 35430
rect 26528 35154 26556 35430
rect 26516 35148 26568 35154
rect 26516 35090 26568 35096
rect 26608 34740 26660 34746
rect 26608 34682 26660 34688
rect 26620 34066 26648 34682
rect 26608 34060 26660 34066
rect 26608 34002 26660 34008
rect 26240 33856 26292 33862
rect 26240 33798 26292 33804
rect 26712 33386 26740 35634
rect 26700 33380 26752 33386
rect 26700 33322 26752 33328
rect 26516 32904 26568 32910
rect 26516 32846 26568 32852
rect 26424 32496 26476 32502
rect 26424 32438 26476 32444
rect 26332 31816 26384 31822
rect 26332 31758 26384 31764
rect 26146 31376 26202 31385
rect 26056 31340 26108 31346
rect 26146 31311 26202 31320
rect 26056 31282 26108 31288
rect 25964 31136 26016 31142
rect 25964 31078 26016 31084
rect 25872 30728 25924 30734
rect 25872 30670 25924 30676
rect 25780 30660 25832 30666
rect 25780 30602 25832 30608
rect 25596 29844 25648 29850
rect 25596 29786 25648 29792
rect 24860 29572 24912 29578
rect 24860 29514 24912 29520
rect 24952 29504 25004 29510
rect 24952 29446 25004 29452
rect 24964 29238 24992 29446
rect 24952 29232 25004 29238
rect 24952 29174 25004 29180
rect 25136 29096 25188 29102
rect 24766 29064 24822 29073
rect 25136 29038 25188 29044
rect 24766 28999 24822 29008
rect 24676 28552 24728 28558
rect 24676 28494 24728 28500
rect 24492 28212 24544 28218
rect 24492 28154 24544 28160
rect 24504 26382 24532 28154
rect 24492 26376 24544 26382
rect 24492 26318 24544 26324
rect 24504 25294 24532 26318
rect 24676 26240 24728 26246
rect 24676 26182 24728 26188
rect 24584 26036 24636 26042
rect 24584 25978 24636 25984
rect 24596 25498 24624 25978
rect 24688 25906 24716 26182
rect 24780 25974 24808 28999
rect 25148 28762 25176 29038
rect 25596 28960 25648 28966
rect 25596 28902 25648 28908
rect 25261 28860 25569 28869
rect 25261 28858 25267 28860
rect 25323 28858 25347 28860
rect 25403 28858 25427 28860
rect 25483 28858 25507 28860
rect 25563 28858 25569 28860
rect 25323 28806 25325 28858
rect 25505 28806 25507 28858
rect 25261 28804 25267 28806
rect 25323 28804 25347 28806
rect 25403 28804 25427 28806
rect 25483 28804 25507 28806
rect 25563 28804 25569 28806
rect 25261 28795 25569 28804
rect 25136 28756 25188 28762
rect 25136 28698 25188 28704
rect 25608 28558 25636 28902
rect 24952 28552 25004 28558
rect 24952 28494 25004 28500
rect 25596 28552 25648 28558
rect 25596 28494 25648 28500
rect 24860 27872 24912 27878
rect 24860 27814 24912 27820
rect 24872 27470 24900 27814
rect 24964 27674 24992 28494
rect 25044 28484 25096 28490
rect 25044 28426 25096 28432
rect 25056 28150 25084 28426
rect 25688 28416 25740 28422
rect 25688 28358 25740 28364
rect 25044 28144 25096 28150
rect 25044 28086 25096 28092
rect 24952 27668 25004 27674
rect 24952 27610 25004 27616
rect 24860 27464 24912 27470
rect 24860 27406 24912 27412
rect 24768 25968 24820 25974
rect 24768 25910 24820 25916
rect 24676 25900 24728 25906
rect 24676 25842 24728 25848
rect 24688 25786 24716 25842
rect 25056 25838 25084 28086
rect 25700 28082 25728 28358
rect 25136 28076 25188 28082
rect 25136 28018 25188 28024
rect 25688 28076 25740 28082
rect 25688 28018 25740 28024
rect 25044 25832 25096 25838
rect 24688 25758 24808 25786
rect 25044 25774 25096 25780
rect 24676 25696 24728 25702
rect 24676 25638 24728 25644
rect 24584 25492 24636 25498
rect 24584 25434 24636 25440
rect 24492 25288 24544 25294
rect 24492 25230 24544 25236
rect 24400 24812 24452 24818
rect 24400 24754 24452 24760
rect 24412 24410 24440 24754
rect 24596 24682 24624 25434
rect 24688 25242 24716 25638
rect 24780 25362 24808 25758
rect 24768 25356 24820 25362
rect 24768 25298 24820 25304
rect 24952 25356 25004 25362
rect 24952 25298 25004 25304
rect 24860 25288 24912 25294
rect 24688 25236 24860 25242
rect 24688 25230 24912 25236
rect 24688 25214 24900 25230
rect 24584 24676 24636 24682
rect 24584 24618 24636 24624
rect 24688 24614 24716 25214
rect 24676 24608 24728 24614
rect 24676 24550 24728 24556
rect 24400 24404 24452 24410
rect 24400 24346 24452 24352
rect 24216 24064 24268 24070
rect 24216 24006 24268 24012
rect 24228 23798 24256 24006
rect 24216 23792 24268 23798
rect 24216 23734 24268 23740
rect 24228 22710 24256 23734
rect 24308 23656 24360 23662
rect 24308 23598 24360 23604
rect 24320 23050 24348 23598
rect 24400 23520 24452 23526
rect 24400 23462 24452 23468
rect 24308 23044 24360 23050
rect 24308 22986 24360 22992
rect 24216 22704 24268 22710
rect 24216 22646 24268 22652
rect 24228 21894 24256 22646
rect 24320 22438 24348 22986
rect 24412 22438 24440 23462
rect 24308 22432 24360 22438
rect 24308 22374 24360 22380
rect 24400 22432 24452 22438
rect 24400 22374 24452 22380
rect 24688 22094 24716 24550
rect 24964 23866 24992 25298
rect 25044 25152 25096 25158
rect 25044 25094 25096 25100
rect 24952 23860 25004 23866
rect 24952 23802 25004 23808
rect 24768 23724 24820 23730
rect 24768 23666 24820 23672
rect 24780 22778 24808 23666
rect 25056 23186 25084 25094
rect 25148 23798 25176 28018
rect 25688 27872 25740 27878
rect 25688 27814 25740 27820
rect 25261 27772 25569 27781
rect 25261 27770 25267 27772
rect 25323 27770 25347 27772
rect 25403 27770 25427 27772
rect 25483 27770 25507 27772
rect 25563 27770 25569 27772
rect 25323 27718 25325 27770
rect 25505 27718 25507 27770
rect 25261 27716 25267 27718
rect 25323 27716 25347 27718
rect 25403 27716 25427 27718
rect 25483 27716 25507 27718
rect 25563 27716 25569 27718
rect 25261 27707 25569 27716
rect 25700 27402 25728 27814
rect 25688 27396 25740 27402
rect 25688 27338 25740 27344
rect 25596 27328 25648 27334
rect 25596 27270 25648 27276
rect 25261 26684 25569 26693
rect 25261 26682 25267 26684
rect 25323 26682 25347 26684
rect 25403 26682 25427 26684
rect 25483 26682 25507 26684
rect 25563 26682 25569 26684
rect 25323 26630 25325 26682
rect 25505 26630 25507 26682
rect 25261 26628 25267 26630
rect 25323 26628 25347 26630
rect 25403 26628 25427 26630
rect 25483 26628 25507 26630
rect 25563 26628 25569 26630
rect 25261 26619 25569 26628
rect 25608 25702 25636 27270
rect 25792 26058 25820 30602
rect 25872 29504 25924 29510
rect 25872 29446 25924 29452
rect 25884 29170 25912 29446
rect 25872 29164 25924 29170
rect 25872 29106 25924 29112
rect 25884 27690 25912 29106
rect 25976 28626 26004 31078
rect 26068 30938 26096 31282
rect 26056 30932 26108 30938
rect 26056 30874 26108 30880
rect 26056 29844 26108 29850
rect 26056 29786 26108 29792
rect 26068 29170 26096 29786
rect 26148 29572 26200 29578
rect 26148 29514 26200 29520
rect 26160 29238 26188 29514
rect 26148 29232 26200 29238
rect 26148 29174 26200 29180
rect 26056 29164 26108 29170
rect 26056 29106 26108 29112
rect 26160 28642 26188 29174
rect 26240 28960 26292 28966
rect 26240 28902 26292 28908
rect 25964 28620 26016 28626
rect 25964 28562 26016 28568
rect 26068 28614 26188 28642
rect 26068 28422 26096 28614
rect 26148 28484 26200 28490
rect 26148 28426 26200 28432
rect 26056 28416 26108 28422
rect 26056 28358 26108 28364
rect 26068 28082 26096 28358
rect 26160 28218 26188 28426
rect 26148 28212 26200 28218
rect 26148 28154 26200 28160
rect 26252 28098 26280 28902
rect 26056 28076 26108 28082
rect 26056 28018 26108 28024
rect 26160 28070 26280 28098
rect 25884 27662 26004 27690
rect 25872 27464 25924 27470
rect 25872 27406 25924 27412
rect 25884 27130 25912 27406
rect 25872 27124 25924 27130
rect 25872 27066 25924 27072
rect 25700 26030 25820 26058
rect 25596 25696 25648 25702
rect 25596 25638 25648 25644
rect 25261 25596 25569 25605
rect 25261 25594 25267 25596
rect 25323 25594 25347 25596
rect 25403 25594 25427 25596
rect 25483 25594 25507 25596
rect 25563 25594 25569 25596
rect 25323 25542 25325 25594
rect 25505 25542 25507 25594
rect 25261 25540 25267 25542
rect 25323 25540 25347 25542
rect 25403 25540 25427 25542
rect 25483 25540 25507 25542
rect 25563 25540 25569 25542
rect 25261 25531 25569 25540
rect 25228 25220 25280 25226
rect 25228 25162 25280 25168
rect 25240 24818 25268 25162
rect 25228 24812 25280 24818
rect 25228 24754 25280 24760
rect 25504 24812 25556 24818
rect 25700 24800 25728 26030
rect 25780 25900 25832 25906
rect 25780 25842 25832 25848
rect 25792 25498 25820 25842
rect 25780 25492 25832 25498
rect 25780 25434 25832 25440
rect 25792 25242 25820 25434
rect 25976 25362 26004 27662
rect 26068 26926 26096 28018
rect 26160 27946 26188 28070
rect 26148 27940 26200 27946
rect 26148 27882 26200 27888
rect 26160 26994 26188 27882
rect 26148 26988 26200 26994
rect 26148 26930 26200 26936
rect 26056 26920 26108 26926
rect 26056 26862 26108 26868
rect 26148 25832 26200 25838
rect 26148 25774 26200 25780
rect 26056 25696 26108 25702
rect 26056 25638 26108 25644
rect 25964 25356 26016 25362
rect 25964 25298 26016 25304
rect 25792 25214 25912 25242
rect 25884 24818 25912 25214
rect 25556 24772 25728 24800
rect 25504 24754 25556 24760
rect 25700 24614 25728 24772
rect 25780 24812 25832 24818
rect 25780 24754 25832 24760
rect 25872 24812 25924 24818
rect 25872 24754 25924 24760
rect 25688 24608 25740 24614
rect 25688 24550 25740 24556
rect 25261 24508 25569 24517
rect 25261 24506 25267 24508
rect 25323 24506 25347 24508
rect 25403 24506 25427 24508
rect 25483 24506 25507 24508
rect 25563 24506 25569 24508
rect 25323 24454 25325 24506
rect 25505 24454 25507 24506
rect 25261 24452 25267 24454
rect 25323 24452 25347 24454
rect 25403 24452 25427 24454
rect 25483 24452 25507 24454
rect 25563 24452 25569 24454
rect 25261 24443 25569 24452
rect 25792 23866 25820 24754
rect 25780 23860 25832 23866
rect 25780 23802 25832 23808
rect 25136 23792 25188 23798
rect 25136 23734 25188 23740
rect 25044 23180 25096 23186
rect 25044 23122 25096 23128
rect 25148 23118 25176 23734
rect 25261 23420 25569 23429
rect 25261 23418 25267 23420
rect 25323 23418 25347 23420
rect 25403 23418 25427 23420
rect 25483 23418 25507 23420
rect 25563 23418 25569 23420
rect 25323 23366 25325 23418
rect 25505 23366 25507 23418
rect 25261 23364 25267 23366
rect 25323 23364 25347 23366
rect 25403 23364 25427 23366
rect 25483 23364 25507 23366
rect 25563 23364 25569 23366
rect 25261 23355 25569 23364
rect 25228 23248 25280 23254
rect 25228 23190 25280 23196
rect 25136 23112 25188 23118
rect 24964 23060 25136 23066
rect 24964 23054 25188 23060
rect 24964 23038 25176 23054
rect 24768 22772 24820 22778
rect 24820 22732 24900 22760
rect 24768 22714 24820 22720
rect 24872 22098 24900 22732
rect 24688 22066 24808 22094
rect 24584 22024 24636 22030
rect 24584 21966 24636 21972
rect 24492 21956 24544 21962
rect 24492 21898 24544 21904
rect 24216 21888 24268 21894
rect 24216 21830 24268 21836
rect 24504 19922 24532 21898
rect 24596 20398 24624 21966
rect 24780 21894 24808 22066
rect 24860 22092 24912 22098
rect 24860 22034 24912 22040
rect 24768 21888 24820 21894
rect 24768 21830 24820 21836
rect 24676 20596 24728 20602
rect 24676 20538 24728 20544
rect 24584 20392 24636 20398
rect 24584 20334 24636 20340
rect 24492 19916 24544 19922
rect 24492 19858 24544 19864
rect 24688 19786 24716 20538
rect 24780 19922 24808 21830
rect 24964 21418 24992 23038
rect 25240 22930 25268 23190
rect 25148 22902 25268 22930
rect 25872 22976 25924 22982
rect 25872 22918 25924 22924
rect 25044 22568 25096 22574
rect 25044 22510 25096 22516
rect 24952 21412 25004 21418
rect 24952 21354 25004 21360
rect 24964 20942 24992 21354
rect 24952 20936 25004 20942
rect 24952 20878 25004 20884
rect 24964 20534 24992 20878
rect 24952 20528 25004 20534
rect 24952 20470 25004 20476
rect 24768 19916 24820 19922
rect 24768 19858 24820 19864
rect 24860 19848 24912 19854
rect 24860 19790 24912 19796
rect 24676 19780 24728 19786
rect 24676 19722 24728 19728
rect 24216 18896 24268 18902
rect 24216 18838 24268 18844
rect 24228 18290 24256 18838
rect 24688 18834 24716 19722
rect 24872 18970 24900 19790
rect 24860 18964 24912 18970
rect 24860 18906 24912 18912
rect 24676 18828 24728 18834
rect 24676 18770 24728 18776
rect 24688 18426 24716 18770
rect 24860 18760 24912 18766
rect 24860 18702 24912 18708
rect 24676 18420 24728 18426
rect 24676 18362 24728 18368
rect 24216 18284 24268 18290
rect 24216 18226 24268 18232
rect 24584 18216 24636 18222
rect 24584 18158 24636 18164
rect 24400 18080 24452 18086
rect 24400 18022 24452 18028
rect 24124 17332 24176 17338
rect 24124 17274 24176 17280
rect 24412 17202 24440 18022
rect 24596 17542 24624 18158
rect 24584 17536 24636 17542
rect 24584 17478 24636 17484
rect 24400 17196 24452 17202
rect 24400 17138 24452 17144
rect 24596 16522 24624 17478
rect 24584 16516 24636 16522
rect 24584 16458 24636 16464
rect 24872 16182 24900 18702
rect 24964 16726 24992 20470
rect 25056 19922 25084 22510
rect 25148 22094 25176 22902
rect 25884 22710 25912 22918
rect 25872 22704 25924 22710
rect 25872 22646 25924 22652
rect 25261 22332 25569 22341
rect 25261 22330 25267 22332
rect 25323 22330 25347 22332
rect 25403 22330 25427 22332
rect 25483 22330 25507 22332
rect 25563 22330 25569 22332
rect 25323 22278 25325 22330
rect 25505 22278 25507 22330
rect 25261 22276 25267 22278
rect 25323 22276 25347 22278
rect 25403 22276 25427 22278
rect 25483 22276 25507 22278
rect 25563 22276 25569 22278
rect 25261 22267 25569 22276
rect 25964 22094 26016 22098
rect 26068 22094 26096 25638
rect 26160 23254 26188 25774
rect 26240 24676 26292 24682
rect 26240 24618 26292 24624
rect 26252 23866 26280 24618
rect 26240 23860 26292 23866
rect 26240 23802 26292 23808
rect 26148 23248 26200 23254
rect 26148 23190 26200 23196
rect 25148 22066 25268 22094
rect 25136 21888 25188 21894
rect 25136 21830 25188 21836
rect 25148 21554 25176 21830
rect 25240 21554 25268 22066
rect 25964 22092 26096 22094
rect 26016 22066 26096 22092
rect 25964 22034 26016 22040
rect 25136 21548 25188 21554
rect 25136 21490 25188 21496
rect 25228 21548 25280 21554
rect 25228 21490 25280 21496
rect 25688 21548 25740 21554
rect 25688 21490 25740 21496
rect 25596 21344 25648 21350
rect 25596 21286 25648 21292
rect 25261 21244 25569 21253
rect 25261 21242 25267 21244
rect 25323 21242 25347 21244
rect 25403 21242 25427 21244
rect 25483 21242 25507 21244
rect 25563 21242 25569 21244
rect 25323 21190 25325 21242
rect 25505 21190 25507 21242
rect 25261 21188 25267 21190
rect 25323 21188 25347 21190
rect 25403 21188 25427 21190
rect 25483 21188 25507 21190
rect 25563 21188 25569 21190
rect 25261 21179 25569 21188
rect 25608 20942 25636 21286
rect 25700 20942 25728 21490
rect 26146 21448 26202 21457
rect 26146 21383 26202 21392
rect 25596 20936 25648 20942
rect 25596 20878 25648 20884
rect 25688 20936 25740 20942
rect 25688 20878 25740 20884
rect 25964 20936 26016 20942
rect 25964 20878 26016 20884
rect 25700 20534 25728 20878
rect 25688 20528 25740 20534
rect 25688 20470 25740 20476
rect 25136 20460 25188 20466
rect 25136 20402 25188 20408
rect 25148 20058 25176 20402
rect 25700 20346 25728 20470
rect 25976 20398 26004 20878
rect 26056 20800 26108 20806
rect 26056 20742 26108 20748
rect 25608 20318 25728 20346
rect 25964 20392 26016 20398
rect 25964 20334 26016 20340
rect 25261 20156 25569 20165
rect 25261 20154 25267 20156
rect 25323 20154 25347 20156
rect 25403 20154 25427 20156
rect 25483 20154 25507 20156
rect 25563 20154 25569 20156
rect 25323 20102 25325 20154
rect 25505 20102 25507 20154
rect 25261 20100 25267 20102
rect 25323 20100 25347 20102
rect 25403 20100 25427 20102
rect 25483 20100 25507 20102
rect 25563 20100 25569 20102
rect 25261 20091 25569 20100
rect 25136 20052 25188 20058
rect 25136 19994 25188 20000
rect 25044 19916 25096 19922
rect 25044 19858 25096 19864
rect 25056 18290 25084 19858
rect 25608 19854 25636 20318
rect 25688 20256 25740 20262
rect 25688 20198 25740 20204
rect 25596 19848 25648 19854
rect 25596 19790 25648 19796
rect 25261 19068 25569 19077
rect 25261 19066 25267 19068
rect 25323 19066 25347 19068
rect 25403 19066 25427 19068
rect 25483 19066 25507 19068
rect 25563 19066 25569 19068
rect 25323 19014 25325 19066
rect 25505 19014 25507 19066
rect 25261 19012 25267 19014
rect 25323 19012 25347 19014
rect 25403 19012 25427 19014
rect 25483 19012 25507 19014
rect 25563 19012 25569 19014
rect 25261 19003 25569 19012
rect 25700 18358 25728 20198
rect 25976 20058 26004 20334
rect 25964 20052 26016 20058
rect 25964 19994 26016 20000
rect 26068 19854 26096 20742
rect 26056 19848 26108 19854
rect 26056 19790 26108 19796
rect 26160 18834 26188 21383
rect 26344 20330 26372 31758
rect 26436 30122 26464 32438
rect 26528 32434 26556 32846
rect 26516 32428 26568 32434
rect 26516 32370 26568 32376
rect 26700 32224 26752 32230
rect 26700 32166 26752 32172
rect 26712 31890 26740 32166
rect 26700 31884 26752 31890
rect 26700 31826 26752 31832
rect 26516 31680 26568 31686
rect 26516 31622 26568 31628
rect 26528 31346 26556 31622
rect 26516 31340 26568 31346
rect 26516 31282 26568 31288
rect 26424 30116 26476 30122
rect 26424 30058 26476 30064
rect 26528 28150 26556 31282
rect 26700 31136 26752 31142
rect 26700 31078 26752 31084
rect 26712 30734 26740 31078
rect 26700 30728 26752 30734
rect 26700 30670 26752 30676
rect 26608 30252 26660 30258
rect 26608 30194 26660 30200
rect 26620 30025 26648 30194
rect 26606 30016 26662 30025
rect 26606 29951 26662 29960
rect 26516 28144 26568 28150
rect 26516 28086 26568 28092
rect 26608 28008 26660 28014
rect 26608 27950 26660 27956
rect 26620 26858 26648 27950
rect 26608 26852 26660 26858
rect 26608 26794 26660 26800
rect 26516 26784 26568 26790
rect 26516 26726 26568 26732
rect 26528 26450 26556 26726
rect 26516 26444 26568 26450
rect 26516 26386 26568 26392
rect 26620 25906 26648 26794
rect 26700 26308 26752 26314
rect 26700 26250 26752 26256
rect 26712 26042 26740 26250
rect 26700 26036 26752 26042
rect 26700 25978 26752 25984
rect 26608 25900 26660 25906
rect 26608 25842 26660 25848
rect 26424 24744 26476 24750
rect 26424 24686 26476 24692
rect 26436 24410 26464 24686
rect 26620 24682 26648 25842
rect 26700 24744 26752 24750
rect 26700 24686 26752 24692
rect 26608 24676 26660 24682
rect 26608 24618 26660 24624
rect 26516 24608 26568 24614
rect 26516 24550 26568 24556
rect 26424 24404 26476 24410
rect 26424 24346 26476 24352
rect 26436 23730 26464 24346
rect 26528 23730 26556 24550
rect 26424 23724 26476 23730
rect 26424 23666 26476 23672
rect 26516 23724 26568 23730
rect 26516 23666 26568 23672
rect 26436 22778 26464 23666
rect 26712 23662 26740 24686
rect 26804 23730 26832 35866
rect 26896 33522 26924 38218
rect 26884 33516 26936 33522
rect 26884 33458 26936 33464
rect 26884 33380 26936 33386
rect 26884 33322 26936 33328
rect 26896 25906 26924 33322
rect 26988 31754 27016 39918
rect 27080 32434 27108 43250
rect 27264 42226 27292 43726
rect 27434 42256 27490 42265
rect 27252 42220 27304 42226
rect 27632 42226 27660 46582
rect 27724 45626 27752 49200
rect 27804 47048 27856 47054
rect 27804 46990 27856 46996
rect 27712 45620 27764 45626
rect 27712 45562 27764 45568
rect 27816 45014 27844 46990
rect 28368 46510 28396 49200
rect 28630 47696 28686 47705
rect 28630 47631 28686 47640
rect 28356 46504 28408 46510
rect 28356 46446 28408 46452
rect 27896 45484 27948 45490
rect 27896 45426 27948 45432
rect 27908 45082 27936 45426
rect 27896 45076 27948 45082
rect 27896 45018 27948 45024
rect 27804 45008 27856 45014
rect 27804 44950 27856 44956
rect 27804 44736 27856 44742
rect 27804 44678 27856 44684
rect 27816 44402 27844 44678
rect 27804 44396 27856 44402
rect 27804 44338 27856 44344
rect 27908 43314 27936 45018
rect 28354 44976 28410 44985
rect 28354 44911 28356 44920
rect 28408 44911 28410 44920
rect 28356 44882 28408 44888
rect 27896 43308 27948 43314
rect 27896 43250 27948 43256
rect 28080 43104 28132 43110
rect 28080 43046 28132 43052
rect 28092 42770 28120 43046
rect 28080 42764 28132 42770
rect 28080 42706 28132 42712
rect 27804 42628 27856 42634
rect 27804 42570 27856 42576
rect 27816 42362 27844 42570
rect 27804 42356 27856 42362
rect 27804 42298 27856 42304
rect 27434 42191 27490 42200
rect 27620 42220 27672 42226
rect 27252 42162 27304 42168
rect 27344 41540 27396 41546
rect 27344 41482 27396 41488
rect 27356 40050 27384 41482
rect 27344 40044 27396 40050
rect 27344 39986 27396 39992
rect 27344 38956 27396 38962
rect 27344 38898 27396 38904
rect 27356 37874 27384 38898
rect 27344 37868 27396 37874
rect 27344 37810 27396 37816
rect 27342 36816 27398 36825
rect 27342 36751 27344 36760
rect 27396 36751 27398 36760
rect 27344 36722 27396 36728
rect 27448 36242 27476 42191
rect 27620 42162 27672 42168
rect 27528 41676 27580 41682
rect 27528 41618 27580 41624
rect 27540 40905 27568 41618
rect 27632 41414 27660 42162
rect 27896 41472 27948 41478
rect 27896 41414 27948 41420
rect 27632 41386 27752 41414
rect 27526 40896 27582 40905
rect 27526 40831 27582 40840
rect 27724 37806 27752 41386
rect 27908 41138 27936 41414
rect 27896 41132 27948 41138
rect 27896 41074 27948 41080
rect 28644 40594 28672 47631
rect 28734 46812 29042 46821
rect 28734 46810 28740 46812
rect 28796 46810 28820 46812
rect 28876 46810 28900 46812
rect 28956 46810 28980 46812
rect 29036 46810 29042 46812
rect 28796 46758 28798 46810
rect 28978 46758 28980 46810
rect 28734 46756 28740 46758
rect 28796 46756 28820 46758
rect 28876 46756 28900 46758
rect 28956 46756 28980 46758
rect 29036 46756 29042 46758
rect 28734 46747 29042 46756
rect 28734 45724 29042 45733
rect 28734 45722 28740 45724
rect 28796 45722 28820 45724
rect 28876 45722 28900 45724
rect 28956 45722 28980 45724
rect 29036 45722 29042 45724
rect 28796 45670 28798 45722
rect 28978 45670 28980 45722
rect 28734 45668 28740 45670
rect 28796 45668 28820 45670
rect 28876 45668 28900 45670
rect 28956 45668 28980 45670
rect 29036 45668 29042 45670
rect 28734 45659 29042 45668
rect 28734 44636 29042 44645
rect 28734 44634 28740 44636
rect 28796 44634 28820 44636
rect 28876 44634 28900 44636
rect 28956 44634 28980 44636
rect 29036 44634 29042 44636
rect 28796 44582 28798 44634
rect 28978 44582 28980 44634
rect 28734 44580 28740 44582
rect 28796 44580 28820 44582
rect 28876 44580 28900 44582
rect 28956 44580 28980 44582
rect 29036 44580 29042 44582
rect 28734 44571 29042 44580
rect 28734 43548 29042 43557
rect 28734 43546 28740 43548
rect 28796 43546 28820 43548
rect 28876 43546 28900 43548
rect 28956 43546 28980 43548
rect 29036 43546 29042 43548
rect 28796 43494 28798 43546
rect 28978 43494 28980 43546
rect 28734 43492 28740 43494
rect 28796 43492 28820 43494
rect 28876 43492 28900 43494
rect 28956 43492 28980 43494
rect 29036 43492 29042 43494
rect 28734 43483 29042 43492
rect 28734 42460 29042 42469
rect 28734 42458 28740 42460
rect 28796 42458 28820 42460
rect 28876 42458 28900 42460
rect 28956 42458 28980 42460
rect 29036 42458 29042 42460
rect 28796 42406 28798 42458
rect 28978 42406 28980 42458
rect 28734 42404 28740 42406
rect 28796 42404 28820 42406
rect 28876 42404 28900 42406
rect 28956 42404 28980 42406
rect 29036 42404 29042 42406
rect 28734 42395 29042 42404
rect 28734 41372 29042 41381
rect 28734 41370 28740 41372
rect 28796 41370 28820 41372
rect 28876 41370 28900 41372
rect 28956 41370 28980 41372
rect 29036 41370 29042 41372
rect 28796 41318 28798 41370
rect 28978 41318 28980 41370
rect 28734 41316 28740 41318
rect 28796 41316 28820 41318
rect 28876 41316 28900 41318
rect 28956 41316 28980 41318
rect 29036 41316 29042 41318
rect 28734 41307 29042 41316
rect 28632 40588 28684 40594
rect 28632 40530 28684 40536
rect 28734 40284 29042 40293
rect 28734 40282 28740 40284
rect 28796 40282 28820 40284
rect 28876 40282 28900 40284
rect 28956 40282 28980 40284
rect 29036 40282 29042 40284
rect 28796 40230 28798 40282
rect 28978 40230 28980 40282
rect 28734 40228 28740 40230
rect 28796 40228 28820 40230
rect 28876 40228 28900 40230
rect 28956 40228 28980 40230
rect 29036 40228 29042 40230
rect 28734 40219 29042 40228
rect 29918 40216 29974 40225
rect 29918 40151 29974 40160
rect 27896 39840 27948 39846
rect 27896 39782 27948 39788
rect 27908 39506 27936 39782
rect 28630 39536 28686 39545
rect 27896 39500 27948 39506
rect 29932 39506 29960 40151
rect 28630 39471 28686 39480
rect 29920 39500 29972 39506
rect 27896 39442 27948 39448
rect 28644 38418 28672 39471
rect 29920 39442 29972 39448
rect 28734 39196 29042 39205
rect 28734 39194 28740 39196
rect 28796 39194 28820 39196
rect 28876 39194 28900 39196
rect 28956 39194 28980 39196
rect 29036 39194 29042 39196
rect 28796 39142 28798 39194
rect 28978 39142 28980 39194
rect 28734 39140 28740 39142
rect 28796 39140 28820 39142
rect 28876 39140 28900 39142
rect 28956 39140 28980 39142
rect 29036 39140 29042 39142
rect 28734 39131 29042 39140
rect 28632 38412 28684 38418
rect 28632 38354 28684 38360
rect 28734 38108 29042 38117
rect 28734 38106 28740 38108
rect 28796 38106 28820 38108
rect 28876 38106 28900 38108
rect 28956 38106 28980 38108
rect 29036 38106 29042 38108
rect 28796 38054 28798 38106
rect 28978 38054 28980 38106
rect 28734 38052 28740 38054
rect 28796 38052 28820 38054
rect 28876 38052 28900 38054
rect 28956 38052 28980 38054
rect 29036 38052 29042 38054
rect 28734 38043 29042 38052
rect 27988 37868 28040 37874
rect 27988 37810 28040 37816
rect 27712 37800 27764 37806
rect 27712 37742 27764 37748
rect 27436 36236 27488 36242
rect 27436 36178 27488 36184
rect 27724 35894 27752 37742
rect 27896 37188 27948 37194
rect 27896 37130 27948 37136
rect 27908 36922 27936 37130
rect 27896 36916 27948 36922
rect 27896 36858 27948 36864
rect 27804 36780 27856 36786
rect 27804 36722 27856 36728
rect 27632 35866 27752 35894
rect 27528 35148 27580 35154
rect 27528 35090 27580 35096
rect 27160 34400 27212 34406
rect 27160 34342 27212 34348
rect 27172 33454 27200 34342
rect 27540 34105 27568 35090
rect 27526 34096 27582 34105
rect 27526 34031 27582 34040
rect 27252 33924 27304 33930
rect 27252 33866 27304 33872
rect 27264 33658 27292 33866
rect 27252 33652 27304 33658
rect 27252 33594 27304 33600
rect 27160 33448 27212 33454
rect 27160 33390 27212 33396
rect 27528 32972 27580 32978
rect 27528 32914 27580 32920
rect 27068 32428 27120 32434
rect 27068 32370 27120 32376
rect 27434 32328 27490 32337
rect 27434 32263 27490 32272
rect 26988 31726 27292 31754
rect 26884 25900 26936 25906
rect 26884 25842 26936 25848
rect 26792 23724 26844 23730
rect 26792 23666 26844 23672
rect 27068 23724 27120 23730
rect 27068 23666 27120 23672
rect 26700 23656 26752 23662
rect 26700 23598 26752 23604
rect 26700 23520 26752 23526
rect 26700 23462 26752 23468
rect 26712 23186 26740 23462
rect 26700 23180 26752 23186
rect 26700 23122 26752 23128
rect 26424 22772 26476 22778
rect 26424 22714 26476 22720
rect 26332 20324 26384 20330
rect 26332 20266 26384 20272
rect 26148 18828 26200 18834
rect 26148 18770 26200 18776
rect 26700 18624 26752 18630
rect 26700 18566 26752 18572
rect 25688 18352 25740 18358
rect 25688 18294 25740 18300
rect 25044 18284 25096 18290
rect 25044 18226 25096 18232
rect 25056 17270 25084 18226
rect 25261 17980 25569 17989
rect 25261 17978 25267 17980
rect 25323 17978 25347 17980
rect 25403 17978 25427 17980
rect 25483 17978 25507 17980
rect 25563 17978 25569 17980
rect 25323 17926 25325 17978
rect 25505 17926 25507 17978
rect 25261 17924 25267 17926
rect 25323 17924 25347 17926
rect 25403 17924 25427 17926
rect 25483 17924 25507 17926
rect 25563 17924 25569 17926
rect 25261 17915 25569 17924
rect 26712 17746 26740 18566
rect 26700 17740 26752 17746
rect 26700 17682 26752 17688
rect 25504 17536 25556 17542
rect 25504 17478 25556 17484
rect 25516 17338 25544 17478
rect 25504 17332 25556 17338
rect 25504 17274 25556 17280
rect 25044 17264 25096 17270
rect 25044 17206 25096 17212
rect 24952 16720 25004 16726
rect 24952 16662 25004 16668
rect 24860 16176 24912 16182
rect 24860 16118 24912 16124
rect 25056 15570 25084 17206
rect 26240 17196 26292 17202
rect 26240 17138 26292 17144
rect 25872 16992 25924 16998
rect 25872 16934 25924 16940
rect 25261 16892 25569 16901
rect 25261 16890 25267 16892
rect 25323 16890 25347 16892
rect 25403 16890 25427 16892
rect 25483 16890 25507 16892
rect 25563 16890 25569 16892
rect 25323 16838 25325 16890
rect 25505 16838 25507 16890
rect 25261 16836 25267 16838
rect 25323 16836 25347 16838
rect 25403 16836 25427 16838
rect 25483 16836 25507 16838
rect 25563 16836 25569 16838
rect 25261 16827 25569 16836
rect 25884 16522 25912 16934
rect 26252 16522 26280 17138
rect 26700 16992 26752 16998
rect 26700 16934 26752 16940
rect 26712 16658 26740 16934
rect 26700 16652 26752 16658
rect 26700 16594 26752 16600
rect 25872 16516 25924 16522
rect 25872 16458 25924 16464
rect 26240 16516 26292 16522
rect 26240 16458 26292 16464
rect 25884 16402 25912 16458
rect 25884 16374 26004 16402
rect 25976 16046 26004 16374
rect 26252 16250 26280 16458
rect 26240 16244 26292 16250
rect 26240 16186 26292 16192
rect 26240 16108 26292 16114
rect 26240 16050 26292 16056
rect 25964 16040 26016 16046
rect 25964 15982 26016 15988
rect 25261 15804 25569 15813
rect 25261 15802 25267 15804
rect 25323 15802 25347 15804
rect 25403 15802 25427 15804
rect 25483 15802 25507 15804
rect 25563 15802 25569 15804
rect 25323 15750 25325 15802
rect 25505 15750 25507 15802
rect 25261 15748 25267 15750
rect 25323 15748 25347 15750
rect 25403 15748 25427 15750
rect 25483 15748 25507 15750
rect 25563 15748 25569 15750
rect 25261 15739 25569 15748
rect 25044 15564 25096 15570
rect 25044 15506 25096 15512
rect 25056 15026 25084 15506
rect 25504 15496 25556 15502
rect 25504 15438 25556 15444
rect 25516 15065 25544 15438
rect 25502 15056 25558 15065
rect 25044 15020 25096 15026
rect 25044 14962 25096 14968
rect 25136 15020 25188 15026
rect 25502 14991 25558 15000
rect 25136 14962 25188 14968
rect 24216 14816 24268 14822
rect 24216 14758 24268 14764
rect 24032 14068 24084 14074
rect 24032 14010 24084 14016
rect 24044 13326 24072 14010
rect 24228 13938 24256 14758
rect 24308 14272 24360 14278
rect 24308 14214 24360 14220
rect 24216 13932 24268 13938
rect 24216 13874 24268 13880
rect 24320 13802 24348 14214
rect 25148 14074 25176 14962
rect 25261 14716 25569 14725
rect 25261 14714 25267 14716
rect 25323 14714 25347 14716
rect 25403 14714 25427 14716
rect 25483 14714 25507 14716
rect 25563 14714 25569 14716
rect 25323 14662 25325 14714
rect 25505 14662 25507 14714
rect 25261 14660 25267 14662
rect 25323 14660 25347 14662
rect 25403 14660 25427 14662
rect 25483 14660 25507 14662
rect 25563 14660 25569 14662
rect 25261 14651 25569 14660
rect 25780 14340 25832 14346
rect 25780 14282 25832 14288
rect 25792 14074 25820 14282
rect 25136 14068 25188 14074
rect 25136 14010 25188 14016
rect 25780 14068 25832 14074
rect 25780 14010 25832 14016
rect 24584 13932 24636 13938
rect 24584 13874 24636 13880
rect 25596 13932 25648 13938
rect 25596 13874 25648 13880
rect 24308 13796 24360 13802
rect 24308 13738 24360 13744
rect 24596 13530 24624 13874
rect 24676 13728 24728 13734
rect 24676 13670 24728 13676
rect 24688 13530 24716 13670
rect 25261 13628 25569 13637
rect 25261 13626 25267 13628
rect 25323 13626 25347 13628
rect 25403 13626 25427 13628
rect 25483 13626 25507 13628
rect 25563 13626 25569 13628
rect 25323 13574 25325 13626
rect 25505 13574 25507 13626
rect 25261 13572 25267 13574
rect 25323 13572 25347 13574
rect 25403 13572 25427 13574
rect 25483 13572 25507 13574
rect 25563 13572 25569 13574
rect 25261 13563 25569 13572
rect 25608 13530 25636 13874
rect 24584 13524 24636 13530
rect 24584 13466 24636 13472
rect 24676 13524 24728 13530
rect 24676 13466 24728 13472
rect 25596 13524 25648 13530
rect 25596 13466 25648 13472
rect 25976 13326 26004 15982
rect 26056 15564 26108 15570
rect 26056 15506 26108 15512
rect 26068 15094 26096 15506
rect 26252 15162 26280 16050
rect 26240 15156 26292 15162
rect 26240 15098 26292 15104
rect 26056 15088 26108 15094
rect 26056 15030 26108 15036
rect 26068 14482 26096 15030
rect 26056 14476 26108 14482
rect 26056 14418 26108 14424
rect 26240 14272 26292 14278
rect 26240 14214 26292 14220
rect 24032 13320 24084 13326
rect 24032 13262 24084 13268
rect 25872 13320 25924 13326
rect 25872 13262 25924 13268
rect 25964 13320 26016 13326
rect 25964 13262 26016 13268
rect 24952 13252 25004 13258
rect 24952 13194 25004 13200
rect 23940 12912 23992 12918
rect 23940 12854 23992 12860
rect 22744 12776 22796 12782
rect 22744 12718 22796 12724
rect 23848 12776 23900 12782
rect 23848 12718 23900 12724
rect 24964 12306 24992 13194
rect 25884 12986 25912 13262
rect 26252 12986 26280 14214
rect 25872 12980 25924 12986
rect 25872 12922 25924 12928
rect 26240 12980 26292 12986
rect 26240 12922 26292 12928
rect 26976 12844 27028 12850
rect 26976 12786 27028 12792
rect 26516 12708 26568 12714
rect 26516 12650 26568 12656
rect 25261 12540 25569 12549
rect 25261 12538 25267 12540
rect 25323 12538 25347 12540
rect 25403 12538 25427 12540
rect 25483 12538 25507 12540
rect 25563 12538 25569 12540
rect 25323 12486 25325 12538
rect 25505 12486 25507 12538
rect 25261 12484 25267 12486
rect 25323 12484 25347 12486
rect 25403 12484 25427 12486
rect 25483 12484 25507 12486
rect 25563 12484 25569 12486
rect 25261 12475 25569 12484
rect 26528 12306 26556 12650
rect 26700 12640 26752 12646
rect 26700 12582 26752 12588
rect 26712 12306 26740 12582
rect 24952 12300 25004 12306
rect 24952 12242 25004 12248
rect 26516 12300 26568 12306
rect 26516 12242 26568 12248
rect 26700 12300 26752 12306
rect 26700 12242 26752 12248
rect 21640 12232 21692 12238
rect 21640 12174 21692 12180
rect 21788 11996 22096 12005
rect 21788 11994 21794 11996
rect 21850 11994 21874 11996
rect 21930 11994 21954 11996
rect 22010 11994 22034 11996
rect 22090 11994 22096 11996
rect 21850 11942 21852 11994
rect 22032 11942 22034 11994
rect 21788 11940 21794 11942
rect 21850 11940 21874 11942
rect 21930 11940 21954 11942
rect 22010 11940 22034 11942
rect 22090 11940 22096 11942
rect 21788 11931 22096 11940
rect 26700 11552 26752 11558
rect 26700 11494 26752 11500
rect 25261 11452 25569 11461
rect 25261 11450 25267 11452
rect 25323 11450 25347 11452
rect 25403 11450 25427 11452
rect 25483 11450 25507 11452
rect 25563 11450 25569 11452
rect 25323 11398 25325 11450
rect 25505 11398 25507 11450
rect 25261 11396 25267 11398
rect 25323 11396 25347 11398
rect 25403 11396 25427 11398
rect 25483 11396 25507 11398
rect 25563 11396 25569 11398
rect 25261 11387 25569 11396
rect 26712 11218 26740 11494
rect 26700 11212 26752 11218
rect 26700 11154 26752 11160
rect 26516 11144 26568 11150
rect 26516 11086 26568 11092
rect 21788 10908 22096 10917
rect 21788 10906 21794 10908
rect 21850 10906 21874 10908
rect 21930 10906 21954 10908
rect 22010 10906 22034 10908
rect 22090 10906 22096 10908
rect 21850 10854 21852 10906
rect 22032 10854 22034 10906
rect 21788 10852 21794 10854
rect 21850 10852 21874 10854
rect 21930 10852 21954 10854
rect 22010 10852 22034 10854
rect 22090 10852 22096 10854
rect 21788 10843 22096 10852
rect 26528 10674 26556 11086
rect 26516 10668 26568 10674
rect 26516 10610 26568 10616
rect 25261 10364 25569 10373
rect 25261 10362 25267 10364
rect 25323 10362 25347 10364
rect 25403 10362 25427 10364
rect 25483 10362 25507 10364
rect 25563 10362 25569 10364
rect 25323 10310 25325 10362
rect 25505 10310 25507 10362
rect 25261 10308 25267 10310
rect 25323 10308 25347 10310
rect 25403 10308 25427 10310
rect 25483 10308 25507 10310
rect 25563 10308 25569 10310
rect 25261 10299 25569 10308
rect 21788 9820 22096 9829
rect 21788 9818 21794 9820
rect 21850 9818 21874 9820
rect 21930 9818 21954 9820
rect 22010 9818 22034 9820
rect 22090 9818 22096 9820
rect 21850 9766 21852 9818
rect 22032 9766 22034 9818
rect 21788 9764 21794 9766
rect 21850 9764 21874 9766
rect 21930 9764 21954 9766
rect 22010 9764 22034 9766
rect 22090 9764 22096 9766
rect 21788 9755 22096 9764
rect 20536 9580 20588 9586
rect 20536 9522 20588 9528
rect 20628 9376 20680 9382
rect 20628 9318 20680 9324
rect 18315 9276 18623 9285
rect 18315 9274 18321 9276
rect 18377 9274 18401 9276
rect 18457 9274 18481 9276
rect 18537 9274 18561 9276
rect 18617 9274 18623 9276
rect 18377 9222 18379 9274
rect 18559 9222 18561 9274
rect 18315 9220 18321 9222
rect 18377 9220 18401 9222
rect 18457 9220 18481 9222
rect 18537 9220 18561 9222
rect 18617 9220 18623 9222
rect 18315 9211 18623 9220
rect 18315 8188 18623 8197
rect 18315 8186 18321 8188
rect 18377 8186 18401 8188
rect 18457 8186 18481 8188
rect 18537 8186 18561 8188
rect 18617 8186 18623 8188
rect 18377 8134 18379 8186
rect 18559 8134 18561 8186
rect 18315 8132 18321 8134
rect 18377 8132 18401 8134
rect 18457 8132 18481 8134
rect 18537 8132 18561 8134
rect 18617 8132 18623 8134
rect 18315 8123 18623 8132
rect 18315 7100 18623 7109
rect 18315 7098 18321 7100
rect 18377 7098 18401 7100
rect 18457 7098 18481 7100
rect 18537 7098 18561 7100
rect 18617 7098 18623 7100
rect 18377 7046 18379 7098
rect 18559 7046 18561 7098
rect 18315 7044 18321 7046
rect 18377 7044 18401 7046
rect 18457 7044 18481 7046
rect 18537 7044 18561 7046
rect 18617 7044 18623 7046
rect 18315 7035 18623 7044
rect 18315 6012 18623 6021
rect 18315 6010 18321 6012
rect 18377 6010 18401 6012
rect 18457 6010 18481 6012
rect 18537 6010 18561 6012
rect 18617 6010 18623 6012
rect 18377 5958 18379 6010
rect 18559 5958 18561 6010
rect 18315 5956 18321 5958
rect 18377 5956 18401 5958
rect 18457 5956 18481 5958
rect 18537 5956 18561 5958
rect 18617 5956 18623 5958
rect 18315 5947 18623 5956
rect 18315 4924 18623 4933
rect 18315 4922 18321 4924
rect 18377 4922 18401 4924
rect 18457 4922 18481 4924
rect 18537 4922 18561 4924
rect 18617 4922 18623 4924
rect 18377 4870 18379 4922
rect 18559 4870 18561 4922
rect 18315 4868 18321 4870
rect 18377 4868 18401 4870
rect 18457 4868 18481 4870
rect 18537 4868 18561 4870
rect 18617 4868 18623 4870
rect 18315 4859 18623 4868
rect 20640 4690 20668 9318
rect 25261 9276 25569 9285
rect 25261 9274 25267 9276
rect 25323 9274 25347 9276
rect 25403 9274 25427 9276
rect 25483 9274 25507 9276
rect 25563 9274 25569 9276
rect 25323 9222 25325 9274
rect 25505 9222 25507 9274
rect 25261 9220 25267 9222
rect 25323 9220 25347 9222
rect 25403 9220 25427 9222
rect 25483 9220 25507 9222
rect 25563 9220 25569 9222
rect 25261 9211 25569 9220
rect 26516 8968 26568 8974
rect 26516 8910 26568 8916
rect 21788 8732 22096 8741
rect 21788 8730 21794 8732
rect 21850 8730 21874 8732
rect 21930 8730 21954 8732
rect 22010 8730 22034 8732
rect 22090 8730 22096 8732
rect 21850 8678 21852 8730
rect 22032 8678 22034 8730
rect 21788 8676 21794 8678
rect 21850 8676 21874 8678
rect 21930 8676 21954 8678
rect 22010 8676 22034 8678
rect 22090 8676 22096 8678
rect 21788 8667 22096 8676
rect 26528 8566 26556 8910
rect 26516 8560 26568 8566
rect 26516 8502 26568 8508
rect 26608 8288 26660 8294
rect 26146 8256 26202 8265
rect 26608 8230 26660 8236
rect 25261 8188 25569 8197
rect 26146 8191 26202 8200
rect 25261 8186 25267 8188
rect 25323 8186 25347 8188
rect 25403 8186 25427 8188
rect 25483 8186 25507 8188
rect 25563 8186 25569 8188
rect 25323 8134 25325 8186
rect 25505 8134 25507 8186
rect 25261 8132 25267 8134
rect 25323 8132 25347 8134
rect 25403 8132 25427 8134
rect 25483 8132 25507 8134
rect 25563 8132 25569 8134
rect 25261 8123 25569 8132
rect 25688 7880 25740 7886
rect 25688 7822 25740 7828
rect 21788 7644 22096 7653
rect 21788 7642 21794 7644
rect 21850 7642 21874 7644
rect 21930 7642 21954 7644
rect 22010 7642 22034 7644
rect 22090 7642 22096 7644
rect 21850 7590 21852 7642
rect 22032 7590 22034 7642
rect 21788 7588 21794 7590
rect 21850 7588 21874 7590
rect 21930 7588 21954 7590
rect 22010 7588 22034 7590
rect 22090 7588 22096 7590
rect 21788 7579 22096 7588
rect 25261 7100 25569 7109
rect 25261 7098 25267 7100
rect 25323 7098 25347 7100
rect 25403 7098 25427 7100
rect 25483 7098 25507 7100
rect 25563 7098 25569 7100
rect 25323 7046 25325 7098
rect 25505 7046 25507 7098
rect 25261 7044 25267 7046
rect 25323 7044 25347 7046
rect 25403 7044 25427 7046
rect 25483 7044 25507 7046
rect 25563 7044 25569 7046
rect 25261 7035 25569 7044
rect 21788 6556 22096 6565
rect 21788 6554 21794 6556
rect 21850 6554 21874 6556
rect 21930 6554 21954 6556
rect 22010 6554 22034 6556
rect 22090 6554 22096 6556
rect 21850 6502 21852 6554
rect 22032 6502 22034 6554
rect 21788 6500 21794 6502
rect 21850 6500 21874 6502
rect 21930 6500 21954 6502
rect 22010 6500 22034 6502
rect 22090 6500 22096 6502
rect 21788 6491 22096 6500
rect 25261 6012 25569 6021
rect 25261 6010 25267 6012
rect 25323 6010 25347 6012
rect 25403 6010 25427 6012
rect 25483 6010 25507 6012
rect 25563 6010 25569 6012
rect 25323 5958 25325 6010
rect 25505 5958 25507 6010
rect 25261 5956 25267 5958
rect 25323 5956 25347 5958
rect 25403 5956 25427 5958
rect 25483 5956 25507 5958
rect 25563 5956 25569 5958
rect 25261 5947 25569 5956
rect 21788 5468 22096 5477
rect 21788 5466 21794 5468
rect 21850 5466 21874 5468
rect 21930 5466 21954 5468
rect 22010 5466 22034 5468
rect 22090 5466 22096 5468
rect 21850 5414 21852 5466
rect 22032 5414 22034 5466
rect 21788 5412 21794 5414
rect 21850 5412 21874 5414
rect 21930 5412 21954 5414
rect 22010 5412 22034 5414
rect 22090 5412 22096 5414
rect 21788 5403 22096 5412
rect 25261 4924 25569 4933
rect 25261 4922 25267 4924
rect 25323 4922 25347 4924
rect 25403 4922 25427 4924
rect 25483 4922 25507 4924
rect 25563 4922 25569 4924
rect 25323 4870 25325 4922
rect 25505 4870 25507 4922
rect 25261 4868 25267 4870
rect 25323 4868 25347 4870
rect 25403 4868 25427 4870
rect 25483 4868 25507 4870
rect 25563 4868 25569 4870
rect 25261 4859 25569 4868
rect 20628 4684 20680 4690
rect 20628 4626 20680 4632
rect 21272 4684 21324 4690
rect 21272 4626 21324 4632
rect 20444 4616 20496 4622
rect 20444 4558 20496 4564
rect 20456 4146 20484 4558
rect 20444 4140 20496 4146
rect 20444 4082 20496 4088
rect 18696 4004 18748 4010
rect 18696 3946 18748 3952
rect 18315 3836 18623 3845
rect 18315 3834 18321 3836
rect 18377 3834 18401 3836
rect 18457 3834 18481 3836
rect 18537 3834 18561 3836
rect 18617 3834 18623 3836
rect 18377 3782 18379 3834
rect 18559 3782 18561 3834
rect 18315 3780 18321 3782
rect 18377 3780 18401 3782
rect 18457 3780 18481 3782
rect 18537 3780 18561 3782
rect 18617 3780 18623 3782
rect 18315 3771 18623 3780
rect 18052 3732 18104 3738
rect 18052 3674 18104 3680
rect 18708 3670 18736 3946
rect 18696 3664 18748 3670
rect 18696 3606 18748 3612
rect 17408 3528 17460 3534
rect 17408 3470 17460 3476
rect 17500 3528 17552 3534
rect 17500 3470 17552 3476
rect 19248 3528 19300 3534
rect 19248 3470 19300 3476
rect 17420 2582 17448 3470
rect 17408 2576 17460 2582
rect 17408 2518 17460 2524
rect 17224 2508 17276 2514
rect 17224 2450 17276 2456
rect 17512 1986 17540 3470
rect 19260 3058 19288 3470
rect 19432 3392 19484 3398
rect 19432 3334 19484 3340
rect 19444 3126 19472 3334
rect 19432 3120 19484 3126
rect 19432 3062 19484 3068
rect 19248 3052 19300 3058
rect 19248 2994 19300 3000
rect 19984 2984 20036 2990
rect 19984 2926 20036 2932
rect 18315 2748 18623 2757
rect 18315 2746 18321 2748
rect 18377 2746 18401 2748
rect 18457 2746 18481 2748
rect 18537 2746 18561 2748
rect 18617 2746 18623 2748
rect 18377 2694 18379 2746
rect 18559 2694 18561 2746
rect 18315 2692 18321 2694
rect 18377 2692 18401 2694
rect 18457 2692 18481 2694
rect 18537 2692 18561 2694
rect 18617 2692 18623 2694
rect 18315 2683 18623 2692
rect 18052 2508 18104 2514
rect 18052 2450 18104 2456
rect 17420 1958 17540 1986
rect 17420 800 17448 1958
rect 18064 800 18092 2450
rect 19996 800 20024 2926
rect 21284 800 21312 4626
rect 21788 4380 22096 4389
rect 21788 4378 21794 4380
rect 21850 4378 21874 4380
rect 21930 4378 21954 4380
rect 22010 4378 22034 4380
rect 22090 4378 22096 4380
rect 21850 4326 21852 4378
rect 22032 4326 22034 4378
rect 21788 4324 21794 4326
rect 21850 4324 21874 4326
rect 21930 4324 21954 4326
rect 22010 4324 22034 4326
rect 22090 4324 22096 4326
rect 21788 4315 22096 4324
rect 25261 3836 25569 3845
rect 25261 3834 25267 3836
rect 25323 3834 25347 3836
rect 25403 3834 25427 3836
rect 25483 3834 25507 3836
rect 25563 3834 25569 3836
rect 25323 3782 25325 3834
rect 25505 3782 25507 3834
rect 25261 3780 25267 3782
rect 25323 3780 25347 3782
rect 25403 3780 25427 3782
rect 25483 3780 25507 3782
rect 25563 3780 25569 3782
rect 25261 3771 25569 3780
rect 25700 3738 25728 7822
rect 26160 7342 26188 8191
rect 26424 7744 26476 7750
rect 26424 7686 26476 7692
rect 26436 7478 26464 7686
rect 26424 7472 26476 7478
rect 26424 7414 26476 7420
rect 26620 7410 26648 8230
rect 26700 7812 26752 7818
rect 26700 7754 26752 7760
rect 26608 7404 26660 7410
rect 26608 7346 26660 7352
rect 26148 7336 26200 7342
rect 26148 7278 26200 7284
rect 26424 6860 26476 6866
rect 26424 6802 26476 6808
rect 25780 6792 25832 6798
rect 25780 6734 25832 6740
rect 25792 4622 25820 6734
rect 26436 6322 26464 6802
rect 26712 6458 26740 7754
rect 26988 6914 27016 12786
rect 27080 11762 27108 23666
rect 27264 22642 27292 31726
rect 27344 31272 27396 31278
rect 27344 31214 27396 31220
rect 27356 25770 27384 31214
rect 27448 30802 27476 32263
rect 27436 30796 27488 30802
rect 27436 30738 27488 30744
rect 27540 30705 27568 32914
rect 27526 30696 27582 30705
rect 27526 30631 27582 30640
rect 27528 29708 27580 29714
rect 27528 29650 27580 29656
rect 27540 28665 27568 29650
rect 27526 28656 27582 28665
rect 27526 28591 27582 28600
rect 27526 27568 27582 27577
rect 27526 27503 27528 27512
rect 27580 27503 27582 27512
rect 27528 27474 27580 27480
rect 27632 26994 27660 35866
rect 27712 31952 27764 31958
rect 27712 31894 27764 31900
rect 27724 31346 27752 31894
rect 27712 31340 27764 31346
rect 27712 31282 27764 31288
rect 27712 29572 27764 29578
rect 27712 29514 27764 29520
rect 27724 29306 27752 29514
rect 27712 29300 27764 29306
rect 27712 29242 27764 29248
rect 27620 26988 27672 26994
rect 27620 26930 27672 26936
rect 27344 25764 27396 25770
rect 27344 25706 27396 25712
rect 27528 25356 27580 25362
rect 27528 25298 27580 25304
rect 27540 25265 27568 25298
rect 27526 25256 27582 25265
rect 27526 25191 27582 25200
rect 27436 24812 27488 24818
rect 27436 24754 27488 24760
rect 27448 24410 27476 24754
rect 27436 24404 27488 24410
rect 27436 24346 27488 24352
rect 27344 24132 27396 24138
rect 27344 24074 27396 24080
rect 27356 22778 27384 24074
rect 27436 23520 27488 23526
rect 27436 23462 27488 23468
rect 27448 23254 27476 23462
rect 27436 23248 27488 23254
rect 27436 23190 27488 23196
rect 27344 22772 27396 22778
rect 27344 22714 27396 22720
rect 27252 22636 27304 22642
rect 27252 22578 27304 22584
rect 27160 15904 27212 15910
rect 27160 15846 27212 15852
rect 27172 15502 27200 15846
rect 27160 15496 27212 15502
rect 27160 15438 27212 15444
rect 27264 12434 27292 22578
rect 27528 22092 27580 22098
rect 27632 22094 27660 26930
rect 27632 22066 27752 22094
rect 27528 22034 27580 22040
rect 27540 21185 27568 22034
rect 27620 21412 27672 21418
rect 27620 21354 27672 21360
rect 27526 21176 27582 21185
rect 27526 21111 27582 21120
rect 27528 21004 27580 21010
rect 27528 20946 27580 20952
rect 27540 20505 27568 20946
rect 27526 20496 27582 20505
rect 27526 20431 27582 20440
rect 27632 18290 27660 21354
rect 27620 18284 27672 18290
rect 27620 18226 27672 18232
rect 27344 15360 27396 15366
rect 27344 15302 27396 15308
rect 27436 15360 27488 15366
rect 27436 15302 27488 15308
rect 27356 15162 27384 15302
rect 27344 15156 27396 15162
rect 27344 15098 27396 15104
rect 27448 15026 27476 15302
rect 27436 15020 27488 15026
rect 27436 14962 27488 14968
rect 27344 14952 27396 14958
rect 27344 14894 27396 14900
rect 27356 12782 27384 14894
rect 27344 12776 27396 12782
rect 27344 12718 27396 12724
rect 27264 12406 27384 12434
rect 27068 11756 27120 11762
rect 27068 11698 27120 11704
rect 27356 9586 27384 12406
rect 27448 10606 27476 14962
rect 27528 14476 27580 14482
rect 27528 14418 27580 14424
rect 27540 14385 27568 14418
rect 27526 14376 27582 14385
rect 27526 14311 27582 14320
rect 27632 12850 27660 18226
rect 27620 12844 27672 12850
rect 27620 12786 27672 12792
rect 27436 10600 27488 10606
rect 27436 10542 27488 10548
rect 27526 10296 27582 10305
rect 27526 10231 27582 10240
rect 27540 10130 27568 10231
rect 27528 10124 27580 10130
rect 27528 10066 27580 10072
rect 27344 9580 27396 9586
rect 27344 9522 27396 9528
rect 27620 9580 27672 9586
rect 27620 9522 27672 9528
rect 27252 8900 27304 8906
rect 27252 8842 27304 8848
rect 27264 8634 27292 8842
rect 27252 8628 27304 8634
rect 27252 8570 27304 8576
rect 27160 7200 27212 7206
rect 27160 7142 27212 7148
rect 26988 6886 27108 6914
rect 26700 6452 26752 6458
rect 26700 6394 26752 6400
rect 26424 6316 26476 6322
rect 26424 6258 26476 6264
rect 25780 4616 25832 4622
rect 25780 4558 25832 4564
rect 26516 4616 26568 4622
rect 26516 4558 26568 4564
rect 25792 4078 25820 4558
rect 25872 4480 25924 4486
rect 25872 4422 25924 4428
rect 25780 4072 25832 4078
rect 25780 4014 25832 4020
rect 25688 3732 25740 3738
rect 25688 3674 25740 3680
rect 25884 3602 25912 4422
rect 26148 4072 26200 4078
rect 26148 4014 26200 4020
rect 26424 4072 26476 4078
rect 26424 4014 26476 4020
rect 25872 3596 25924 3602
rect 25872 3538 25924 3544
rect 21548 3528 21600 3534
rect 21548 3470 21600 3476
rect 23848 3528 23900 3534
rect 23848 3470 23900 3476
rect 24308 3528 24360 3534
rect 26160 3505 26188 4014
rect 26436 3738 26464 4014
rect 26424 3732 26476 3738
rect 26424 3674 26476 3680
rect 24308 3470 24360 3476
rect 26146 3496 26202 3505
rect 21560 3058 21588 3470
rect 22192 3392 22244 3398
rect 22192 3334 22244 3340
rect 21788 3292 22096 3301
rect 21788 3290 21794 3292
rect 21850 3290 21874 3292
rect 21930 3290 21954 3292
rect 22010 3290 22034 3292
rect 22090 3290 22096 3292
rect 21850 3238 21852 3290
rect 22032 3238 22034 3290
rect 21788 3236 21794 3238
rect 21850 3236 21874 3238
rect 21930 3236 21954 3238
rect 22010 3236 22034 3238
rect 22090 3236 22096 3238
rect 21788 3227 22096 3236
rect 22204 3126 22232 3334
rect 22192 3120 22244 3126
rect 22192 3062 22244 3068
rect 21548 3052 21600 3058
rect 21548 2994 21600 3000
rect 21640 2916 21692 2922
rect 21640 2858 21692 2864
rect 21652 1714 21680 2858
rect 23860 2650 23888 3470
rect 24320 3058 24348 3470
rect 26146 3431 26202 3440
rect 24492 3392 24544 3398
rect 24492 3334 24544 3340
rect 24504 3126 24532 3334
rect 24492 3120 24544 3126
rect 24492 3062 24544 3068
rect 26528 3058 26556 4558
rect 26700 4548 26752 4554
rect 26700 4490 26752 4496
rect 26712 4282 26740 4490
rect 26700 4276 26752 4282
rect 26700 4218 26752 4224
rect 24308 3052 24360 3058
rect 24308 2994 24360 3000
rect 26516 3052 26568 3058
rect 26516 2994 26568 3000
rect 25136 2984 25188 2990
rect 25136 2926 25188 2932
rect 23848 2644 23900 2650
rect 23848 2586 23900 2592
rect 21788 2204 22096 2213
rect 21788 2202 21794 2204
rect 21850 2202 21874 2204
rect 21930 2202 21954 2204
rect 22010 2202 22034 2204
rect 22090 2202 22096 2204
rect 21850 2150 21852 2202
rect 22032 2150 22034 2202
rect 21788 2148 21794 2150
rect 21850 2148 21874 2150
rect 21930 2148 21954 2150
rect 22010 2148 22034 2150
rect 22090 2148 22096 2150
rect 21788 2139 22096 2148
rect 21652 1686 21956 1714
rect 21928 800 21956 1686
rect 25148 800 25176 2926
rect 26424 2848 26476 2854
rect 26146 2816 26202 2825
rect 26424 2790 26476 2796
rect 25261 2748 25569 2757
rect 26146 2751 26202 2760
rect 25261 2746 25267 2748
rect 25323 2746 25347 2748
rect 25403 2746 25427 2748
rect 25483 2746 25507 2748
rect 25563 2746 25569 2748
rect 25323 2694 25325 2746
rect 25505 2694 25507 2746
rect 25261 2692 25267 2694
rect 25323 2692 25347 2694
rect 25403 2692 25427 2694
rect 25483 2692 25507 2694
rect 25563 2692 25569 2694
rect 25261 2683 25569 2692
rect 26160 2514 26188 2751
rect 26436 2514 26464 2790
rect 27080 2650 27108 6886
rect 27172 6866 27200 7142
rect 27160 6860 27212 6866
rect 27160 6802 27212 6808
rect 27528 5772 27580 5778
rect 27528 5714 27580 5720
rect 27540 5273 27568 5714
rect 27526 5264 27582 5273
rect 27526 5199 27582 5208
rect 27528 4684 27580 4690
rect 27528 4626 27580 4632
rect 27436 3460 27488 3466
rect 27436 3402 27488 3408
rect 27068 2644 27120 2650
rect 27068 2586 27120 2592
rect 27448 2553 27476 3402
rect 27434 2544 27490 2553
rect 26148 2508 26200 2514
rect 26148 2450 26200 2456
rect 26424 2508 26476 2514
rect 27434 2479 27490 2488
rect 26424 2450 26476 2456
rect 27068 2440 27120 2446
rect 27068 2382 27120 2388
rect 27080 800 27108 2382
rect 27540 1465 27568 4626
rect 27632 4146 27660 9522
rect 27724 7954 27752 22066
rect 27816 8362 27844 36722
rect 27896 34944 27948 34950
rect 27896 34886 27948 34892
rect 27908 29170 27936 34886
rect 28000 32434 28028 37810
rect 28356 37256 28408 37262
rect 28356 37198 28408 37204
rect 28368 36378 28396 37198
rect 28734 37020 29042 37029
rect 28734 37018 28740 37020
rect 28796 37018 28820 37020
rect 28876 37018 28900 37020
rect 28956 37018 28980 37020
rect 29036 37018 29042 37020
rect 28796 36966 28798 37018
rect 28978 36966 28980 37018
rect 28734 36964 28740 36966
rect 28796 36964 28820 36966
rect 28876 36964 28900 36966
rect 28956 36964 28980 36966
rect 29036 36964 29042 36966
rect 28734 36955 29042 36964
rect 28356 36372 28408 36378
rect 28356 36314 28408 36320
rect 28734 35932 29042 35941
rect 28734 35930 28740 35932
rect 28796 35930 28820 35932
rect 28876 35930 28900 35932
rect 28956 35930 28980 35932
rect 29036 35930 29042 35932
rect 28796 35878 28798 35930
rect 28978 35878 28980 35930
rect 28734 35876 28740 35878
rect 28796 35876 28820 35878
rect 28876 35876 28900 35878
rect 28956 35876 28980 35878
rect 29036 35876 29042 35878
rect 28734 35867 29042 35876
rect 28734 34844 29042 34853
rect 28734 34842 28740 34844
rect 28796 34842 28820 34844
rect 28876 34842 28900 34844
rect 28956 34842 28980 34844
rect 29036 34842 29042 34844
rect 28796 34790 28798 34842
rect 28978 34790 28980 34842
rect 28734 34788 28740 34790
rect 28796 34788 28820 34790
rect 28876 34788 28900 34790
rect 28956 34788 28980 34790
rect 29036 34788 29042 34790
rect 28734 34779 29042 34788
rect 28734 33756 29042 33765
rect 28734 33754 28740 33756
rect 28796 33754 28820 33756
rect 28876 33754 28900 33756
rect 28956 33754 28980 33756
rect 29036 33754 29042 33756
rect 28796 33702 28798 33754
rect 28978 33702 28980 33754
rect 28734 33700 28740 33702
rect 28796 33700 28820 33702
rect 28876 33700 28900 33702
rect 28956 33700 28980 33702
rect 29036 33700 29042 33702
rect 28734 33691 29042 33700
rect 28172 33516 28224 33522
rect 28172 33458 28224 33464
rect 28080 32836 28132 32842
rect 28080 32778 28132 32784
rect 28092 32570 28120 32778
rect 28080 32564 28132 32570
rect 28080 32506 28132 32512
rect 28184 32450 28212 33458
rect 28264 33312 28316 33318
rect 28264 33254 28316 33260
rect 27988 32428 28040 32434
rect 27988 32370 28040 32376
rect 28092 32422 28212 32450
rect 27896 29164 27948 29170
rect 27896 29106 27948 29112
rect 27896 27396 27948 27402
rect 27896 27338 27948 27344
rect 27908 27130 27936 27338
rect 27896 27124 27948 27130
rect 27896 27066 27948 27072
rect 27896 24268 27948 24274
rect 27896 24210 27948 24216
rect 27908 22642 27936 24210
rect 27896 22636 27948 22642
rect 27896 22578 27948 22584
rect 28000 22094 28028 32370
rect 28092 24818 28120 32422
rect 28172 31136 28224 31142
rect 28172 31078 28224 31084
rect 28184 30802 28212 31078
rect 28276 30870 28304 33254
rect 28734 32668 29042 32677
rect 28734 32666 28740 32668
rect 28796 32666 28820 32668
rect 28876 32666 28900 32668
rect 28956 32666 28980 32668
rect 29036 32666 29042 32668
rect 28796 32614 28798 32666
rect 28978 32614 28980 32666
rect 28734 32612 28740 32614
rect 28796 32612 28820 32614
rect 28876 32612 28900 32614
rect 28956 32612 28980 32614
rect 29036 32612 29042 32614
rect 28734 32603 29042 32612
rect 28354 32056 28410 32065
rect 28354 31991 28410 32000
rect 28368 31890 28396 31991
rect 28356 31884 28408 31890
rect 28356 31826 28408 31832
rect 28734 31580 29042 31589
rect 28734 31578 28740 31580
rect 28796 31578 28820 31580
rect 28876 31578 28900 31580
rect 28956 31578 28980 31580
rect 29036 31578 29042 31580
rect 28796 31526 28798 31578
rect 28978 31526 28980 31578
rect 28734 31524 28740 31526
rect 28796 31524 28820 31526
rect 28876 31524 28900 31526
rect 28956 31524 28980 31526
rect 29036 31524 29042 31526
rect 28734 31515 29042 31524
rect 28356 31340 28408 31346
rect 28356 31282 28408 31288
rect 28368 30938 28396 31282
rect 28356 30932 28408 30938
rect 28356 30874 28408 30880
rect 28264 30864 28316 30870
rect 28264 30806 28316 30812
rect 28172 30796 28224 30802
rect 28172 30738 28224 30744
rect 28368 30682 28396 30874
rect 28276 30654 28396 30682
rect 28172 27872 28224 27878
rect 28172 27814 28224 27820
rect 28184 27538 28212 27814
rect 28172 27532 28224 27538
rect 28172 27474 28224 27480
rect 28172 25220 28224 25226
rect 28172 25162 28224 25168
rect 28184 24954 28212 25162
rect 28172 24948 28224 24954
rect 28172 24890 28224 24896
rect 28080 24812 28132 24818
rect 28080 24754 28132 24760
rect 28000 22066 28120 22094
rect 28092 20992 28120 22066
rect 28172 21956 28224 21962
rect 28172 21898 28224 21904
rect 28184 21690 28212 21898
rect 28172 21684 28224 21690
rect 28172 21626 28224 21632
rect 28276 21554 28304 30654
rect 28734 30492 29042 30501
rect 28734 30490 28740 30492
rect 28796 30490 28820 30492
rect 28876 30490 28900 30492
rect 28956 30490 28980 30492
rect 29036 30490 29042 30492
rect 28796 30438 28798 30490
rect 28978 30438 28980 30490
rect 28734 30436 28740 30438
rect 28796 30436 28820 30438
rect 28876 30436 28900 30438
rect 28956 30436 28980 30438
rect 29036 30436 29042 30438
rect 28734 30427 29042 30436
rect 28356 30048 28408 30054
rect 28356 29990 28408 29996
rect 28368 29714 28396 29990
rect 28356 29708 28408 29714
rect 28356 29650 28408 29656
rect 28734 29404 29042 29413
rect 28734 29402 28740 29404
rect 28796 29402 28820 29404
rect 28876 29402 28900 29404
rect 28956 29402 28980 29404
rect 29036 29402 29042 29404
rect 28796 29350 28798 29402
rect 28978 29350 28980 29402
rect 28734 29348 28740 29350
rect 28796 29348 28820 29350
rect 28876 29348 28900 29350
rect 28956 29348 28980 29350
rect 29036 29348 29042 29350
rect 28734 29339 29042 29348
rect 28734 28316 29042 28325
rect 28734 28314 28740 28316
rect 28796 28314 28820 28316
rect 28876 28314 28900 28316
rect 28956 28314 28980 28316
rect 29036 28314 29042 28316
rect 28796 28262 28798 28314
rect 28978 28262 28980 28314
rect 28734 28260 28740 28262
rect 28796 28260 28820 28262
rect 28876 28260 28900 28262
rect 28956 28260 28980 28262
rect 29036 28260 29042 28262
rect 28734 28251 29042 28260
rect 28734 27228 29042 27237
rect 28734 27226 28740 27228
rect 28796 27226 28820 27228
rect 28876 27226 28900 27228
rect 28956 27226 28980 27228
rect 29036 27226 29042 27228
rect 28796 27174 28798 27226
rect 28978 27174 28980 27226
rect 28734 27172 28740 27174
rect 28796 27172 28820 27174
rect 28876 27172 28900 27174
rect 28956 27172 28980 27174
rect 29036 27172 29042 27174
rect 28734 27163 29042 27172
rect 28354 26616 28410 26625
rect 28354 26551 28410 26560
rect 28368 26450 28396 26551
rect 28356 26444 28408 26450
rect 28356 26386 28408 26392
rect 28734 26140 29042 26149
rect 28734 26138 28740 26140
rect 28796 26138 28820 26140
rect 28876 26138 28900 26140
rect 28956 26138 28980 26140
rect 29036 26138 29042 26140
rect 28796 26086 28798 26138
rect 28978 26086 28980 26138
rect 28734 26084 28740 26086
rect 28796 26084 28820 26086
rect 28876 26084 28900 26086
rect 28956 26084 28980 26086
rect 29036 26084 29042 26086
rect 28734 26075 29042 26084
rect 28356 25696 28408 25702
rect 28356 25638 28408 25644
rect 28368 25362 28396 25638
rect 28356 25356 28408 25362
rect 28356 25298 28408 25304
rect 28734 25052 29042 25061
rect 28734 25050 28740 25052
rect 28796 25050 28820 25052
rect 28876 25050 28900 25052
rect 28956 25050 28980 25052
rect 29036 25050 29042 25052
rect 28796 24998 28798 25050
rect 28978 24998 28980 25050
rect 28734 24996 28740 24998
rect 28796 24996 28820 24998
rect 28876 24996 28900 24998
rect 28956 24996 28980 24998
rect 29036 24996 29042 24998
rect 28734 24987 29042 24996
rect 28354 24576 28410 24585
rect 28354 24511 28410 24520
rect 28368 24274 28396 24511
rect 28356 24268 28408 24274
rect 28356 24210 28408 24216
rect 28734 23964 29042 23973
rect 28734 23962 28740 23964
rect 28796 23962 28820 23964
rect 28876 23962 28900 23964
rect 28956 23962 28980 23964
rect 29036 23962 29042 23964
rect 28796 23910 28798 23962
rect 28978 23910 28980 23962
rect 28734 23908 28740 23910
rect 28796 23908 28820 23910
rect 28876 23908 28900 23910
rect 28956 23908 28980 23910
rect 29036 23908 29042 23910
rect 28734 23899 29042 23908
rect 29918 23896 29974 23905
rect 29918 23831 29974 23840
rect 29932 23186 29960 23831
rect 29920 23180 29972 23186
rect 29920 23122 29972 23128
rect 28734 22876 29042 22885
rect 28734 22874 28740 22876
rect 28796 22874 28820 22876
rect 28876 22874 28900 22876
rect 28956 22874 28980 22876
rect 29036 22874 29042 22876
rect 28796 22822 28798 22874
rect 28978 22822 28980 22874
rect 28734 22820 28740 22822
rect 28796 22820 28820 22822
rect 28876 22820 28900 22822
rect 28956 22820 28980 22822
rect 29036 22820 29042 22822
rect 28734 22811 29042 22820
rect 28356 22024 28408 22030
rect 28356 21966 28408 21972
rect 28368 21622 28396 21966
rect 28734 21788 29042 21797
rect 28734 21786 28740 21788
rect 28796 21786 28820 21788
rect 28876 21786 28900 21788
rect 28956 21786 28980 21788
rect 29036 21786 29042 21788
rect 28796 21734 28798 21786
rect 28978 21734 28980 21786
rect 28734 21732 28740 21734
rect 28796 21732 28820 21734
rect 28876 21732 28900 21734
rect 28956 21732 28980 21734
rect 29036 21732 29042 21734
rect 28734 21723 29042 21732
rect 28356 21616 28408 21622
rect 28356 21558 28408 21564
rect 28264 21548 28316 21554
rect 28264 21490 28316 21496
rect 28092 20964 28304 20992
rect 28172 20868 28224 20874
rect 28172 20810 28224 20816
rect 28184 20602 28212 20810
rect 28172 20596 28224 20602
rect 28172 20538 28224 20544
rect 28080 20460 28132 20466
rect 28080 20402 28132 20408
rect 27896 19848 27948 19854
rect 27896 19790 27948 19796
rect 27908 17814 27936 19790
rect 27988 18692 28040 18698
rect 27988 18634 28040 18640
rect 28000 18426 28028 18634
rect 27988 18420 28040 18426
rect 27988 18362 28040 18368
rect 27896 17808 27948 17814
rect 27896 17750 27948 17756
rect 27896 16992 27948 16998
rect 27896 16934 27948 16940
rect 27908 16726 27936 16934
rect 27896 16720 27948 16726
rect 27896 16662 27948 16668
rect 28092 15502 28120 20402
rect 28276 17202 28304 20964
rect 28356 20936 28408 20942
rect 28356 20878 28408 20884
rect 28368 20398 28396 20878
rect 28734 20700 29042 20709
rect 28734 20698 28740 20700
rect 28796 20698 28820 20700
rect 28876 20698 28900 20700
rect 28956 20698 28980 20700
rect 29036 20698 29042 20700
rect 28796 20646 28798 20698
rect 28978 20646 28980 20698
rect 28734 20644 28740 20646
rect 28796 20644 28820 20646
rect 28876 20644 28900 20646
rect 28956 20644 28980 20646
rect 29036 20644 29042 20646
rect 28734 20635 29042 20644
rect 28356 20392 28408 20398
rect 28356 20334 28408 20340
rect 28630 19816 28686 19825
rect 28630 19751 28686 19760
rect 28356 19168 28408 19174
rect 28356 19110 28408 19116
rect 28368 18834 28396 19110
rect 28356 18828 28408 18834
rect 28356 18770 28408 18776
rect 28644 17746 28672 19751
rect 28734 19612 29042 19621
rect 28734 19610 28740 19612
rect 28796 19610 28820 19612
rect 28876 19610 28900 19612
rect 28956 19610 28980 19612
rect 29036 19610 29042 19612
rect 28796 19558 28798 19610
rect 28978 19558 28980 19610
rect 28734 19556 28740 19558
rect 28796 19556 28820 19558
rect 28876 19556 28900 19558
rect 28956 19556 28980 19558
rect 29036 19556 29042 19558
rect 28734 19547 29042 19556
rect 28734 18524 29042 18533
rect 28734 18522 28740 18524
rect 28796 18522 28820 18524
rect 28876 18522 28900 18524
rect 28956 18522 28980 18524
rect 29036 18522 29042 18524
rect 28796 18470 28798 18522
rect 28978 18470 28980 18522
rect 28734 18468 28740 18470
rect 28796 18468 28820 18470
rect 28876 18468 28900 18470
rect 28956 18468 28980 18470
rect 29036 18468 29042 18470
rect 28734 18459 29042 18468
rect 28632 17740 28684 17746
rect 28632 17682 28684 17688
rect 28734 17436 29042 17445
rect 28734 17434 28740 17436
rect 28796 17434 28820 17436
rect 28876 17434 28900 17436
rect 28956 17434 28980 17436
rect 29036 17434 29042 17436
rect 28796 17382 28798 17434
rect 28978 17382 28980 17434
rect 28734 17380 28740 17382
rect 28796 17380 28820 17382
rect 28876 17380 28900 17382
rect 28956 17380 28980 17382
rect 29036 17380 29042 17382
rect 28734 17371 29042 17380
rect 28264 17196 28316 17202
rect 28264 17138 28316 17144
rect 28632 16516 28684 16522
rect 28632 16458 28684 16464
rect 28644 15745 28672 16458
rect 29918 16416 29974 16425
rect 28734 16348 29042 16357
rect 29918 16351 29974 16360
rect 28734 16346 28740 16348
rect 28796 16346 28820 16348
rect 28876 16346 28900 16348
rect 28956 16346 28980 16348
rect 29036 16346 29042 16348
rect 28796 16294 28798 16346
rect 28978 16294 28980 16346
rect 28734 16292 28740 16294
rect 28796 16292 28820 16294
rect 28876 16292 28900 16294
rect 28956 16292 28980 16294
rect 29036 16292 29042 16294
rect 28734 16283 29042 16292
rect 29932 16114 29960 16351
rect 29920 16108 29972 16114
rect 29920 16050 29972 16056
rect 28630 15736 28686 15745
rect 28630 15671 28686 15680
rect 28080 15496 28132 15502
rect 28080 15438 28132 15444
rect 27804 8356 27856 8362
rect 27804 8298 27856 8304
rect 27816 8242 27844 8298
rect 27816 8214 27936 8242
rect 27712 7948 27764 7954
rect 27712 7890 27764 7896
rect 27804 7744 27856 7750
rect 27804 7686 27856 7692
rect 27816 7410 27844 7686
rect 27804 7404 27856 7410
rect 27804 7346 27856 7352
rect 27620 4140 27672 4146
rect 27620 4082 27672 4088
rect 27632 3534 27660 4082
rect 27908 3534 27936 8214
rect 28092 6914 28120 15438
rect 28172 15360 28224 15366
rect 28172 15302 28224 15308
rect 28184 14482 28212 15302
rect 28734 15260 29042 15269
rect 28734 15258 28740 15260
rect 28796 15258 28820 15260
rect 28876 15258 28900 15260
rect 28956 15258 28980 15260
rect 29036 15258 29042 15260
rect 28796 15206 28798 15258
rect 28978 15206 28980 15258
rect 28734 15204 28740 15206
rect 28796 15204 28820 15206
rect 28876 15204 28900 15206
rect 28956 15204 28980 15206
rect 29036 15204 29042 15206
rect 28734 15195 29042 15204
rect 28172 14476 28224 14482
rect 28172 14418 28224 14424
rect 28356 14408 28408 14414
rect 28356 14350 28408 14356
rect 28368 13938 28396 14350
rect 28734 14172 29042 14181
rect 28734 14170 28740 14172
rect 28796 14170 28820 14172
rect 28876 14170 28900 14172
rect 28956 14170 28980 14172
rect 29036 14170 29042 14172
rect 28796 14118 28798 14170
rect 28978 14118 28980 14170
rect 28734 14116 28740 14118
rect 28796 14116 28820 14118
rect 28876 14116 28900 14118
rect 28956 14116 28980 14118
rect 29036 14116 29042 14118
rect 28734 14107 29042 14116
rect 28356 13932 28408 13938
rect 28356 13874 28408 13880
rect 28734 13084 29042 13093
rect 28734 13082 28740 13084
rect 28796 13082 28820 13084
rect 28876 13082 28900 13084
rect 28956 13082 28980 13084
rect 29036 13082 29042 13084
rect 28796 13030 28798 13082
rect 28978 13030 28980 13082
rect 28734 13028 28740 13030
rect 28796 13028 28820 13030
rect 28876 13028 28900 13030
rect 28956 13028 28980 13030
rect 29036 13028 29042 13030
rect 28734 13019 29042 13028
rect 28354 12336 28410 12345
rect 28354 12271 28356 12280
rect 28408 12271 28410 12280
rect 28356 12242 28408 12248
rect 28734 11996 29042 12005
rect 28734 11994 28740 11996
rect 28796 11994 28820 11996
rect 28876 11994 28900 11996
rect 28956 11994 28980 11996
rect 29036 11994 29042 11996
rect 28796 11942 28798 11994
rect 28978 11942 28980 11994
rect 28734 11940 28740 11942
rect 28796 11940 28820 11942
rect 28876 11940 28900 11942
rect 28956 11940 28980 11942
rect 29036 11940 29042 11942
rect 28734 11931 29042 11940
rect 29920 11076 29972 11082
rect 29920 11018 29972 11024
rect 29932 10985 29960 11018
rect 29918 10976 29974 10985
rect 28734 10908 29042 10917
rect 29918 10911 29974 10920
rect 28734 10906 28740 10908
rect 28796 10906 28820 10908
rect 28876 10906 28900 10908
rect 28956 10906 28980 10908
rect 29036 10906 29042 10908
rect 28796 10854 28798 10906
rect 28978 10854 28980 10906
rect 28734 10852 28740 10854
rect 28796 10852 28820 10854
rect 28876 10852 28900 10854
rect 28956 10852 28980 10854
rect 29036 10852 29042 10854
rect 28734 10843 29042 10852
rect 28356 10464 28408 10470
rect 28356 10406 28408 10412
rect 28368 10130 28396 10406
rect 28356 10124 28408 10130
rect 28356 10066 28408 10072
rect 28172 9988 28224 9994
rect 28172 9930 28224 9936
rect 28184 9722 28212 9930
rect 28734 9820 29042 9829
rect 28734 9818 28740 9820
rect 28796 9818 28820 9820
rect 28876 9818 28900 9820
rect 28956 9818 28980 9820
rect 29036 9818 29042 9820
rect 28796 9766 28798 9818
rect 28978 9766 28980 9818
rect 28734 9764 28740 9766
rect 28796 9764 28820 9766
rect 28876 9764 28900 9766
rect 28956 9764 28980 9766
rect 29036 9764 29042 9766
rect 28734 9755 29042 9764
rect 28172 9716 28224 9722
rect 28172 9658 28224 9664
rect 28356 8968 28408 8974
rect 28354 8936 28356 8945
rect 28408 8936 28410 8945
rect 28354 8871 28410 8880
rect 28734 8732 29042 8741
rect 28734 8730 28740 8732
rect 28796 8730 28820 8732
rect 28876 8730 28900 8732
rect 28956 8730 28980 8732
rect 29036 8730 29042 8732
rect 28796 8678 28798 8730
rect 28978 8678 28980 8730
rect 28734 8676 28740 8678
rect 28796 8676 28820 8678
rect 28876 8676 28900 8678
rect 28956 8676 28980 8678
rect 29036 8676 29042 8678
rect 28734 8667 29042 8676
rect 29920 7812 29972 7818
rect 29920 7754 29972 7760
rect 28734 7644 29042 7653
rect 28734 7642 28740 7644
rect 28796 7642 28820 7644
rect 28876 7642 28900 7644
rect 28956 7642 28980 7644
rect 29036 7642 29042 7644
rect 28796 7590 28798 7642
rect 28978 7590 28980 7642
rect 28734 7588 28740 7590
rect 28796 7588 28820 7590
rect 28876 7588 28900 7590
rect 28956 7588 28980 7590
rect 29036 7588 29042 7590
rect 28734 7579 29042 7588
rect 29932 7585 29960 7754
rect 29918 7576 29974 7585
rect 29918 7511 29974 7520
rect 28000 6886 28120 6914
rect 28354 6896 28410 6905
rect 28000 6322 28028 6886
rect 28354 6831 28356 6840
rect 28408 6831 28410 6840
rect 28356 6802 28408 6808
rect 28734 6556 29042 6565
rect 28734 6554 28740 6556
rect 28796 6554 28820 6556
rect 28876 6554 28900 6556
rect 28956 6554 28980 6556
rect 29036 6554 29042 6556
rect 28796 6502 28798 6554
rect 28978 6502 28980 6554
rect 28734 6500 28740 6502
rect 28796 6500 28820 6502
rect 28876 6500 28900 6502
rect 28956 6500 28980 6502
rect 29036 6500 29042 6502
rect 28734 6491 29042 6500
rect 27988 6316 28040 6322
rect 27988 6258 28040 6264
rect 28172 6112 28224 6118
rect 28172 6054 28224 6060
rect 28184 5778 28212 6054
rect 28172 5772 28224 5778
rect 28172 5714 28224 5720
rect 28356 5704 28408 5710
rect 28356 5646 28408 5652
rect 28368 5234 28396 5646
rect 28734 5468 29042 5477
rect 28734 5466 28740 5468
rect 28796 5466 28820 5468
rect 28876 5466 28900 5468
rect 28956 5466 28980 5468
rect 29036 5466 29042 5468
rect 28796 5414 28798 5466
rect 28978 5414 28980 5466
rect 28734 5412 28740 5414
rect 28796 5412 28820 5414
rect 28876 5412 28900 5414
rect 28956 5412 28980 5414
rect 29036 5412 29042 5414
rect 28734 5403 29042 5412
rect 28356 5228 28408 5234
rect 28356 5170 28408 5176
rect 28734 4380 29042 4389
rect 28734 4378 28740 4380
rect 28796 4378 28820 4380
rect 28876 4378 28900 4380
rect 28956 4378 28980 4380
rect 29036 4378 29042 4380
rect 28796 4326 28798 4378
rect 28978 4326 28980 4378
rect 28734 4324 28740 4326
rect 28796 4324 28820 4326
rect 28876 4324 28900 4326
rect 28956 4324 28980 4326
rect 29036 4324 29042 4326
rect 28734 4315 29042 4324
rect 27620 3528 27672 3534
rect 27620 3470 27672 3476
rect 27896 3528 27948 3534
rect 27896 3470 27948 3476
rect 27908 3058 27936 3470
rect 28734 3292 29042 3301
rect 28734 3290 28740 3292
rect 28796 3290 28820 3292
rect 28876 3290 28900 3292
rect 28956 3290 28980 3292
rect 29036 3290 29042 3292
rect 28796 3238 28798 3290
rect 28978 3238 28980 3290
rect 28734 3236 28740 3238
rect 28796 3236 28820 3238
rect 28876 3236 28900 3238
rect 28956 3236 28980 3238
rect 29036 3236 29042 3238
rect 28734 3227 29042 3236
rect 27896 3052 27948 3058
rect 27896 2994 27948 3000
rect 28734 2204 29042 2213
rect 28734 2202 28740 2204
rect 28796 2202 28820 2204
rect 28876 2202 28900 2204
rect 28956 2202 28980 2204
rect 29036 2202 29042 2204
rect 28796 2150 28798 2202
rect 28978 2150 28980 2202
rect 28734 2148 28740 2150
rect 28796 2148 28820 2150
rect 28876 2148 28900 2150
rect 28956 2148 28980 2150
rect 29036 2148 29042 2150
rect 28734 2139 29042 2148
rect 27526 1456 27582 1465
rect 27526 1391 27582 1400
rect -10 200 102 800
rect 634 200 746 800
rect 1278 200 1390 800
rect 1922 200 2034 800
rect 2566 200 2678 800
rect 3210 200 3322 800
rect 3854 200 3966 800
rect 4498 200 4610 800
rect 5786 200 5898 800
rect 6430 200 6542 800
rect 7074 200 7186 800
rect 7718 200 7830 800
rect 8362 200 8474 800
rect 9006 200 9118 800
rect 9650 200 9762 800
rect 10938 200 11050 800
rect 11582 200 11694 800
rect 12226 200 12338 800
rect 12870 200 12982 800
rect 13514 200 13626 800
rect 14158 200 14270 800
rect 14802 200 14914 800
rect 16090 200 16202 800
rect 16734 200 16846 800
rect 17378 200 17490 800
rect 18022 200 18134 800
rect 18666 200 18778 800
rect 19310 200 19422 800
rect 19954 200 20066 800
rect 21242 200 21354 800
rect 21886 200 21998 800
rect 22530 200 22642 800
rect 23174 200 23286 800
rect 23818 200 23930 800
rect 24462 200 24574 800
rect 25106 200 25218 800
rect 26394 200 26506 800
rect 27038 200 27150 800
rect 27682 200 27794 800
rect 28326 200 28438 800
rect 28970 200 29082 800
rect 29614 200 29726 800
<< via2 >>
rect 2962 49680 3018 49736
rect 4429 47354 4485 47356
rect 4509 47354 4565 47356
rect 4589 47354 4645 47356
rect 4669 47354 4725 47356
rect 4429 47302 4475 47354
rect 4475 47302 4485 47354
rect 4509 47302 4539 47354
rect 4539 47302 4551 47354
rect 4551 47302 4565 47354
rect 4589 47302 4603 47354
rect 4603 47302 4615 47354
rect 4615 47302 4645 47354
rect 4669 47302 4679 47354
rect 4679 47302 4725 47354
rect 4429 47300 4485 47302
rect 4509 47300 4565 47302
rect 4589 47300 4645 47302
rect 4669 47300 4725 47302
rect 4429 46266 4485 46268
rect 4509 46266 4565 46268
rect 4589 46266 4645 46268
rect 4669 46266 4725 46268
rect 4429 46214 4475 46266
rect 4475 46214 4485 46266
rect 4509 46214 4539 46266
rect 4539 46214 4551 46266
rect 4551 46214 4565 46266
rect 4589 46214 4603 46266
rect 4603 46214 4615 46266
rect 4615 46214 4645 46266
rect 4669 46214 4679 46266
rect 4679 46214 4725 46266
rect 4429 46212 4485 46214
rect 4509 46212 4565 46214
rect 4589 46212 4645 46214
rect 4669 46212 4725 46214
rect 1582 42200 1638 42256
rect 1674 37440 1730 37496
rect 4429 45178 4485 45180
rect 4509 45178 4565 45180
rect 4589 45178 4645 45180
rect 4669 45178 4725 45180
rect 4429 45126 4475 45178
rect 4475 45126 4485 45178
rect 4509 45126 4539 45178
rect 4539 45126 4551 45178
rect 4551 45126 4565 45178
rect 4589 45126 4603 45178
rect 4603 45126 4615 45178
rect 4615 45126 4645 45178
rect 4669 45126 4679 45178
rect 4679 45126 4725 45178
rect 4429 45124 4485 45126
rect 4509 45124 4565 45126
rect 4589 45124 4645 45126
rect 4669 45124 4725 45126
rect 4250 44920 4306 44976
rect 3606 44276 3608 44296
rect 3608 44276 3660 44296
rect 3660 44276 3662 44296
rect 3606 44240 3662 44276
rect 1674 36080 1730 36136
rect 1582 29960 1638 30016
rect 1582 27920 1638 27976
rect 1582 25236 1584 25256
rect 1584 25236 1636 25256
rect 1636 25236 1638 25256
rect 1582 25200 1638 25236
rect 1582 18400 1638 18456
rect 1582 14340 1638 14376
rect 1582 14320 1584 14340
rect 1584 14320 1636 14340
rect 1636 14320 1638 14340
rect 1582 13640 1638 13696
rect 2134 19080 2190 19136
rect 2778 41520 2834 41576
rect 2778 38800 2834 38856
rect 2870 36760 2926 36816
rect 4429 44090 4485 44092
rect 4509 44090 4565 44092
rect 4589 44090 4645 44092
rect 4669 44090 4725 44092
rect 4429 44038 4475 44090
rect 4475 44038 4485 44090
rect 4509 44038 4539 44090
rect 4539 44038 4551 44090
rect 4551 44038 4565 44090
rect 4589 44038 4603 44090
rect 4603 44038 4615 44090
rect 4615 44038 4645 44090
rect 4669 44038 4679 44090
rect 4679 44038 4725 44090
rect 4429 44036 4485 44038
rect 4509 44036 4565 44038
rect 4589 44036 4645 44038
rect 4669 44036 4725 44038
rect 4429 43002 4485 43004
rect 4509 43002 4565 43004
rect 4589 43002 4645 43004
rect 4669 43002 4725 43004
rect 4429 42950 4475 43002
rect 4475 42950 4485 43002
rect 4509 42950 4539 43002
rect 4539 42950 4551 43002
rect 4551 42950 4565 43002
rect 4589 42950 4603 43002
rect 4603 42950 4615 43002
rect 4615 42950 4645 43002
rect 4669 42950 4679 43002
rect 4679 42950 4725 43002
rect 4429 42948 4485 42950
rect 4509 42948 4565 42950
rect 4589 42948 4645 42950
rect 4669 42948 4725 42950
rect 4429 41914 4485 41916
rect 4509 41914 4565 41916
rect 4589 41914 4645 41916
rect 4669 41914 4725 41916
rect 4429 41862 4475 41914
rect 4475 41862 4485 41914
rect 4509 41862 4539 41914
rect 4539 41862 4551 41914
rect 4551 41862 4565 41914
rect 4589 41862 4603 41914
rect 4603 41862 4615 41914
rect 4615 41862 4645 41914
rect 4669 41862 4679 41914
rect 4679 41862 4725 41914
rect 4429 41860 4485 41862
rect 4509 41860 4565 41862
rect 4589 41860 4645 41862
rect 4669 41860 4725 41862
rect 4429 40826 4485 40828
rect 4509 40826 4565 40828
rect 4589 40826 4645 40828
rect 4669 40826 4725 40828
rect 4429 40774 4475 40826
rect 4475 40774 4485 40826
rect 4509 40774 4539 40826
rect 4539 40774 4551 40826
rect 4551 40774 4565 40826
rect 4589 40774 4603 40826
rect 4603 40774 4615 40826
rect 4615 40774 4645 40826
rect 4669 40774 4679 40826
rect 4679 40774 4725 40826
rect 4429 40772 4485 40774
rect 4509 40772 4565 40774
rect 4589 40772 4645 40774
rect 4669 40772 4725 40774
rect 4429 39738 4485 39740
rect 4509 39738 4565 39740
rect 4589 39738 4645 39740
rect 4669 39738 4725 39740
rect 4429 39686 4475 39738
rect 4475 39686 4485 39738
rect 4509 39686 4539 39738
rect 4539 39686 4551 39738
rect 4551 39686 4565 39738
rect 4589 39686 4603 39738
rect 4603 39686 4615 39738
rect 4615 39686 4645 39738
rect 4669 39686 4679 39738
rect 4679 39686 4725 39738
rect 4429 39684 4485 39686
rect 4509 39684 4565 39686
rect 4589 39684 4645 39686
rect 4669 39684 4725 39686
rect 4429 38650 4485 38652
rect 4509 38650 4565 38652
rect 4589 38650 4645 38652
rect 4669 38650 4725 38652
rect 4429 38598 4475 38650
rect 4475 38598 4485 38650
rect 4509 38598 4539 38650
rect 4539 38598 4551 38650
rect 4551 38598 4565 38650
rect 4589 38598 4603 38650
rect 4603 38598 4615 38650
rect 4615 38598 4645 38650
rect 4669 38598 4679 38650
rect 4679 38598 4725 38650
rect 4429 38596 4485 38598
rect 4509 38596 4565 38598
rect 4589 38596 4645 38598
rect 4669 38596 4725 38598
rect 4429 37562 4485 37564
rect 4509 37562 4565 37564
rect 4589 37562 4645 37564
rect 4669 37562 4725 37564
rect 4429 37510 4475 37562
rect 4475 37510 4485 37562
rect 4509 37510 4539 37562
rect 4539 37510 4551 37562
rect 4551 37510 4565 37562
rect 4589 37510 4603 37562
rect 4603 37510 4615 37562
rect 4615 37510 4645 37562
rect 4669 37510 4679 37562
rect 4679 37510 4725 37562
rect 4429 37508 4485 37510
rect 4509 37508 4565 37510
rect 4589 37508 4645 37510
rect 4669 37508 4725 37510
rect 2778 34720 2834 34776
rect 2778 32000 2834 32056
rect 2778 25880 2834 25936
rect 2778 19760 2834 19816
rect 1582 2760 1638 2816
rect 2778 17740 2834 17776
rect 2778 17720 2780 17740
rect 2780 17720 2832 17740
rect 2832 17720 2834 17740
rect 2778 15680 2834 15736
rect 3514 33380 3570 33416
rect 3514 33360 3516 33380
rect 3516 33360 3568 33380
rect 3568 33360 3570 33380
rect 2778 11636 2780 11656
rect 2780 11636 2832 11656
rect 2832 11636 2834 11656
rect 2778 11600 2834 11636
rect 3514 12280 3570 12336
rect 2778 8880 2834 8936
rect 2962 8200 3018 8256
rect 3054 7520 3110 7576
rect 3146 4800 3202 4856
rect 2778 4120 2834 4176
rect 2778 3440 2834 3496
rect 4429 36474 4485 36476
rect 4509 36474 4565 36476
rect 4589 36474 4645 36476
rect 4669 36474 4725 36476
rect 4429 36422 4475 36474
rect 4475 36422 4485 36474
rect 4509 36422 4539 36474
rect 4539 36422 4551 36474
rect 4551 36422 4565 36474
rect 4589 36422 4603 36474
rect 4603 36422 4615 36474
rect 4615 36422 4645 36474
rect 4669 36422 4679 36474
rect 4679 36422 4725 36474
rect 4429 36420 4485 36422
rect 4509 36420 4565 36422
rect 4589 36420 4645 36422
rect 4669 36420 4725 36422
rect 7902 46810 7958 46812
rect 7982 46810 8038 46812
rect 8062 46810 8118 46812
rect 8142 46810 8198 46812
rect 7902 46758 7948 46810
rect 7948 46758 7958 46810
rect 7982 46758 8012 46810
rect 8012 46758 8024 46810
rect 8024 46758 8038 46810
rect 8062 46758 8076 46810
rect 8076 46758 8088 46810
rect 8088 46758 8118 46810
rect 8142 46758 8152 46810
rect 8152 46758 8198 46810
rect 7902 46756 7958 46758
rect 7982 46756 8038 46758
rect 8062 46756 8118 46758
rect 8142 46756 8198 46758
rect 4429 35386 4485 35388
rect 4509 35386 4565 35388
rect 4589 35386 4645 35388
rect 4669 35386 4725 35388
rect 4429 35334 4475 35386
rect 4475 35334 4485 35386
rect 4509 35334 4539 35386
rect 4539 35334 4551 35386
rect 4551 35334 4565 35386
rect 4589 35334 4603 35386
rect 4603 35334 4615 35386
rect 4615 35334 4645 35386
rect 4669 35334 4679 35386
rect 4679 35334 4725 35386
rect 4429 35332 4485 35334
rect 4509 35332 4565 35334
rect 4589 35332 4645 35334
rect 4669 35332 4725 35334
rect 7902 45722 7958 45724
rect 7982 45722 8038 45724
rect 8062 45722 8118 45724
rect 8142 45722 8198 45724
rect 7902 45670 7948 45722
rect 7948 45670 7958 45722
rect 7982 45670 8012 45722
rect 8012 45670 8024 45722
rect 8024 45670 8038 45722
rect 8062 45670 8076 45722
rect 8076 45670 8088 45722
rect 8088 45670 8118 45722
rect 8142 45670 8152 45722
rect 8152 45670 8198 45722
rect 7902 45668 7958 45670
rect 7982 45668 8038 45670
rect 8062 45668 8118 45670
rect 8142 45668 8198 45670
rect 11375 47354 11431 47356
rect 11455 47354 11511 47356
rect 11535 47354 11591 47356
rect 11615 47354 11671 47356
rect 11375 47302 11421 47354
rect 11421 47302 11431 47354
rect 11455 47302 11485 47354
rect 11485 47302 11497 47354
rect 11497 47302 11511 47354
rect 11535 47302 11549 47354
rect 11549 47302 11561 47354
rect 11561 47302 11591 47354
rect 11615 47302 11625 47354
rect 11625 47302 11671 47354
rect 11375 47300 11431 47302
rect 11455 47300 11511 47302
rect 11535 47300 11591 47302
rect 11615 47300 11671 47302
rect 11375 46266 11431 46268
rect 11455 46266 11511 46268
rect 11535 46266 11591 46268
rect 11615 46266 11671 46268
rect 11375 46214 11421 46266
rect 11421 46214 11431 46266
rect 11455 46214 11485 46266
rect 11485 46214 11497 46266
rect 11497 46214 11511 46266
rect 11535 46214 11549 46266
rect 11549 46214 11561 46266
rect 11561 46214 11591 46266
rect 11615 46214 11625 46266
rect 11625 46214 11671 46266
rect 11375 46212 11431 46214
rect 11455 46212 11511 46214
rect 11535 46212 11591 46214
rect 11615 46212 11671 46214
rect 14848 46810 14904 46812
rect 14928 46810 14984 46812
rect 15008 46810 15064 46812
rect 15088 46810 15144 46812
rect 14848 46758 14894 46810
rect 14894 46758 14904 46810
rect 14928 46758 14958 46810
rect 14958 46758 14970 46810
rect 14970 46758 14984 46810
rect 15008 46758 15022 46810
rect 15022 46758 15034 46810
rect 15034 46758 15064 46810
rect 15088 46758 15098 46810
rect 15098 46758 15144 46810
rect 14848 46756 14904 46758
rect 14928 46756 14984 46758
rect 15008 46756 15064 46758
rect 15088 46756 15144 46758
rect 18321 47354 18377 47356
rect 18401 47354 18457 47356
rect 18481 47354 18537 47356
rect 18561 47354 18617 47356
rect 18321 47302 18367 47354
rect 18367 47302 18377 47354
rect 18401 47302 18431 47354
rect 18431 47302 18443 47354
rect 18443 47302 18457 47354
rect 18481 47302 18495 47354
rect 18495 47302 18507 47354
rect 18507 47302 18537 47354
rect 18561 47302 18571 47354
rect 18571 47302 18617 47354
rect 18321 47300 18377 47302
rect 18401 47300 18457 47302
rect 18481 47300 18537 47302
rect 18561 47300 18617 47302
rect 18321 46266 18377 46268
rect 18401 46266 18457 46268
rect 18481 46266 18537 46268
rect 18561 46266 18617 46268
rect 18321 46214 18367 46266
rect 18367 46214 18377 46266
rect 18401 46214 18431 46266
rect 18431 46214 18443 46266
rect 18443 46214 18457 46266
rect 18481 46214 18495 46266
rect 18495 46214 18507 46266
rect 18507 46214 18537 46266
rect 18561 46214 18571 46266
rect 18571 46214 18617 46266
rect 18321 46212 18377 46214
rect 18401 46212 18457 46214
rect 18481 46212 18537 46214
rect 18561 46212 18617 46214
rect 21794 46810 21850 46812
rect 21874 46810 21930 46812
rect 21954 46810 22010 46812
rect 22034 46810 22090 46812
rect 21794 46758 21840 46810
rect 21840 46758 21850 46810
rect 21874 46758 21904 46810
rect 21904 46758 21916 46810
rect 21916 46758 21930 46810
rect 21954 46758 21968 46810
rect 21968 46758 21980 46810
rect 21980 46758 22010 46810
rect 22034 46758 22044 46810
rect 22044 46758 22090 46810
rect 21794 46756 21850 46758
rect 21874 46756 21930 46758
rect 21954 46756 22010 46758
rect 22034 46756 22090 46758
rect 11375 45178 11431 45180
rect 11455 45178 11511 45180
rect 11535 45178 11591 45180
rect 11615 45178 11671 45180
rect 11375 45126 11421 45178
rect 11421 45126 11431 45178
rect 11455 45126 11485 45178
rect 11485 45126 11497 45178
rect 11497 45126 11511 45178
rect 11535 45126 11549 45178
rect 11549 45126 11561 45178
rect 11561 45126 11591 45178
rect 11615 45126 11625 45178
rect 11625 45126 11671 45178
rect 11375 45124 11431 45126
rect 11455 45124 11511 45126
rect 11535 45124 11591 45126
rect 11615 45124 11671 45126
rect 7902 44634 7958 44636
rect 7982 44634 8038 44636
rect 8062 44634 8118 44636
rect 8142 44634 8198 44636
rect 7902 44582 7948 44634
rect 7948 44582 7958 44634
rect 7982 44582 8012 44634
rect 8012 44582 8024 44634
rect 8024 44582 8038 44634
rect 8062 44582 8076 44634
rect 8076 44582 8088 44634
rect 8088 44582 8118 44634
rect 8142 44582 8152 44634
rect 8152 44582 8198 44634
rect 7902 44580 7958 44582
rect 7982 44580 8038 44582
rect 8062 44580 8118 44582
rect 8142 44580 8198 44582
rect 11375 44090 11431 44092
rect 11455 44090 11511 44092
rect 11535 44090 11591 44092
rect 11615 44090 11671 44092
rect 11375 44038 11421 44090
rect 11421 44038 11431 44090
rect 11455 44038 11485 44090
rect 11485 44038 11497 44090
rect 11497 44038 11511 44090
rect 11535 44038 11549 44090
rect 11549 44038 11561 44090
rect 11561 44038 11591 44090
rect 11615 44038 11625 44090
rect 11625 44038 11671 44090
rect 11375 44036 11431 44038
rect 11455 44036 11511 44038
rect 11535 44036 11591 44038
rect 11615 44036 11671 44038
rect 7902 43546 7958 43548
rect 7982 43546 8038 43548
rect 8062 43546 8118 43548
rect 8142 43546 8198 43548
rect 7902 43494 7948 43546
rect 7948 43494 7958 43546
rect 7982 43494 8012 43546
rect 8012 43494 8024 43546
rect 8024 43494 8038 43546
rect 8062 43494 8076 43546
rect 8076 43494 8088 43546
rect 8088 43494 8118 43546
rect 8142 43494 8152 43546
rect 8152 43494 8198 43546
rect 7902 43492 7958 43494
rect 7982 43492 8038 43494
rect 8062 43492 8118 43494
rect 8142 43492 8198 43494
rect 11375 43002 11431 43004
rect 11455 43002 11511 43004
rect 11535 43002 11591 43004
rect 11615 43002 11671 43004
rect 11375 42950 11421 43002
rect 11421 42950 11431 43002
rect 11455 42950 11485 43002
rect 11485 42950 11497 43002
rect 11497 42950 11511 43002
rect 11535 42950 11549 43002
rect 11549 42950 11561 43002
rect 11561 42950 11591 43002
rect 11615 42950 11625 43002
rect 11625 42950 11671 43002
rect 11375 42948 11431 42950
rect 11455 42948 11511 42950
rect 11535 42948 11591 42950
rect 11615 42948 11671 42950
rect 7902 42458 7958 42460
rect 7982 42458 8038 42460
rect 8062 42458 8118 42460
rect 8142 42458 8198 42460
rect 7902 42406 7948 42458
rect 7948 42406 7958 42458
rect 7982 42406 8012 42458
rect 8012 42406 8024 42458
rect 8024 42406 8038 42458
rect 8062 42406 8076 42458
rect 8076 42406 8088 42458
rect 8088 42406 8118 42458
rect 8142 42406 8152 42458
rect 8152 42406 8198 42458
rect 7902 42404 7958 42406
rect 7982 42404 8038 42406
rect 8062 42404 8118 42406
rect 8142 42404 8198 42406
rect 11375 41914 11431 41916
rect 11455 41914 11511 41916
rect 11535 41914 11591 41916
rect 11615 41914 11671 41916
rect 11375 41862 11421 41914
rect 11421 41862 11431 41914
rect 11455 41862 11485 41914
rect 11485 41862 11497 41914
rect 11497 41862 11511 41914
rect 11535 41862 11549 41914
rect 11549 41862 11561 41914
rect 11561 41862 11591 41914
rect 11615 41862 11625 41914
rect 11625 41862 11671 41914
rect 11375 41860 11431 41862
rect 11455 41860 11511 41862
rect 11535 41860 11591 41862
rect 11615 41860 11671 41862
rect 7902 41370 7958 41372
rect 7982 41370 8038 41372
rect 8062 41370 8118 41372
rect 8142 41370 8198 41372
rect 7902 41318 7948 41370
rect 7948 41318 7958 41370
rect 7982 41318 8012 41370
rect 8012 41318 8024 41370
rect 8024 41318 8038 41370
rect 8062 41318 8076 41370
rect 8076 41318 8088 41370
rect 8088 41318 8118 41370
rect 8142 41318 8152 41370
rect 8152 41318 8198 41370
rect 7902 41316 7958 41318
rect 7982 41316 8038 41318
rect 8062 41316 8118 41318
rect 8142 41316 8198 41318
rect 11375 40826 11431 40828
rect 11455 40826 11511 40828
rect 11535 40826 11591 40828
rect 11615 40826 11671 40828
rect 11375 40774 11421 40826
rect 11421 40774 11431 40826
rect 11455 40774 11485 40826
rect 11485 40774 11497 40826
rect 11497 40774 11511 40826
rect 11535 40774 11549 40826
rect 11549 40774 11561 40826
rect 11561 40774 11591 40826
rect 11615 40774 11625 40826
rect 11625 40774 11671 40826
rect 11375 40772 11431 40774
rect 11455 40772 11511 40774
rect 11535 40772 11591 40774
rect 11615 40772 11671 40774
rect 7902 40282 7958 40284
rect 7982 40282 8038 40284
rect 8062 40282 8118 40284
rect 8142 40282 8198 40284
rect 7902 40230 7948 40282
rect 7948 40230 7958 40282
rect 7982 40230 8012 40282
rect 8012 40230 8024 40282
rect 8024 40230 8038 40282
rect 8062 40230 8076 40282
rect 8076 40230 8088 40282
rect 8088 40230 8118 40282
rect 8142 40230 8152 40282
rect 8152 40230 8198 40282
rect 7902 40228 7958 40230
rect 7982 40228 8038 40230
rect 8062 40228 8118 40230
rect 8142 40228 8198 40230
rect 11375 39738 11431 39740
rect 11455 39738 11511 39740
rect 11535 39738 11591 39740
rect 11615 39738 11671 39740
rect 11375 39686 11421 39738
rect 11421 39686 11431 39738
rect 11455 39686 11485 39738
rect 11485 39686 11497 39738
rect 11497 39686 11511 39738
rect 11535 39686 11549 39738
rect 11549 39686 11561 39738
rect 11561 39686 11591 39738
rect 11615 39686 11625 39738
rect 11625 39686 11671 39738
rect 11375 39684 11431 39686
rect 11455 39684 11511 39686
rect 11535 39684 11591 39686
rect 11615 39684 11671 39686
rect 7902 39194 7958 39196
rect 7982 39194 8038 39196
rect 8062 39194 8118 39196
rect 8142 39194 8198 39196
rect 7902 39142 7948 39194
rect 7948 39142 7958 39194
rect 7982 39142 8012 39194
rect 8012 39142 8024 39194
rect 8024 39142 8038 39194
rect 8062 39142 8076 39194
rect 8076 39142 8088 39194
rect 8088 39142 8118 39194
rect 8142 39142 8152 39194
rect 8152 39142 8198 39194
rect 7902 39140 7958 39142
rect 7982 39140 8038 39142
rect 8062 39140 8118 39142
rect 8142 39140 8198 39142
rect 11375 38650 11431 38652
rect 11455 38650 11511 38652
rect 11535 38650 11591 38652
rect 11615 38650 11671 38652
rect 11375 38598 11421 38650
rect 11421 38598 11431 38650
rect 11455 38598 11485 38650
rect 11485 38598 11497 38650
rect 11497 38598 11511 38650
rect 11535 38598 11549 38650
rect 11549 38598 11561 38650
rect 11561 38598 11591 38650
rect 11615 38598 11625 38650
rect 11625 38598 11671 38650
rect 11375 38596 11431 38598
rect 11455 38596 11511 38598
rect 11535 38596 11591 38598
rect 11615 38596 11671 38598
rect 7902 38106 7958 38108
rect 7982 38106 8038 38108
rect 8062 38106 8118 38108
rect 8142 38106 8198 38108
rect 7902 38054 7948 38106
rect 7948 38054 7958 38106
rect 7982 38054 8012 38106
rect 8012 38054 8024 38106
rect 8024 38054 8038 38106
rect 8062 38054 8076 38106
rect 8076 38054 8088 38106
rect 8088 38054 8118 38106
rect 8142 38054 8152 38106
rect 8152 38054 8198 38106
rect 7902 38052 7958 38054
rect 7982 38052 8038 38054
rect 8062 38052 8118 38054
rect 8142 38052 8198 38054
rect 11375 37562 11431 37564
rect 11455 37562 11511 37564
rect 11535 37562 11591 37564
rect 11615 37562 11671 37564
rect 11375 37510 11421 37562
rect 11421 37510 11431 37562
rect 11455 37510 11485 37562
rect 11485 37510 11497 37562
rect 11497 37510 11511 37562
rect 11535 37510 11549 37562
rect 11549 37510 11561 37562
rect 11561 37510 11591 37562
rect 11615 37510 11625 37562
rect 11625 37510 11671 37562
rect 11375 37508 11431 37510
rect 11455 37508 11511 37510
rect 11535 37508 11591 37510
rect 11615 37508 11671 37510
rect 7902 37018 7958 37020
rect 7982 37018 8038 37020
rect 8062 37018 8118 37020
rect 8142 37018 8198 37020
rect 7902 36966 7948 37018
rect 7948 36966 7958 37018
rect 7982 36966 8012 37018
rect 8012 36966 8024 37018
rect 8024 36966 8038 37018
rect 8062 36966 8076 37018
rect 8076 36966 8088 37018
rect 8088 36966 8118 37018
rect 8142 36966 8152 37018
rect 8152 36966 8198 37018
rect 7902 36964 7958 36966
rect 7982 36964 8038 36966
rect 8062 36964 8118 36966
rect 8142 36964 8198 36966
rect 7902 35930 7958 35932
rect 7982 35930 8038 35932
rect 8062 35930 8118 35932
rect 8142 35930 8198 35932
rect 7902 35878 7948 35930
rect 7948 35878 7958 35930
rect 7982 35878 8012 35930
rect 8012 35878 8024 35930
rect 8024 35878 8038 35930
rect 8062 35878 8076 35930
rect 8076 35878 8088 35930
rect 8088 35878 8118 35930
rect 8142 35878 8152 35930
rect 8152 35878 8198 35930
rect 7902 35876 7958 35878
rect 7982 35876 8038 35878
rect 8062 35876 8118 35878
rect 8142 35876 8198 35878
rect 7902 34842 7958 34844
rect 7982 34842 8038 34844
rect 8062 34842 8118 34844
rect 8142 34842 8198 34844
rect 7902 34790 7948 34842
rect 7948 34790 7958 34842
rect 7982 34790 8012 34842
rect 8012 34790 8024 34842
rect 8024 34790 8038 34842
rect 8062 34790 8076 34842
rect 8076 34790 8088 34842
rect 8088 34790 8118 34842
rect 8142 34790 8152 34842
rect 8152 34790 8198 34842
rect 7902 34788 7958 34790
rect 7982 34788 8038 34790
rect 8062 34788 8118 34790
rect 8142 34788 8198 34790
rect 4429 34298 4485 34300
rect 4509 34298 4565 34300
rect 4589 34298 4645 34300
rect 4669 34298 4725 34300
rect 4429 34246 4475 34298
rect 4475 34246 4485 34298
rect 4509 34246 4539 34298
rect 4539 34246 4551 34298
rect 4551 34246 4565 34298
rect 4589 34246 4603 34298
rect 4603 34246 4615 34298
rect 4615 34246 4645 34298
rect 4669 34246 4679 34298
rect 4679 34246 4725 34298
rect 4429 34244 4485 34246
rect 4509 34244 4565 34246
rect 4589 34244 4645 34246
rect 4669 34244 4725 34246
rect 7902 33754 7958 33756
rect 7982 33754 8038 33756
rect 8062 33754 8118 33756
rect 8142 33754 8198 33756
rect 7902 33702 7948 33754
rect 7948 33702 7958 33754
rect 7982 33702 8012 33754
rect 8012 33702 8024 33754
rect 8024 33702 8038 33754
rect 8062 33702 8076 33754
rect 8076 33702 8088 33754
rect 8088 33702 8118 33754
rect 8142 33702 8152 33754
rect 8152 33702 8198 33754
rect 7902 33700 7958 33702
rect 7982 33700 8038 33702
rect 8062 33700 8118 33702
rect 8142 33700 8198 33702
rect 4429 33210 4485 33212
rect 4509 33210 4565 33212
rect 4589 33210 4645 33212
rect 4669 33210 4725 33212
rect 4429 33158 4475 33210
rect 4475 33158 4485 33210
rect 4509 33158 4539 33210
rect 4539 33158 4551 33210
rect 4551 33158 4565 33210
rect 4589 33158 4603 33210
rect 4603 33158 4615 33210
rect 4615 33158 4645 33210
rect 4669 33158 4679 33210
rect 4679 33158 4725 33210
rect 4429 33156 4485 33158
rect 4509 33156 4565 33158
rect 4589 33156 4645 33158
rect 4669 33156 4725 33158
rect 7902 32666 7958 32668
rect 7982 32666 8038 32668
rect 8062 32666 8118 32668
rect 8142 32666 8198 32668
rect 7902 32614 7948 32666
rect 7948 32614 7958 32666
rect 7982 32614 8012 32666
rect 8012 32614 8024 32666
rect 8024 32614 8038 32666
rect 8062 32614 8076 32666
rect 8076 32614 8088 32666
rect 8088 32614 8118 32666
rect 8142 32614 8152 32666
rect 8152 32614 8198 32666
rect 7902 32612 7958 32614
rect 7982 32612 8038 32614
rect 8062 32612 8118 32614
rect 8142 32612 8198 32614
rect 4429 32122 4485 32124
rect 4509 32122 4565 32124
rect 4589 32122 4645 32124
rect 4669 32122 4725 32124
rect 4429 32070 4475 32122
rect 4475 32070 4485 32122
rect 4509 32070 4539 32122
rect 4539 32070 4551 32122
rect 4551 32070 4565 32122
rect 4589 32070 4603 32122
rect 4603 32070 4615 32122
rect 4615 32070 4645 32122
rect 4669 32070 4679 32122
rect 4679 32070 4725 32122
rect 4429 32068 4485 32070
rect 4509 32068 4565 32070
rect 4589 32068 4645 32070
rect 4669 32068 4725 32070
rect 7902 31578 7958 31580
rect 7982 31578 8038 31580
rect 8062 31578 8118 31580
rect 8142 31578 8198 31580
rect 7902 31526 7948 31578
rect 7948 31526 7958 31578
rect 7982 31526 8012 31578
rect 8012 31526 8024 31578
rect 8024 31526 8038 31578
rect 8062 31526 8076 31578
rect 8076 31526 8088 31578
rect 8088 31526 8118 31578
rect 8142 31526 8152 31578
rect 8152 31526 8198 31578
rect 7902 31524 7958 31526
rect 7982 31524 8038 31526
rect 8062 31524 8118 31526
rect 8142 31524 8198 31526
rect 4429 31034 4485 31036
rect 4509 31034 4565 31036
rect 4589 31034 4645 31036
rect 4669 31034 4725 31036
rect 4429 30982 4475 31034
rect 4475 30982 4485 31034
rect 4509 30982 4539 31034
rect 4539 30982 4551 31034
rect 4551 30982 4565 31034
rect 4589 30982 4603 31034
rect 4603 30982 4615 31034
rect 4615 30982 4645 31034
rect 4669 30982 4679 31034
rect 4679 30982 4725 31034
rect 4429 30980 4485 30982
rect 4509 30980 4565 30982
rect 4589 30980 4645 30982
rect 4669 30980 4725 30982
rect 7902 30490 7958 30492
rect 7982 30490 8038 30492
rect 8062 30490 8118 30492
rect 8142 30490 8198 30492
rect 7902 30438 7948 30490
rect 7948 30438 7958 30490
rect 7982 30438 8012 30490
rect 8012 30438 8024 30490
rect 8024 30438 8038 30490
rect 8062 30438 8076 30490
rect 8076 30438 8088 30490
rect 8088 30438 8118 30490
rect 8142 30438 8152 30490
rect 8152 30438 8198 30490
rect 7902 30436 7958 30438
rect 7982 30436 8038 30438
rect 8062 30436 8118 30438
rect 8142 30436 8198 30438
rect 4429 29946 4485 29948
rect 4509 29946 4565 29948
rect 4589 29946 4645 29948
rect 4669 29946 4725 29948
rect 4429 29894 4475 29946
rect 4475 29894 4485 29946
rect 4509 29894 4539 29946
rect 4539 29894 4551 29946
rect 4551 29894 4565 29946
rect 4589 29894 4603 29946
rect 4603 29894 4615 29946
rect 4615 29894 4645 29946
rect 4669 29894 4679 29946
rect 4679 29894 4725 29946
rect 4429 29892 4485 29894
rect 4509 29892 4565 29894
rect 4589 29892 4645 29894
rect 4669 29892 4725 29894
rect 7902 29402 7958 29404
rect 7982 29402 8038 29404
rect 8062 29402 8118 29404
rect 8142 29402 8198 29404
rect 7902 29350 7948 29402
rect 7948 29350 7958 29402
rect 7982 29350 8012 29402
rect 8012 29350 8024 29402
rect 8024 29350 8038 29402
rect 8062 29350 8076 29402
rect 8076 29350 8088 29402
rect 8088 29350 8118 29402
rect 8142 29350 8152 29402
rect 8152 29350 8198 29402
rect 7902 29348 7958 29350
rect 7982 29348 8038 29350
rect 8062 29348 8118 29350
rect 8142 29348 8198 29350
rect 4429 28858 4485 28860
rect 4509 28858 4565 28860
rect 4589 28858 4645 28860
rect 4669 28858 4725 28860
rect 4429 28806 4475 28858
rect 4475 28806 4485 28858
rect 4509 28806 4539 28858
rect 4539 28806 4551 28858
rect 4551 28806 4565 28858
rect 4589 28806 4603 28858
rect 4603 28806 4615 28858
rect 4615 28806 4645 28858
rect 4669 28806 4679 28858
rect 4679 28806 4725 28858
rect 4429 28804 4485 28806
rect 4509 28804 4565 28806
rect 4589 28804 4645 28806
rect 4669 28804 4725 28806
rect 7902 28314 7958 28316
rect 7982 28314 8038 28316
rect 8062 28314 8118 28316
rect 8142 28314 8198 28316
rect 7902 28262 7948 28314
rect 7948 28262 7958 28314
rect 7982 28262 8012 28314
rect 8012 28262 8024 28314
rect 8024 28262 8038 28314
rect 8062 28262 8076 28314
rect 8076 28262 8088 28314
rect 8088 28262 8118 28314
rect 8142 28262 8152 28314
rect 8152 28262 8198 28314
rect 7902 28260 7958 28262
rect 7982 28260 8038 28262
rect 8062 28260 8118 28262
rect 8142 28260 8198 28262
rect 4429 27770 4485 27772
rect 4509 27770 4565 27772
rect 4589 27770 4645 27772
rect 4669 27770 4725 27772
rect 4429 27718 4475 27770
rect 4475 27718 4485 27770
rect 4509 27718 4539 27770
rect 4539 27718 4551 27770
rect 4551 27718 4565 27770
rect 4589 27718 4603 27770
rect 4603 27718 4615 27770
rect 4615 27718 4645 27770
rect 4669 27718 4679 27770
rect 4679 27718 4725 27770
rect 4429 27716 4485 27718
rect 4509 27716 4565 27718
rect 4589 27716 4645 27718
rect 4669 27716 4725 27718
rect 7902 27226 7958 27228
rect 7982 27226 8038 27228
rect 8062 27226 8118 27228
rect 8142 27226 8198 27228
rect 7902 27174 7948 27226
rect 7948 27174 7958 27226
rect 7982 27174 8012 27226
rect 8012 27174 8024 27226
rect 8024 27174 8038 27226
rect 8062 27174 8076 27226
rect 8076 27174 8088 27226
rect 8088 27174 8118 27226
rect 8142 27174 8152 27226
rect 8152 27174 8198 27226
rect 7902 27172 7958 27174
rect 7982 27172 8038 27174
rect 8062 27172 8118 27174
rect 8142 27172 8198 27174
rect 4429 26682 4485 26684
rect 4509 26682 4565 26684
rect 4589 26682 4645 26684
rect 4669 26682 4725 26684
rect 4429 26630 4475 26682
rect 4475 26630 4485 26682
rect 4509 26630 4539 26682
rect 4539 26630 4551 26682
rect 4551 26630 4565 26682
rect 4589 26630 4603 26682
rect 4603 26630 4615 26682
rect 4615 26630 4645 26682
rect 4669 26630 4679 26682
rect 4679 26630 4725 26682
rect 4429 26628 4485 26630
rect 4509 26628 4565 26630
rect 4589 26628 4645 26630
rect 4669 26628 4725 26630
rect 7902 26138 7958 26140
rect 7982 26138 8038 26140
rect 8062 26138 8118 26140
rect 8142 26138 8198 26140
rect 7902 26086 7948 26138
rect 7948 26086 7958 26138
rect 7982 26086 8012 26138
rect 8012 26086 8024 26138
rect 8024 26086 8038 26138
rect 8062 26086 8076 26138
rect 8076 26086 8088 26138
rect 8088 26086 8118 26138
rect 8142 26086 8152 26138
rect 8152 26086 8198 26138
rect 7902 26084 7958 26086
rect 7982 26084 8038 26086
rect 8062 26084 8118 26086
rect 8142 26084 8198 26086
rect 4429 25594 4485 25596
rect 4509 25594 4565 25596
rect 4589 25594 4645 25596
rect 4669 25594 4725 25596
rect 4429 25542 4475 25594
rect 4475 25542 4485 25594
rect 4509 25542 4539 25594
rect 4539 25542 4551 25594
rect 4551 25542 4565 25594
rect 4589 25542 4603 25594
rect 4603 25542 4615 25594
rect 4615 25542 4645 25594
rect 4669 25542 4679 25594
rect 4679 25542 4725 25594
rect 4429 25540 4485 25542
rect 4509 25540 4565 25542
rect 4589 25540 4645 25542
rect 4669 25540 4725 25542
rect 7902 25050 7958 25052
rect 7982 25050 8038 25052
rect 8062 25050 8118 25052
rect 8142 25050 8198 25052
rect 7902 24998 7948 25050
rect 7948 24998 7958 25050
rect 7982 24998 8012 25050
rect 8012 24998 8024 25050
rect 8024 24998 8038 25050
rect 8062 24998 8076 25050
rect 8076 24998 8088 25050
rect 8088 24998 8118 25050
rect 8142 24998 8152 25050
rect 8152 24998 8198 25050
rect 7902 24996 7958 24998
rect 7982 24996 8038 24998
rect 8062 24996 8118 24998
rect 8142 24996 8198 24998
rect 4429 24506 4485 24508
rect 4509 24506 4565 24508
rect 4589 24506 4645 24508
rect 4669 24506 4725 24508
rect 4429 24454 4475 24506
rect 4475 24454 4485 24506
rect 4509 24454 4539 24506
rect 4539 24454 4551 24506
rect 4551 24454 4565 24506
rect 4589 24454 4603 24506
rect 4603 24454 4615 24506
rect 4615 24454 4645 24506
rect 4669 24454 4679 24506
rect 4679 24454 4725 24506
rect 4429 24452 4485 24454
rect 4509 24452 4565 24454
rect 4589 24452 4645 24454
rect 4669 24452 4725 24454
rect 7902 23962 7958 23964
rect 7982 23962 8038 23964
rect 8062 23962 8118 23964
rect 8142 23962 8198 23964
rect 7902 23910 7948 23962
rect 7948 23910 7958 23962
rect 7982 23910 8012 23962
rect 8012 23910 8024 23962
rect 8024 23910 8038 23962
rect 8062 23910 8076 23962
rect 8076 23910 8088 23962
rect 8088 23910 8118 23962
rect 8142 23910 8152 23962
rect 8152 23910 8198 23962
rect 7902 23908 7958 23910
rect 7982 23908 8038 23910
rect 8062 23908 8118 23910
rect 8142 23908 8198 23910
rect 4429 23418 4485 23420
rect 4509 23418 4565 23420
rect 4589 23418 4645 23420
rect 4669 23418 4725 23420
rect 4429 23366 4475 23418
rect 4475 23366 4485 23418
rect 4509 23366 4539 23418
rect 4539 23366 4551 23418
rect 4551 23366 4565 23418
rect 4589 23366 4603 23418
rect 4603 23366 4615 23418
rect 4615 23366 4645 23418
rect 4669 23366 4679 23418
rect 4679 23366 4725 23418
rect 4429 23364 4485 23366
rect 4509 23364 4565 23366
rect 4589 23364 4645 23366
rect 4669 23364 4725 23366
rect 7902 22874 7958 22876
rect 7982 22874 8038 22876
rect 8062 22874 8118 22876
rect 8142 22874 8198 22876
rect 7902 22822 7948 22874
rect 7948 22822 7958 22874
rect 7982 22822 8012 22874
rect 8012 22822 8024 22874
rect 8024 22822 8038 22874
rect 8062 22822 8076 22874
rect 8076 22822 8088 22874
rect 8088 22822 8118 22874
rect 8142 22822 8152 22874
rect 8152 22822 8198 22874
rect 7902 22820 7958 22822
rect 7982 22820 8038 22822
rect 8062 22820 8118 22822
rect 8142 22820 8198 22822
rect 4429 22330 4485 22332
rect 4509 22330 4565 22332
rect 4589 22330 4645 22332
rect 4669 22330 4725 22332
rect 4429 22278 4475 22330
rect 4475 22278 4485 22330
rect 4509 22278 4539 22330
rect 4539 22278 4551 22330
rect 4551 22278 4565 22330
rect 4589 22278 4603 22330
rect 4603 22278 4615 22330
rect 4615 22278 4645 22330
rect 4669 22278 4679 22330
rect 4679 22278 4725 22330
rect 4429 22276 4485 22278
rect 4509 22276 4565 22278
rect 4589 22276 4645 22278
rect 4669 22276 4725 22278
rect 7902 21786 7958 21788
rect 7982 21786 8038 21788
rect 8062 21786 8118 21788
rect 8142 21786 8198 21788
rect 7902 21734 7948 21786
rect 7948 21734 7958 21786
rect 7982 21734 8012 21786
rect 8012 21734 8024 21786
rect 8024 21734 8038 21786
rect 8062 21734 8076 21786
rect 8076 21734 8088 21786
rect 8088 21734 8118 21786
rect 8142 21734 8152 21786
rect 8152 21734 8198 21786
rect 7902 21732 7958 21734
rect 7982 21732 8038 21734
rect 8062 21732 8118 21734
rect 8142 21732 8198 21734
rect 4429 21242 4485 21244
rect 4509 21242 4565 21244
rect 4589 21242 4645 21244
rect 4669 21242 4725 21244
rect 4429 21190 4475 21242
rect 4475 21190 4485 21242
rect 4509 21190 4539 21242
rect 4539 21190 4551 21242
rect 4551 21190 4565 21242
rect 4589 21190 4603 21242
rect 4603 21190 4615 21242
rect 4615 21190 4645 21242
rect 4669 21190 4679 21242
rect 4679 21190 4725 21242
rect 4429 21188 4485 21190
rect 4509 21188 4565 21190
rect 4589 21188 4645 21190
rect 4669 21188 4725 21190
rect 7902 20698 7958 20700
rect 7982 20698 8038 20700
rect 8062 20698 8118 20700
rect 8142 20698 8198 20700
rect 7902 20646 7948 20698
rect 7948 20646 7958 20698
rect 7982 20646 8012 20698
rect 8012 20646 8024 20698
rect 8024 20646 8038 20698
rect 8062 20646 8076 20698
rect 8076 20646 8088 20698
rect 8088 20646 8118 20698
rect 8142 20646 8152 20698
rect 8152 20646 8198 20698
rect 7902 20644 7958 20646
rect 7982 20644 8038 20646
rect 8062 20644 8118 20646
rect 8142 20644 8198 20646
rect 4429 20154 4485 20156
rect 4509 20154 4565 20156
rect 4589 20154 4645 20156
rect 4669 20154 4725 20156
rect 4429 20102 4475 20154
rect 4475 20102 4485 20154
rect 4509 20102 4539 20154
rect 4539 20102 4551 20154
rect 4551 20102 4565 20154
rect 4589 20102 4603 20154
rect 4603 20102 4615 20154
rect 4615 20102 4645 20154
rect 4669 20102 4679 20154
rect 4679 20102 4725 20154
rect 4429 20100 4485 20102
rect 4509 20100 4565 20102
rect 4589 20100 4645 20102
rect 4669 20100 4725 20102
rect 7902 19610 7958 19612
rect 7982 19610 8038 19612
rect 8062 19610 8118 19612
rect 8142 19610 8198 19612
rect 7902 19558 7948 19610
rect 7948 19558 7958 19610
rect 7982 19558 8012 19610
rect 8012 19558 8024 19610
rect 8024 19558 8038 19610
rect 8062 19558 8076 19610
rect 8076 19558 8088 19610
rect 8088 19558 8118 19610
rect 8142 19558 8152 19610
rect 8152 19558 8198 19610
rect 7902 19556 7958 19558
rect 7982 19556 8038 19558
rect 8062 19556 8118 19558
rect 8142 19556 8198 19558
rect 4429 19066 4485 19068
rect 4509 19066 4565 19068
rect 4589 19066 4645 19068
rect 4669 19066 4725 19068
rect 4429 19014 4475 19066
rect 4475 19014 4485 19066
rect 4509 19014 4539 19066
rect 4539 19014 4551 19066
rect 4551 19014 4565 19066
rect 4589 19014 4603 19066
rect 4603 19014 4615 19066
rect 4615 19014 4645 19066
rect 4669 19014 4679 19066
rect 4679 19014 4725 19066
rect 4429 19012 4485 19014
rect 4509 19012 4565 19014
rect 4589 19012 4645 19014
rect 4669 19012 4725 19014
rect 7902 18522 7958 18524
rect 7982 18522 8038 18524
rect 8062 18522 8118 18524
rect 8142 18522 8198 18524
rect 7902 18470 7948 18522
rect 7948 18470 7958 18522
rect 7982 18470 8012 18522
rect 8012 18470 8024 18522
rect 8024 18470 8038 18522
rect 8062 18470 8076 18522
rect 8076 18470 8088 18522
rect 8088 18470 8118 18522
rect 8142 18470 8152 18522
rect 8152 18470 8198 18522
rect 7902 18468 7958 18470
rect 7982 18468 8038 18470
rect 8062 18468 8118 18470
rect 8142 18468 8198 18470
rect 4429 17978 4485 17980
rect 4509 17978 4565 17980
rect 4589 17978 4645 17980
rect 4669 17978 4725 17980
rect 4429 17926 4475 17978
rect 4475 17926 4485 17978
rect 4509 17926 4539 17978
rect 4539 17926 4551 17978
rect 4551 17926 4565 17978
rect 4589 17926 4603 17978
rect 4603 17926 4615 17978
rect 4615 17926 4645 17978
rect 4669 17926 4679 17978
rect 4679 17926 4725 17978
rect 4429 17924 4485 17926
rect 4509 17924 4565 17926
rect 4589 17924 4645 17926
rect 4669 17924 4725 17926
rect 4429 16890 4485 16892
rect 4509 16890 4565 16892
rect 4589 16890 4645 16892
rect 4669 16890 4725 16892
rect 4429 16838 4475 16890
rect 4475 16838 4485 16890
rect 4509 16838 4539 16890
rect 4539 16838 4551 16890
rect 4551 16838 4565 16890
rect 4589 16838 4603 16890
rect 4603 16838 4615 16890
rect 4615 16838 4645 16890
rect 4669 16838 4679 16890
rect 4679 16838 4725 16890
rect 4429 16836 4485 16838
rect 4509 16836 4565 16838
rect 4589 16836 4645 16838
rect 4669 16836 4725 16838
rect 4429 15802 4485 15804
rect 4509 15802 4565 15804
rect 4589 15802 4645 15804
rect 4669 15802 4725 15804
rect 4429 15750 4475 15802
rect 4475 15750 4485 15802
rect 4509 15750 4539 15802
rect 4539 15750 4551 15802
rect 4551 15750 4565 15802
rect 4589 15750 4603 15802
rect 4603 15750 4615 15802
rect 4615 15750 4645 15802
rect 4669 15750 4679 15802
rect 4679 15750 4725 15802
rect 4429 15748 4485 15750
rect 4509 15748 4565 15750
rect 4589 15748 4645 15750
rect 4669 15748 4725 15750
rect 4429 14714 4485 14716
rect 4509 14714 4565 14716
rect 4589 14714 4645 14716
rect 4669 14714 4725 14716
rect 4429 14662 4475 14714
rect 4475 14662 4485 14714
rect 4509 14662 4539 14714
rect 4539 14662 4551 14714
rect 4551 14662 4565 14714
rect 4589 14662 4603 14714
rect 4603 14662 4615 14714
rect 4615 14662 4645 14714
rect 4669 14662 4679 14714
rect 4679 14662 4725 14714
rect 4429 14660 4485 14662
rect 4509 14660 4565 14662
rect 4589 14660 4645 14662
rect 4669 14660 4725 14662
rect 4429 13626 4485 13628
rect 4509 13626 4565 13628
rect 4589 13626 4645 13628
rect 4669 13626 4725 13628
rect 4429 13574 4475 13626
rect 4475 13574 4485 13626
rect 4509 13574 4539 13626
rect 4539 13574 4551 13626
rect 4551 13574 4565 13626
rect 4589 13574 4603 13626
rect 4603 13574 4615 13626
rect 4615 13574 4645 13626
rect 4669 13574 4679 13626
rect 4679 13574 4725 13626
rect 4429 13572 4485 13574
rect 4509 13572 4565 13574
rect 4589 13572 4645 13574
rect 4669 13572 4725 13574
rect 4429 12538 4485 12540
rect 4509 12538 4565 12540
rect 4589 12538 4645 12540
rect 4669 12538 4725 12540
rect 4429 12486 4475 12538
rect 4475 12486 4485 12538
rect 4509 12486 4539 12538
rect 4539 12486 4551 12538
rect 4551 12486 4565 12538
rect 4589 12486 4603 12538
rect 4603 12486 4615 12538
rect 4615 12486 4645 12538
rect 4669 12486 4679 12538
rect 4679 12486 4725 12538
rect 4429 12484 4485 12486
rect 4509 12484 4565 12486
rect 4589 12484 4645 12486
rect 4669 12484 4725 12486
rect 4429 11450 4485 11452
rect 4509 11450 4565 11452
rect 4589 11450 4645 11452
rect 4669 11450 4725 11452
rect 4429 11398 4475 11450
rect 4475 11398 4485 11450
rect 4509 11398 4539 11450
rect 4539 11398 4551 11450
rect 4551 11398 4565 11450
rect 4589 11398 4603 11450
rect 4603 11398 4615 11450
rect 4615 11398 4645 11450
rect 4669 11398 4679 11450
rect 4679 11398 4725 11450
rect 4429 11396 4485 11398
rect 4509 11396 4565 11398
rect 4589 11396 4645 11398
rect 4669 11396 4725 11398
rect 4429 10362 4485 10364
rect 4509 10362 4565 10364
rect 4589 10362 4645 10364
rect 4669 10362 4725 10364
rect 4429 10310 4475 10362
rect 4475 10310 4485 10362
rect 4509 10310 4539 10362
rect 4539 10310 4551 10362
rect 4551 10310 4565 10362
rect 4589 10310 4603 10362
rect 4603 10310 4615 10362
rect 4615 10310 4645 10362
rect 4669 10310 4679 10362
rect 4679 10310 4725 10362
rect 4429 10308 4485 10310
rect 4509 10308 4565 10310
rect 4589 10308 4645 10310
rect 4669 10308 4725 10310
rect 4429 9274 4485 9276
rect 4509 9274 4565 9276
rect 4589 9274 4645 9276
rect 4669 9274 4725 9276
rect 4429 9222 4475 9274
rect 4475 9222 4485 9274
rect 4509 9222 4539 9274
rect 4539 9222 4551 9274
rect 4551 9222 4565 9274
rect 4589 9222 4603 9274
rect 4603 9222 4615 9274
rect 4615 9222 4645 9274
rect 4669 9222 4679 9274
rect 4679 9222 4725 9274
rect 4429 9220 4485 9222
rect 4509 9220 4565 9222
rect 4589 9220 4645 9222
rect 4669 9220 4725 9222
rect 4429 8186 4485 8188
rect 4509 8186 4565 8188
rect 4589 8186 4645 8188
rect 4669 8186 4725 8188
rect 4429 8134 4475 8186
rect 4475 8134 4485 8186
rect 4509 8134 4539 8186
rect 4539 8134 4551 8186
rect 4551 8134 4565 8186
rect 4589 8134 4603 8186
rect 4603 8134 4615 8186
rect 4615 8134 4645 8186
rect 4669 8134 4679 8186
rect 4679 8134 4725 8186
rect 4429 8132 4485 8134
rect 4509 8132 4565 8134
rect 4589 8132 4645 8134
rect 4669 8132 4725 8134
rect 4429 7098 4485 7100
rect 4509 7098 4565 7100
rect 4589 7098 4645 7100
rect 4669 7098 4725 7100
rect 4429 7046 4475 7098
rect 4475 7046 4485 7098
rect 4509 7046 4539 7098
rect 4539 7046 4551 7098
rect 4551 7046 4565 7098
rect 4589 7046 4603 7098
rect 4603 7046 4615 7098
rect 4615 7046 4645 7098
rect 4669 7046 4679 7098
rect 4679 7046 4725 7098
rect 4429 7044 4485 7046
rect 4509 7044 4565 7046
rect 4589 7044 4645 7046
rect 4669 7044 4725 7046
rect 4066 6160 4122 6216
rect 3330 1400 3386 1456
rect 4066 2080 4122 2136
rect 4429 6010 4485 6012
rect 4509 6010 4565 6012
rect 4589 6010 4645 6012
rect 4669 6010 4725 6012
rect 4429 5958 4475 6010
rect 4475 5958 4485 6010
rect 4509 5958 4539 6010
rect 4539 5958 4551 6010
rect 4551 5958 4565 6010
rect 4589 5958 4603 6010
rect 4603 5958 4615 6010
rect 4615 5958 4645 6010
rect 4669 5958 4679 6010
rect 4679 5958 4725 6010
rect 4429 5956 4485 5958
rect 4509 5956 4565 5958
rect 4589 5956 4645 5958
rect 4669 5956 4725 5958
rect 4429 4922 4485 4924
rect 4509 4922 4565 4924
rect 4589 4922 4645 4924
rect 4669 4922 4725 4924
rect 4429 4870 4475 4922
rect 4475 4870 4485 4922
rect 4509 4870 4539 4922
rect 4539 4870 4551 4922
rect 4551 4870 4565 4922
rect 4589 4870 4603 4922
rect 4603 4870 4615 4922
rect 4615 4870 4645 4922
rect 4669 4870 4679 4922
rect 4679 4870 4725 4922
rect 4429 4868 4485 4870
rect 4509 4868 4565 4870
rect 4589 4868 4645 4870
rect 4669 4868 4725 4870
rect 4429 3834 4485 3836
rect 4509 3834 4565 3836
rect 4589 3834 4645 3836
rect 4669 3834 4725 3836
rect 4429 3782 4475 3834
rect 4475 3782 4485 3834
rect 4509 3782 4539 3834
rect 4539 3782 4551 3834
rect 4551 3782 4565 3834
rect 4589 3782 4603 3834
rect 4603 3782 4615 3834
rect 4615 3782 4645 3834
rect 4669 3782 4679 3834
rect 4679 3782 4725 3834
rect 4429 3780 4485 3782
rect 4509 3780 4565 3782
rect 4589 3780 4645 3782
rect 4669 3780 4725 3782
rect 7902 17434 7958 17436
rect 7982 17434 8038 17436
rect 8062 17434 8118 17436
rect 8142 17434 8198 17436
rect 7902 17382 7948 17434
rect 7948 17382 7958 17434
rect 7982 17382 8012 17434
rect 8012 17382 8024 17434
rect 8024 17382 8038 17434
rect 8062 17382 8076 17434
rect 8076 17382 8088 17434
rect 8088 17382 8118 17434
rect 8142 17382 8152 17434
rect 8152 17382 8198 17434
rect 7902 17380 7958 17382
rect 7982 17380 8038 17382
rect 8062 17380 8118 17382
rect 8142 17380 8198 17382
rect 7902 16346 7958 16348
rect 7982 16346 8038 16348
rect 8062 16346 8118 16348
rect 8142 16346 8198 16348
rect 7902 16294 7948 16346
rect 7948 16294 7958 16346
rect 7982 16294 8012 16346
rect 8012 16294 8024 16346
rect 8024 16294 8038 16346
rect 8062 16294 8076 16346
rect 8076 16294 8088 16346
rect 8088 16294 8118 16346
rect 8142 16294 8152 16346
rect 8152 16294 8198 16346
rect 7902 16292 7958 16294
rect 7982 16292 8038 16294
rect 8062 16292 8118 16294
rect 8142 16292 8198 16294
rect 7902 15258 7958 15260
rect 7982 15258 8038 15260
rect 8062 15258 8118 15260
rect 8142 15258 8198 15260
rect 7902 15206 7948 15258
rect 7948 15206 7958 15258
rect 7982 15206 8012 15258
rect 8012 15206 8024 15258
rect 8024 15206 8038 15258
rect 8062 15206 8076 15258
rect 8076 15206 8088 15258
rect 8088 15206 8118 15258
rect 8142 15206 8152 15258
rect 8152 15206 8198 15258
rect 7902 15204 7958 15206
rect 7982 15204 8038 15206
rect 8062 15204 8118 15206
rect 8142 15204 8198 15206
rect 7902 14170 7958 14172
rect 7982 14170 8038 14172
rect 8062 14170 8118 14172
rect 8142 14170 8198 14172
rect 7902 14118 7948 14170
rect 7948 14118 7958 14170
rect 7982 14118 8012 14170
rect 8012 14118 8024 14170
rect 8024 14118 8038 14170
rect 8062 14118 8076 14170
rect 8076 14118 8088 14170
rect 8088 14118 8118 14170
rect 8142 14118 8152 14170
rect 8152 14118 8198 14170
rect 7902 14116 7958 14118
rect 7982 14116 8038 14118
rect 8062 14116 8118 14118
rect 8142 14116 8198 14118
rect 7902 13082 7958 13084
rect 7982 13082 8038 13084
rect 8062 13082 8118 13084
rect 8142 13082 8198 13084
rect 7902 13030 7948 13082
rect 7948 13030 7958 13082
rect 7982 13030 8012 13082
rect 8012 13030 8024 13082
rect 8024 13030 8038 13082
rect 8062 13030 8076 13082
rect 8076 13030 8088 13082
rect 8088 13030 8118 13082
rect 8142 13030 8152 13082
rect 8152 13030 8198 13082
rect 7902 13028 7958 13030
rect 7982 13028 8038 13030
rect 8062 13028 8118 13030
rect 8142 13028 8198 13030
rect 7902 11994 7958 11996
rect 7982 11994 8038 11996
rect 8062 11994 8118 11996
rect 8142 11994 8198 11996
rect 7902 11942 7948 11994
rect 7948 11942 7958 11994
rect 7982 11942 8012 11994
rect 8012 11942 8024 11994
rect 8024 11942 8038 11994
rect 8062 11942 8076 11994
rect 8076 11942 8088 11994
rect 8088 11942 8118 11994
rect 8142 11942 8152 11994
rect 8152 11942 8198 11994
rect 7902 11940 7958 11942
rect 7982 11940 8038 11942
rect 8062 11940 8118 11942
rect 8142 11940 8198 11942
rect 7902 10906 7958 10908
rect 7982 10906 8038 10908
rect 8062 10906 8118 10908
rect 8142 10906 8198 10908
rect 7902 10854 7948 10906
rect 7948 10854 7958 10906
rect 7982 10854 8012 10906
rect 8012 10854 8024 10906
rect 8024 10854 8038 10906
rect 8062 10854 8076 10906
rect 8076 10854 8088 10906
rect 8088 10854 8118 10906
rect 8142 10854 8152 10906
rect 8152 10854 8198 10906
rect 7902 10852 7958 10854
rect 7982 10852 8038 10854
rect 8062 10852 8118 10854
rect 8142 10852 8198 10854
rect 7902 9818 7958 9820
rect 7982 9818 8038 9820
rect 8062 9818 8118 9820
rect 8142 9818 8198 9820
rect 7902 9766 7948 9818
rect 7948 9766 7958 9818
rect 7982 9766 8012 9818
rect 8012 9766 8024 9818
rect 8024 9766 8038 9818
rect 8062 9766 8076 9818
rect 8076 9766 8088 9818
rect 8088 9766 8118 9818
rect 8142 9766 8152 9818
rect 8152 9766 8198 9818
rect 7902 9764 7958 9766
rect 7982 9764 8038 9766
rect 8062 9764 8118 9766
rect 8142 9764 8198 9766
rect 7902 8730 7958 8732
rect 7982 8730 8038 8732
rect 8062 8730 8118 8732
rect 8142 8730 8198 8732
rect 7902 8678 7948 8730
rect 7948 8678 7958 8730
rect 7982 8678 8012 8730
rect 8012 8678 8024 8730
rect 8024 8678 8038 8730
rect 8062 8678 8076 8730
rect 8076 8678 8088 8730
rect 8088 8678 8118 8730
rect 8142 8678 8152 8730
rect 8152 8678 8198 8730
rect 7902 8676 7958 8678
rect 7982 8676 8038 8678
rect 8062 8676 8118 8678
rect 8142 8676 8198 8678
rect 7902 7642 7958 7644
rect 7982 7642 8038 7644
rect 8062 7642 8118 7644
rect 8142 7642 8198 7644
rect 7902 7590 7948 7642
rect 7948 7590 7958 7642
rect 7982 7590 8012 7642
rect 8012 7590 8024 7642
rect 8024 7590 8038 7642
rect 8062 7590 8076 7642
rect 8076 7590 8088 7642
rect 8088 7590 8118 7642
rect 8142 7590 8152 7642
rect 8152 7590 8198 7642
rect 7902 7588 7958 7590
rect 7982 7588 8038 7590
rect 8062 7588 8118 7590
rect 8142 7588 8198 7590
rect 7902 6554 7958 6556
rect 7982 6554 8038 6556
rect 8062 6554 8118 6556
rect 8142 6554 8198 6556
rect 7902 6502 7948 6554
rect 7948 6502 7958 6554
rect 7982 6502 8012 6554
rect 8012 6502 8024 6554
rect 8024 6502 8038 6554
rect 8062 6502 8076 6554
rect 8076 6502 8088 6554
rect 8088 6502 8118 6554
rect 8142 6502 8152 6554
rect 8152 6502 8198 6554
rect 7902 6500 7958 6502
rect 7982 6500 8038 6502
rect 8062 6500 8118 6502
rect 8142 6500 8198 6502
rect 7902 5466 7958 5468
rect 7982 5466 8038 5468
rect 8062 5466 8118 5468
rect 8142 5466 8198 5468
rect 7902 5414 7948 5466
rect 7948 5414 7958 5466
rect 7982 5414 8012 5466
rect 8012 5414 8024 5466
rect 8024 5414 8038 5466
rect 8062 5414 8076 5466
rect 8076 5414 8088 5466
rect 8088 5414 8118 5466
rect 8142 5414 8152 5466
rect 8152 5414 8198 5466
rect 7902 5412 7958 5414
rect 7982 5412 8038 5414
rect 8062 5412 8118 5414
rect 8142 5412 8198 5414
rect 4429 2746 4485 2748
rect 4509 2746 4565 2748
rect 4589 2746 4645 2748
rect 4669 2746 4725 2748
rect 4429 2694 4475 2746
rect 4475 2694 4485 2746
rect 4509 2694 4539 2746
rect 4539 2694 4551 2746
rect 4551 2694 4565 2746
rect 4589 2694 4603 2746
rect 4603 2694 4615 2746
rect 4615 2694 4645 2746
rect 4669 2694 4679 2746
rect 4679 2694 4725 2746
rect 4429 2692 4485 2694
rect 4509 2692 4565 2694
rect 4589 2692 4645 2694
rect 4669 2692 4725 2694
rect 7902 4378 7958 4380
rect 7982 4378 8038 4380
rect 8062 4378 8118 4380
rect 8142 4378 8198 4380
rect 7902 4326 7948 4378
rect 7948 4326 7958 4378
rect 7982 4326 8012 4378
rect 8012 4326 8024 4378
rect 8024 4326 8038 4378
rect 8062 4326 8076 4378
rect 8076 4326 8088 4378
rect 8088 4326 8118 4378
rect 8142 4326 8152 4378
rect 8152 4326 8198 4378
rect 7902 4324 7958 4326
rect 7982 4324 8038 4326
rect 8062 4324 8118 4326
rect 8142 4324 8198 4326
rect 7902 3290 7958 3292
rect 7982 3290 8038 3292
rect 8062 3290 8118 3292
rect 8142 3290 8198 3292
rect 7902 3238 7948 3290
rect 7948 3238 7958 3290
rect 7982 3238 8012 3290
rect 8012 3238 8024 3290
rect 8024 3238 8038 3290
rect 8062 3238 8076 3290
rect 8076 3238 8088 3290
rect 8088 3238 8118 3290
rect 8142 3238 8152 3290
rect 8152 3238 8198 3290
rect 7902 3236 7958 3238
rect 7982 3236 8038 3238
rect 8062 3236 8118 3238
rect 8142 3236 8198 3238
rect 7902 2202 7958 2204
rect 7982 2202 8038 2204
rect 8062 2202 8118 2204
rect 8142 2202 8198 2204
rect 7902 2150 7948 2202
rect 7948 2150 7958 2202
rect 7982 2150 8012 2202
rect 8012 2150 8024 2202
rect 8024 2150 8038 2202
rect 8062 2150 8076 2202
rect 8076 2150 8088 2202
rect 8088 2150 8118 2202
rect 8142 2150 8152 2202
rect 8152 2150 8198 2202
rect 7902 2148 7958 2150
rect 7982 2148 8038 2150
rect 8062 2148 8118 2150
rect 8142 2148 8198 2150
rect 11375 36474 11431 36476
rect 11455 36474 11511 36476
rect 11535 36474 11591 36476
rect 11615 36474 11671 36476
rect 11375 36422 11421 36474
rect 11421 36422 11431 36474
rect 11455 36422 11485 36474
rect 11485 36422 11497 36474
rect 11497 36422 11511 36474
rect 11535 36422 11549 36474
rect 11549 36422 11561 36474
rect 11561 36422 11591 36474
rect 11615 36422 11625 36474
rect 11625 36422 11671 36474
rect 11375 36420 11431 36422
rect 11455 36420 11511 36422
rect 11535 36420 11591 36422
rect 11615 36420 11671 36422
rect 14848 45722 14904 45724
rect 14928 45722 14984 45724
rect 15008 45722 15064 45724
rect 15088 45722 15144 45724
rect 14848 45670 14894 45722
rect 14894 45670 14904 45722
rect 14928 45670 14958 45722
rect 14958 45670 14970 45722
rect 14970 45670 14984 45722
rect 15008 45670 15022 45722
rect 15022 45670 15034 45722
rect 15034 45670 15064 45722
rect 15088 45670 15098 45722
rect 15098 45670 15144 45722
rect 14848 45668 14904 45670
rect 14928 45668 14984 45670
rect 15008 45668 15064 45670
rect 15088 45668 15144 45670
rect 21794 45722 21850 45724
rect 21874 45722 21930 45724
rect 21954 45722 22010 45724
rect 22034 45722 22090 45724
rect 21794 45670 21840 45722
rect 21840 45670 21850 45722
rect 21874 45670 21904 45722
rect 21904 45670 21916 45722
rect 21916 45670 21930 45722
rect 21954 45670 21968 45722
rect 21968 45670 21980 45722
rect 21980 45670 22010 45722
rect 22034 45670 22044 45722
rect 22044 45670 22090 45722
rect 21794 45668 21850 45670
rect 21874 45668 21930 45670
rect 21954 45668 22010 45670
rect 22034 45668 22090 45670
rect 18321 45178 18377 45180
rect 18401 45178 18457 45180
rect 18481 45178 18537 45180
rect 18561 45178 18617 45180
rect 18321 45126 18367 45178
rect 18367 45126 18377 45178
rect 18401 45126 18431 45178
rect 18431 45126 18443 45178
rect 18443 45126 18457 45178
rect 18481 45126 18495 45178
rect 18495 45126 18507 45178
rect 18507 45126 18537 45178
rect 18561 45126 18571 45178
rect 18571 45126 18617 45178
rect 18321 45124 18377 45126
rect 18401 45124 18457 45126
rect 18481 45124 18537 45126
rect 18561 45124 18617 45126
rect 14848 44634 14904 44636
rect 14928 44634 14984 44636
rect 15008 44634 15064 44636
rect 15088 44634 15144 44636
rect 14848 44582 14894 44634
rect 14894 44582 14904 44634
rect 14928 44582 14958 44634
rect 14958 44582 14970 44634
rect 14970 44582 14984 44634
rect 15008 44582 15022 44634
rect 15022 44582 15034 44634
rect 15034 44582 15064 44634
rect 15088 44582 15098 44634
rect 15098 44582 15144 44634
rect 14848 44580 14904 44582
rect 14928 44580 14984 44582
rect 15008 44580 15064 44582
rect 15088 44580 15144 44582
rect 18321 44090 18377 44092
rect 18401 44090 18457 44092
rect 18481 44090 18537 44092
rect 18561 44090 18617 44092
rect 18321 44038 18367 44090
rect 18367 44038 18377 44090
rect 18401 44038 18431 44090
rect 18431 44038 18443 44090
rect 18443 44038 18457 44090
rect 18481 44038 18495 44090
rect 18495 44038 18507 44090
rect 18507 44038 18537 44090
rect 18561 44038 18571 44090
rect 18571 44038 18617 44090
rect 18321 44036 18377 44038
rect 18401 44036 18457 44038
rect 18481 44036 18537 44038
rect 18561 44036 18617 44038
rect 14848 43546 14904 43548
rect 14928 43546 14984 43548
rect 15008 43546 15064 43548
rect 15088 43546 15144 43548
rect 14848 43494 14894 43546
rect 14894 43494 14904 43546
rect 14928 43494 14958 43546
rect 14958 43494 14970 43546
rect 14970 43494 14984 43546
rect 15008 43494 15022 43546
rect 15022 43494 15034 43546
rect 15034 43494 15064 43546
rect 15088 43494 15098 43546
rect 15098 43494 15144 43546
rect 14848 43492 14904 43494
rect 14928 43492 14984 43494
rect 15008 43492 15064 43494
rect 15088 43492 15144 43494
rect 18321 43002 18377 43004
rect 18401 43002 18457 43004
rect 18481 43002 18537 43004
rect 18561 43002 18617 43004
rect 18321 42950 18367 43002
rect 18367 42950 18377 43002
rect 18401 42950 18431 43002
rect 18431 42950 18443 43002
rect 18443 42950 18457 43002
rect 18481 42950 18495 43002
rect 18495 42950 18507 43002
rect 18507 42950 18537 43002
rect 18561 42950 18571 43002
rect 18571 42950 18617 43002
rect 18321 42948 18377 42950
rect 18401 42948 18457 42950
rect 18481 42948 18537 42950
rect 18561 42948 18617 42950
rect 14848 42458 14904 42460
rect 14928 42458 14984 42460
rect 15008 42458 15064 42460
rect 15088 42458 15144 42460
rect 14848 42406 14894 42458
rect 14894 42406 14904 42458
rect 14928 42406 14958 42458
rect 14958 42406 14970 42458
rect 14970 42406 14984 42458
rect 15008 42406 15022 42458
rect 15022 42406 15034 42458
rect 15034 42406 15064 42458
rect 15088 42406 15098 42458
rect 15098 42406 15144 42458
rect 14848 42404 14904 42406
rect 14928 42404 14984 42406
rect 15008 42404 15064 42406
rect 15088 42404 15144 42406
rect 18321 41914 18377 41916
rect 18401 41914 18457 41916
rect 18481 41914 18537 41916
rect 18561 41914 18617 41916
rect 18321 41862 18367 41914
rect 18367 41862 18377 41914
rect 18401 41862 18431 41914
rect 18431 41862 18443 41914
rect 18443 41862 18457 41914
rect 18481 41862 18495 41914
rect 18495 41862 18507 41914
rect 18507 41862 18537 41914
rect 18561 41862 18571 41914
rect 18571 41862 18617 41914
rect 18321 41860 18377 41862
rect 18401 41860 18457 41862
rect 18481 41860 18537 41862
rect 18561 41860 18617 41862
rect 14848 41370 14904 41372
rect 14928 41370 14984 41372
rect 15008 41370 15064 41372
rect 15088 41370 15144 41372
rect 14848 41318 14894 41370
rect 14894 41318 14904 41370
rect 14928 41318 14958 41370
rect 14958 41318 14970 41370
rect 14970 41318 14984 41370
rect 15008 41318 15022 41370
rect 15022 41318 15034 41370
rect 15034 41318 15064 41370
rect 15088 41318 15098 41370
rect 15098 41318 15144 41370
rect 14848 41316 14904 41318
rect 14928 41316 14984 41318
rect 15008 41316 15064 41318
rect 15088 41316 15144 41318
rect 18321 40826 18377 40828
rect 18401 40826 18457 40828
rect 18481 40826 18537 40828
rect 18561 40826 18617 40828
rect 18321 40774 18367 40826
rect 18367 40774 18377 40826
rect 18401 40774 18431 40826
rect 18431 40774 18443 40826
rect 18443 40774 18457 40826
rect 18481 40774 18495 40826
rect 18495 40774 18507 40826
rect 18507 40774 18537 40826
rect 18561 40774 18571 40826
rect 18571 40774 18617 40826
rect 18321 40772 18377 40774
rect 18401 40772 18457 40774
rect 18481 40772 18537 40774
rect 18561 40772 18617 40774
rect 14848 40282 14904 40284
rect 14928 40282 14984 40284
rect 15008 40282 15064 40284
rect 15088 40282 15144 40284
rect 14848 40230 14894 40282
rect 14894 40230 14904 40282
rect 14928 40230 14958 40282
rect 14958 40230 14970 40282
rect 14970 40230 14984 40282
rect 15008 40230 15022 40282
rect 15022 40230 15034 40282
rect 15034 40230 15064 40282
rect 15088 40230 15098 40282
rect 15098 40230 15144 40282
rect 14848 40228 14904 40230
rect 14928 40228 14984 40230
rect 15008 40228 15064 40230
rect 15088 40228 15144 40230
rect 18321 39738 18377 39740
rect 18401 39738 18457 39740
rect 18481 39738 18537 39740
rect 18561 39738 18617 39740
rect 18321 39686 18367 39738
rect 18367 39686 18377 39738
rect 18401 39686 18431 39738
rect 18431 39686 18443 39738
rect 18443 39686 18457 39738
rect 18481 39686 18495 39738
rect 18495 39686 18507 39738
rect 18507 39686 18537 39738
rect 18561 39686 18571 39738
rect 18571 39686 18617 39738
rect 18321 39684 18377 39686
rect 18401 39684 18457 39686
rect 18481 39684 18537 39686
rect 18561 39684 18617 39686
rect 14848 39194 14904 39196
rect 14928 39194 14984 39196
rect 15008 39194 15064 39196
rect 15088 39194 15144 39196
rect 14848 39142 14894 39194
rect 14894 39142 14904 39194
rect 14928 39142 14958 39194
rect 14958 39142 14970 39194
rect 14970 39142 14984 39194
rect 15008 39142 15022 39194
rect 15022 39142 15034 39194
rect 15034 39142 15064 39194
rect 15088 39142 15098 39194
rect 15098 39142 15144 39194
rect 14848 39140 14904 39142
rect 14928 39140 14984 39142
rect 15008 39140 15064 39142
rect 15088 39140 15144 39142
rect 18321 38650 18377 38652
rect 18401 38650 18457 38652
rect 18481 38650 18537 38652
rect 18561 38650 18617 38652
rect 18321 38598 18367 38650
rect 18367 38598 18377 38650
rect 18401 38598 18431 38650
rect 18431 38598 18443 38650
rect 18443 38598 18457 38650
rect 18481 38598 18495 38650
rect 18495 38598 18507 38650
rect 18507 38598 18537 38650
rect 18561 38598 18571 38650
rect 18571 38598 18617 38650
rect 18321 38596 18377 38598
rect 18401 38596 18457 38598
rect 18481 38596 18537 38598
rect 18561 38596 18617 38598
rect 14848 38106 14904 38108
rect 14928 38106 14984 38108
rect 15008 38106 15064 38108
rect 15088 38106 15144 38108
rect 14848 38054 14894 38106
rect 14894 38054 14904 38106
rect 14928 38054 14958 38106
rect 14958 38054 14970 38106
rect 14970 38054 14984 38106
rect 15008 38054 15022 38106
rect 15022 38054 15034 38106
rect 15034 38054 15064 38106
rect 15088 38054 15098 38106
rect 15098 38054 15144 38106
rect 14848 38052 14904 38054
rect 14928 38052 14984 38054
rect 15008 38052 15064 38054
rect 15088 38052 15144 38054
rect 14848 37018 14904 37020
rect 14928 37018 14984 37020
rect 15008 37018 15064 37020
rect 15088 37018 15144 37020
rect 14848 36966 14894 37018
rect 14894 36966 14904 37018
rect 14928 36966 14958 37018
rect 14958 36966 14970 37018
rect 14970 36966 14984 37018
rect 15008 36966 15022 37018
rect 15022 36966 15034 37018
rect 15034 36966 15064 37018
rect 15088 36966 15098 37018
rect 15098 36966 15144 37018
rect 14848 36964 14904 36966
rect 14928 36964 14984 36966
rect 15008 36964 15064 36966
rect 15088 36964 15144 36966
rect 14848 35930 14904 35932
rect 14928 35930 14984 35932
rect 15008 35930 15064 35932
rect 15088 35930 15144 35932
rect 14848 35878 14894 35930
rect 14894 35878 14904 35930
rect 14928 35878 14958 35930
rect 14958 35878 14970 35930
rect 14970 35878 14984 35930
rect 15008 35878 15022 35930
rect 15022 35878 15034 35930
rect 15034 35878 15064 35930
rect 15088 35878 15098 35930
rect 15098 35878 15144 35930
rect 14848 35876 14904 35878
rect 14928 35876 14984 35878
rect 15008 35876 15064 35878
rect 15088 35876 15144 35878
rect 11375 35386 11431 35388
rect 11455 35386 11511 35388
rect 11535 35386 11591 35388
rect 11615 35386 11671 35388
rect 11375 35334 11421 35386
rect 11421 35334 11431 35386
rect 11455 35334 11485 35386
rect 11485 35334 11497 35386
rect 11497 35334 11511 35386
rect 11535 35334 11549 35386
rect 11549 35334 11561 35386
rect 11561 35334 11591 35386
rect 11615 35334 11625 35386
rect 11625 35334 11671 35386
rect 11375 35332 11431 35334
rect 11455 35332 11511 35334
rect 11535 35332 11591 35334
rect 11615 35332 11671 35334
rect 14848 34842 14904 34844
rect 14928 34842 14984 34844
rect 15008 34842 15064 34844
rect 15088 34842 15144 34844
rect 14848 34790 14894 34842
rect 14894 34790 14904 34842
rect 14928 34790 14958 34842
rect 14958 34790 14970 34842
rect 14970 34790 14984 34842
rect 15008 34790 15022 34842
rect 15022 34790 15034 34842
rect 15034 34790 15064 34842
rect 15088 34790 15098 34842
rect 15098 34790 15144 34842
rect 14848 34788 14904 34790
rect 14928 34788 14984 34790
rect 15008 34788 15064 34790
rect 15088 34788 15144 34790
rect 11375 34298 11431 34300
rect 11455 34298 11511 34300
rect 11535 34298 11591 34300
rect 11615 34298 11671 34300
rect 11375 34246 11421 34298
rect 11421 34246 11431 34298
rect 11455 34246 11485 34298
rect 11485 34246 11497 34298
rect 11497 34246 11511 34298
rect 11535 34246 11549 34298
rect 11549 34246 11561 34298
rect 11561 34246 11591 34298
rect 11615 34246 11625 34298
rect 11625 34246 11671 34298
rect 11375 34244 11431 34246
rect 11455 34244 11511 34246
rect 11535 34244 11591 34246
rect 11615 34244 11671 34246
rect 11375 33210 11431 33212
rect 11455 33210 11511 33212
rect 11535 33210 11591 33212
rect 11615 33210 11671 33212
rect 11375 33158 11421 33210
rect 11421 33158 11431 33210
rect 11455 33158 11485 33210
rect 11485 33158 11497 33210
rect 11497 33158 11511 33210
rect 11535 33158 11549 33210
rect 11549 33158 11561 33210
rect 11561 33158 11591 33210
rect 11615 33158 11625 33210
rect 11625 33158 11671 33210
rect 11375 33156 11431 33158
rect 11455 33156 11511 33158
rect 11535 33156 11591 33158
rect 11615 33156 11671 33158
rect 11375 32122 11431 32124
rect 11455 32122 11511 32124
rect 11535 32122 11591 32124
rect 11615 32122 11671 32124
rect 11375 32070 11421 32122
rect 11421 32070 11431 32122
rect 11455 32070 11485 32122
rect 11485 32070 11497 32122
rect 11497 32070 11511 32122
rect 11535 32070 11549 32122
rect 11549 32070 11561 32122
rect 11561 32070 11591 32122
rect 11615 32070 11625 32122
rect 11625 32070 11671 32122
rect 11375 32068 11431 32070
rect 11455 32068 11511 32070
rect 11535 32068 11591 32070
rect 11615 32068 11671 32070
rect 11375 31034 11431 31036
rect 11455 31034 11511 31036
rect 11535 31034 11591 31036
rect 11615 31034 11671 31036
rect 11375 30982 11421 31034
rect 11421 30982 11431 31034
rect 11455 30982 11485 31034
rect 11485 30982 11497 31034
rect 11497 30982 11511 31034
rect 11535 30982 11549 31034
rect 11549 30982 11561 31034
rect 11561 30982 11591 31034
rect 11615 30982 11625 31034
rect 11625 30982 11671 31034
rect 11375 30980 11431 30982
rect 11455 30980 11511 30982
rect 11535 30980 11591 30982
rect 11615 30980 11671 30982
rect 11375 29946 11431 29948
rect 11455 29946 11511 29948
rect 11535 29946 11591 29948
rect 11615 29946 11671 29948
rect 11375 29894 11421 29946
rect 11421 29894 11431 29946
rect 11455 29894 11485 29946
rect 11485 29894 11497 29946
rect 11497 29894 11511 29946
rect 11535 29894 11549 29946
rect 11549 29894 11561 29946
rect 11561 29894 11591 29946
rect 11615 29894 11625 29946
rect 11625 29894 11671 29946
rect 11375 29892 11431 29894
rect 11455 29892 11511 29894
rect 11535 29892 11591 29894
rect 11615 29892 11671 29894
rect 11375 28858 11431 28860
rect 11455 28858 11511 28860
rect 11535 28858 11591 28860
rect 11615 28858 11671 28860
rect 11375 28806 11421 28858
rect 11421 28806 11431 28858
rect 11455 28806 11485 28858
rect 11485 28806 11497 28858
rect 11497 28806 11511 28858
rect 11535 28806 11549 28858
rect 11549 28806 11561 28858
rect 11561 28806 11591 28858
rect 11615 28806 11625 28858
rect 11625 28806 11671 28858
rect 11375 28804 11431 28806
rect 11455 28804 11511 28806
rect 11535 28804 11591 28806
rect 11615 28804 11671 28806
rect 11375 27770 11431 27772
rect 11455 27770 11511 27772
rect 11535 27770 11591 27772
rect 11615 27770 11671 27772
rect 11375 27718 11421 27770
rect 11421 27718 11431 27770
rect 11455 27718 11485 27770
rect 11485 27718 11497 27770
rect 11497 27718 11511 27770
rect 11535 27718 11549 27770
rect 11549 27718 11561 27770
rect 11561 27718 11591 27770
rect 11615 27718 11625 27770
rect 11625 27718 11671 27770
rect 11375 27716 11431 27718
rect 11455 27716 11511 27718
rect 11535 27716 11591 27718
rect 11615 27716 11671 27718
rect 11375 26682 11431 26684
rect 11455 26682 11511 26684
rect 11535 26682 11591 26684
rect 11615 26682 11671 26684
rect 11375 26630 11421 26682
rect 11421 26630 11431 26682
rect 11455 26630 11485 26682
rect 11485 26630 11497 26682
rect 11497 26630 11511 26682
rect 11535 26630 11549 26682
rect 11549 26630 11561 26682
rect 11561 26630 11591 26682
rect 11615 26630 11625 26682
rect 11625 26630 11671 26682
rect 11375 26628 11431 26630
rect 11455 26628 11511 26630
rect 11535 26628 11591 26630
rect 11615 26628 11671 26630
rect 11375 25594 11431 25596
rect 11455 25594 11511 25596
rect 11535 25594 11591 25596
rect 11615 25594 11671 25596
rect 11375 25542 11421 25594
rect 11421 25542 11431 25594
rect 11455 25542 11485 25594
rect 11485 25542 11497 25594
rect 11497 25542 11511 25594
rect 11535 25542 11549 25594
rect 11549 25542 11561 25594
rect 11561 25542 11591 25594
rect 11615 25542 11625 25594
rect 11625 25542 11671 25594
rect 11375 25540 11431 25542
rect 11455 25540 11511 25542
rect 11535 25540 11591 25542
rect 11615 25540 11671 25542
rect 11375 24506 11431 24508
rect 11455 24506 11511 24508
rect 11535 24506 11591 24508
rect 11615 24506 11671 24508
rect 11375 24454 11421 24506
rect 11421 24454 11431 24506
rect 11455 24454 11485 24506
rect 11485 24454 11497 24506
rect 11497 24454 11511 24506
rect 11535 24454 11549 24506
rect 11549 24454 11561 24506
rect 11561 24454 11591 24506
rect 11615 24454 11625 24506
rect 11625 24454 11671 24506
rect 11375 24452 11431 24454
rect 11455 24452 11511 24454
rect 11535 24452 11591 24454
rect 11615 24452 11671 24454
rect 11375 23418 11431 23420
rect 11455 23418 11511 23420
rect 11535 23418 11591 23420
rect 11615 23418 11671 23420
rect 11375 23366 11421 23418
rect 11421 23366 11431 23418
rect 11455 23366 11485 23418
rect 11485 23366 11497 23418
rect 11497 23366 11511 23418
rect 11535 23366 11549 23418
rect 11549 23366 11561 23418
rect 11561 23366 11591 23418
rect 11615 23366 11625 23418
rect 11625 23366 11671 23418
rect 11375 23364 11431 23366
rect 11455 23364 11511 23366
rect 11535 23364 11591 23366
rect 11615 23364 11671 23366
rect 11375 22330 11431 22332
rect 11455 22330 11511 22332
rect 11535 22330 11591 22332
rect 11615 22330 11671 22332
rect 11375 22278 11421 22330
rect 11421 22278 11431 22330
rect 11455 22278 11485 22330
rect 11485 22278 11497 22330
rect 11497 22278 11511 22330
rect 11535 22278 11549 22330
rect 11549 22278 11561 22330
rect 11561 22278 11591 22330
rect 11615 22278 11625 22330
rect 11625 22278 11671 22330
rect 11375 22276 11431 22278
rect 11455 22276 11511 22278
rect 11535 22276 11591 22278
rect 11615 22276 11671 22278
rect 11375 21242 11431 21244
rect 11455 21242 11511 21244
rect 11535 21242 11591 21244
rect 11615 21242 11671 21244
rect 11375 21190 11421 21242
rect 11421 21190 11431 21242
rect 11455 21190 11485 21242
rect 11485 21190 11497 21242
rect 11497 21190 11511 21242
rect 11535 21190 11549 21242
rect 11549 21190 11561 21242
rect 11561 21190 11591 21242
rect 11615 21190 11625 21242
rect 11625 21190 11671 21242
rect 11375 21188 11431 21190
rect 11455 21188 11511 21190
rect 11535 21188 11591 21190
rect 11615 21188 11671 21190
rect 14848 33754 14904 33756
rect 14928 33754 14984 33756
rect 15008 33754 15064 33756
rect 15088 33754 15144 33756
rect 14848 33702 14894 33754
rect 14894 33702 14904 33754
rect 14928 33702 14958 33754
rect 14958 33702 14970 33754
rect 14970 33702 14984 33754
rect 15008 33702 15022 33754
rect 15022 33702 15034 33754
rect 15034 33702 15064 33754
rect 15088 33702 15098 33754
rect 15098 33702 15144 33754
rect 14848 33700 14904 33702
rect 14928 33700 14984 33702
rect 15008 33700 15064 33702
rect 15088 33700 15144 33702
rect 14848 32666 14904 32668
rect 14928 32666 14984 32668
rect 15008 32666 15064 32668
rect 15088 32666 15144 32668
rect 14848 32614 14894 32666
rect 14894 32614 14904 32666
rect 14928 32614 14958 32666
rect 14958 32614 14970 32666
rect 14970 32614 14984 32666
rect 15008 32614 15022 32666
rect 15022 32614 15034 32666
rect 15034 32614 15064 32666
rect 15088 32614 15098 32666
rect 15098 32614 15144 32666
rect 14848 32612 14904 32614
rect 14928 32612 14984 32614
rect 15008 32612 15064 32614
rect 15088 32612 15144 32614
rect 18321 37562 18377 37564
rect 18401 37562 18457 37564
rect 18481 37562 18537 37564
rect 18561 37562 18617 37564
rect 18321 37510 18367 37562
rect 18367 37510 18377 37562
rect 18401 37510 18431 37562
rect 18431 37510 18443 37562
rect 18443 37510 18457 37562
rect 18481 37510 18495 37562
rect 18495 37510 18507 37562
rect 18507 37510 18537 37562
rect 18561 37510 18571 37562
rect 18571 37510 18617 37562
rect 18321 37508 18377 37510
rect 18401 37508 18457 37510
rect 18481 37508 18537 37510
rect 18561 37508 18617 37510
rect 14848 31578 14904 31580
rect 14928 31578 14984 31580
rect 15008 31578 15064 31580
rect 15088 31578 15144 31580
rect 14848 31526 14894 31578
rect 14894 31526 14904 31578
rect 14928 31526 14958 31578
rect 14958 31526 14970 31578
rect 14970 31526 14984 31578
rect 15008 31526 15022 31578
rect 15022 31526 15034 31578
rect 15034 31526 15064 31578
rect 15088 31526 15098 31578
rect 15098 31526 15144 31578
rect 14848 31524 14904 31526
rect 14928 31524 14984 31526
rect 15008 31524 15064 31526
rect 15088 31524 15144 31526
rect 14848 30490 14904 30492
rect 14928 30490 14984 30492
rect 15008 30490 15064 30492
rect 15088 30490 15144 30492
rect 14848 30438 14894 30490
rect 14894 30438 14904 30490
rect 14928 30438 14958 30490
rect 14958 30438 14970 30490
rect 14970 30438 14984 30490
rect 15008 30438 15022 30490
rect 15022 30438 15034 30490
rect 15034 30438 15064 30490
rect 15088 30438 15098 30490
rect 15098 30438 15144 30490
rect 14848 30436 14904 30438
rect 14928 30436 14984 30438
rect 15008 30436 15064 30438
rect 15088 30436 15144 30438
rect 14848 29402 14904 29404
rect 14928 29402 14984 29404
rect 15008 29402 15064 29404
rect 15088 29402 15144 29404
rect 14848 29350 14894 29402
rect 14894 29350 14904 29402
rect 14928 29350 14958 29402
rect 14958 29350 14970 29402
rect 14970 29350 14984 29402
rect 15008 29350 15022 29402
rect 15022 29350 15034 29402
rect 15034 29350 15064 29402
rect 15088 29350 15098 29402
rect 15098 29350 15144 29402
rect 14848 29348 14904 29350
rect 14928 29348 14984 29350
rect 15008 29348 15064 29350
rect 15088 29348 15144 29350
rect 14848 28314 14904 28316
rect 14928 28314 14984 28316
rect 15008 28314 15064 28316
rect 15088 28314 15144 28316
rect 14848 28262 14894 28314
rect 14894 28262 14904 28314
rect 14928 28262 14958 28314
rect 14958 28262 14970 28314
rect 14970 28262 14984 28314
rect 15008 28262 15022 28314
rect 15022 28262 15034 28314
rect 15034 28262 15064 28314
rect 15088 28262 15098 28314
rect 15098 28262 15144 28314
rect 14848 28260 14904 28262
rect 14928 28260 14984 28262
rect 15008 28260 15064 28262
rect 15088 28260 15144 28262
rect 14848 27226 14904 27228
rect 14928 27226 14984 27228
rect 15008 27226 15064 27228
rect 15088 27226 15144 27228
rect 14848 27174 14894 27226
rect 14894 27174 14904 27226
rect 14928 27174 14958 27226
rect 14958 27174 14970 27226
rect 14970 27174 14984 27226
rect 15008 27174 15022 27226
rect 15022 27174 15034 27226
rect 15034 27174 15064 27226
rect 15088 27174 15098 27226
rect 15098 27174 15144 27226
rect 14848 27172 14904 27174
rect 14928 27172 14984 27174
rect 15008 27172 15064 27174
rect 15088 27172 15144 27174
rect 14848 26138 14904 26140
rect 14928 26138 14984 26140
rect 15008 26138 15064 26140
rect 15088 26138 15144 26140
rect 14848 26086 14894 26138
rect 14894 26086 14904 26138
rect 14928 26086 14958 26138
rect 14958 26086 14970 26138
rect 14970 26086 14984 26138
rect 15008 26086 15022 26138
rect 15022 26086 15034 26138
rect 15034 26086 15064 26138
rect 15088 26086 15098 26138
rect 15098 26086 15144 26138
rect 14848 26084 14904 26086
rect 14928 26084 14984 26086
rect 15008 26084 15064 26086
rect 15088 26084 15144 26086
rect 14848 25050 14904 25052
rect 14928 25050 14984 25052
rect 15008 25050 15064 25052
rect 15088 25050 15144 25052
rect 14848 24998 14894 25050
rect 14894 24998 14904 25050
rect 14928 24998 14958 25050
rect 14958 24998 14970 25050
rect 14970 24998 14984 25050
rect 15008 24998 15022 25050
rect 15022 24998 15034 25050
rect 15034 24998 15064 25050
rect 15088 24998 15098 25050
rect 15098 24998 15144 25050
rect 14848 24996 14904 24998
rect 14928 24996 14984 24998
rect 15008 24996 15064 24998
rect 15088 24996 15144 24998
rect 14848 23962 14904 23964
rect 14928 23962 14984 23964
rect 15008 23962 15064 23964
rect 15088 23962 15144 23964
rect 14848 23910 14894 23962
rect 14894 23910 14904 23962
rect 14928 23910 14958 23962
rect 14958 23910 14970 23962
rect 14970 23910 14984 23962
rect 15008 23910 15022 23962
rect 15022 23910 15034 23962
rect 15034 23910 15064 23962
rect 15088 23910 15098 23962
rect 15098 23910 15144 23962
rect 14848 23908 14904 23910
rect 14928 23908 14984 23910
rect 15008 23908 15064 23910
rect 15088 23908 15144 23910
rect 14848 22874 14904 22876
rect 14928 22874 14984 22876
rect 15008 22874 15064 22876
rect 15088 22874 15144 22876
rect 14848 22822 14894 22874
rect 14894 22822 14904 22874
rect 14928 22822 14958 22874
rect 14958 22822 14970 22874
rect 14970 22822 14984 22874
rect 15008 22822 15022 22874
rect 15022 22822 15034 22874
rect 15034 22822 15064 22874
rect 15088 22822 15098 22874
rect 15098 22822 15144 22874
rect 14848 22820 14904 22822
rect 14928 22820 14984 22822
rect 15008 22820 15064 22822
rect 15088 22820 15144 22822
rect 18321 36474 18377 36476
rect 18401 36474 18457 36476
rect 18481 36474 18537 36476
rect 18561 36474 18617 36476
rect 18321 36422 18367 36474
rect 18367 36422 18377 36474
rect 18401 36422 18431 36474
rect 18431 36422 18443 36474
rect 18443 36422 18457 36474
rect 18481 36422 18495 36474
rect 18495 36422 18507 36474
rect 18507 36422 18537 36474
rect 18561 36422 18571 36474
rect 18571 36422 18617 36474
rect 18321 36420 18377 36422
rect 18401 36420 18457 36422
rect 18481 36420 18537 36422
rect 18561 36420 18617 36422
rect 19522 38392 19578 38448
rect 18321 35386 18377 35388
rect 18401 35386 18457 35388
rect 18481 35386 18537 35388
rect 18561 35386 18617 35388
rect 18321 35334 18367 35386
rect 18367 35334 18377 35386
rect 18401 35334 18431 35386
rect 18431 35334 18443 35386
rect 18443 35334 18457 35386
rect 18481 35334 18495 35386
rect 18495 35334 18507 35386
rect 18507 35334 18537 35386
rect 18561 35334 18571 35386
rect 18571 35334 18617 35386
rect 18321 35332 18377 35334
rect 18401 35332 18457 35334
rect 18481 35332 18537 35334
rect 18561 35332 18617 35334
rect 18321 34298 18377 34300
rect 18401 34298 18457 34300
rect 18481 34298 18537 34300
rect 18561 34298 18617 34300
rect 18321 34246 18367 34298
rect 18367 34246 18377 34298
rect 18401 34246 18431 34298
rect 18431 34246 18443 34298
rect 18443 34246 18457 34298
rect 18481 34246 18495 34298
rect 18495 34246 18507 34298
rect 18507 34246 18537 34298
rect 18561 34246 18571 34298
rect 18571 34246 18617 34298
rect 18321 34244 18377 34246
rect 18401 34244 18457 34246
rect 18481 34244 18537 34246
rect 18561 34244 18617 34246
rect 18321 33210 18377 33212
rect 18401 33210 18457 33212
rect 18481 33210 18537 33212
rect 18561 33210 18617 33212
rect 18321 33158 18367 33210
rect 18367 33158 18377 33210
rect 18401 33158 18431 33210
rect 18431 33158 18443 33210
rect 18443 33158 18457 33210
rect 18481 33158 18495 33210
rect 18495 33158 18507 33210
rect 18507 33158 18537 33210
rect 18561 33158 18571 33210
rect 18571 33158 18617 33210
rect 18321 33156 18377 33158
rect 18401 33156 18457 33158
rect 18481 33156 18537 33158
rect 18561 33156 18617 33158
rect 26606 49000 26662 49056
rect 25267 47354 25323 47356
rect 25347 47354 25403 47356
rect 25427 47354 25483 47356
rect 25507 47354 25563 47356
rect 25267 47302 25313 47354
rect 25313 47302 25323 47354
rect 25347 47302 25377 47354
rect 25377 47302 25389 47354
rect 25389 47302 25403 47354
rect 25427 47302 25441 47354
rect 25441 47302 25453 47354
rect 25453 47302 25483 47354
rect 25507 47302 25517 47354
rect 25517 47302 25563 47354
rect 25267 47300 25323 47302
rect 25347 47300 25403 47302
rect 25427 47300 25483 47302
rect 25507 47300 25563 47302
rect 21794 44634 21850 44636
rect 21874 44634 21930 44636
rect 21954 44634 22010 44636
rect 22034 44634 22090 44636
rect 21794 44582 21840 44634
rect 21840 44582 21850 44634
rect 21874 44582 21904 44634
rect 21904 44582 21916 44634
rect 21916 44582 21930 44634
rect 21954 44582 21968 44634
rect 21968 44582 21980 44634
rect 21980 44582 22010 44634
rect 22034 44582 22044 44634
rect 22044 44582 22090 44634
rect 21794 44580 21850 44582
rect 21874 44580 21930 44582
rect 21954 44580 22010 44582
rect 22034 44580 22090 44582
rect 21794 43546 21850 43548
rect 21874 43546 21930 43548
rect 21954 43546 22010 43548
rect 22034 43546 22090 43548
rect 21794 43494 21840 43546
rect 21840 43494 21850 43546
rect 21874 43494 21904 43546
rect 21904 43494 21916 43546
rect 21916 43494 21930 43546
rect 21954 43494 21968 43546
rect 21968 43494 21980 43546
rect 21980 43494 22010 43546
rect 22034 43494 22044 43546
rect 22044 43494 22090 43546
rect 21794 43492 21850 43494
rect 21874 43492 21930 43494
rect 21954 43492 22010 43494
rect 22034 43492 22090 43494
rect 21794 42458 21850 42460
rect 21874 42458 21930 42460
rect 21954 42458 22010 42460
rect 22034 42458 22090 42460
rect 21794 42406 21840 42458
rect 21840 42406 21850 42458
rect 21874 42406 21904 42458
rect 21904 42406 21916 42458
rect 21916 42406 21930 42458
rect 21954 42406 21968 42458
rect 21968 42406 21980 42458
rect 21980 42406 22010 42458
rect 22034 42406 22044 42458
rect 22044 42406 22090 42458
rect 21794 42404 21850 42406
rect 21874 42404 21930 42406
rect 21954 42404 22010 42406
rect 22034 42404 22090 42406
rect 21794 41370 21850 41372
rect 21874 41370 21930 41372
rect 21954 41370 22010 41372
rect 22034 41370 22090 41372
rect 21794 41318 21840 41370
rect 21840 41318 21850 41370
rect 21874 41318 21904 41370
rect 21904 41318 21916 41370
rect 21916 41318 21930 41370
rect 21954 41318 21968 41370
rect 21968 41318 21980 41370
rect 21980 41318 22010 41370
rect 22034 41318 22044 41370
rect 22044 41318 22090 41370
rect 21794 41316 21850 41318
rect 21874 41316 21930 41318
rect 21954 41316 22010 41318
rect 22034 41316 22090 41318
rect 21794 40282 21850 40284
rect 21874 40282 21930 40284
rect 21954 40282 22010 40284
rect 22034 40282 22090 40284
rect 21794 40230 21840 40282
rect 21840 40230 21850 40282
rect 21874 40230 21904 40282
rect 21904 40230 21916 40282
rect 21916 40230 21930 40282
rect 21954 40230 21968 40282
rect 21968 40230 21980 40282
rect 21980 40230 22010 40282
rect 22034 40230 22044 40282
rect 22044 40230 22090 40282
rect 21794 40228 21850 40230
rect 21874 40228 21930 40230
rect 21954 40228 22010 40230
rect 22034 40228 22090 40230
rect 21794 39194 21850 39196
rect 21874 39194 21930 39196
rect 21954 39194 22010 39196
rect 22034 39194 22090 39196
rect 21794 39142 21840 39194
rect 21840 39142 21850 39194
rect 21874 39142 21904 39194
rect 21904 39142 21916 39194
rect 21916 39142 21930 39194
rect 21954 39142 21968 39194
rect 21968 39142 21980 39194
rect 21980 39142 22010 39194
rect 22034 39142 22044 39194
rect 22044 39142 22090 39194
rect 21794 39140 21850 39142
rect 21874 39140 21930 39142
rect 21954 39140 22010 39142
rect 22034 39140 22090 39142
rect 20626 38392 20682 38448
rect 21794 38106 21850 38108
rect 21874 38106 21930 38108
rect 21954 38106 22010 38108
rect 22034 38106 22090 38108
rect 21794 38054 21840 38106
rect 21840 38054 21850 38106
rect 21874 38054 21904 38106
rect 21904 38054 21916 38106
rect 21916 38054 21930 38106
rect 21954 38054 21968 38106
rect 21968 38054 21980 38106
rect 21980 38054 22010 38106
rect 22034 38054 22044 38106
rect 22044 38054 22090 38106
rect 21794 38052 21850 38054
rect 21874 38052 21930 38054
rect 21954 38052 22010 38054
rect 22034 38052 22090 38054
rect 18321 32122 18377 32124
rect 18401 32122 18457 32124
rect 18481 32122 18537 32124
rect 18561 32122 18617 32124
rect 18321 32070 18367 32122
rect 18367 32070 18377 32122
rect 18401 32070 18431 32122
rect 18431 32070 18443 32122
rect 18443 32070 18457 32122
rect 18481 32070 18495 32122
rect 18495 32070 18507 32122
rect 18507 32070 18537 32122
rect 18561 32070 18571 32122
rect 18571 32070 18617 32122
rect 18321 32068 18377 32070
rect 18401 32068 18457 32070
rect 18481 32068 18537 32070
rect 18561 32068 18617 32070
rect 14848 21786 14904 21788
rect 14928 21786 14984 21788
rect 15008 21786 15064 21788
rect 15088 21786 15144 21788
rect 14848 21734 14894 21786
rect 14894 21734 14904 21786
rect 14928 21734 14958 21786
rect 14958 21734 14970 21786
rect 14970 21734 14984 21786
rect 15008 21734 15022 21786
rect 15022 21734 15034 21786
rect 15034 21734 15064 21786
rect 15088 21734 15098 21786
rect 15098 21734 15144 21786
rect 14848 21732 14904 21734
rect 14928 21732 14984 21734
rect 15008 21732 15064 21734
rect 15088 21732 15144 21734
rect 14848 20698 14904 20700
rect 14928 20698 14984 20700
rect 15008 20698 15064 20700
rect 15088 20698 15144 20700
rect 14848 20646 14894 20698
rect 14894 20646 14904 20698
rect 14928 20646 14958 20698
rect 14958 20646 14970 20698
rect 14970 20646 14984 20698
rect 15008 20646 15022 20698
rect 15022 20646 15034 20698
rect 15034 20646 15064 20698
rect 15088 20646 15098 20698
rect 15098 20646 15144 20698
rect 14848 20644 14904 20646
rect 14928 20644 14984 20646
rect 15008 20644 15064 20646
rect 15088 20644 15144 20646
rect 11375 20154 11431 20156
rect 11455 20154 11511 20156
rect 11535 20154 11591 20156
rect 11615 20154 11671 20156
rect 11375 20102 11421 20154
rect 11421 20102 11431 20154
rect 11455 20102 11485 20154
rect 11485 20102 11497 20154
rect 11497 20102 11511 20154
rect 11535 20102 11549 20154
rect 11549 20102 11561 20154
rect 11561 20102 11591 20154
rect 11615 20102 11625 20154
rect 11625 20102 11671 20154
rect 11375 20100 11431 20102
rect 11455 20100 11511 20102
rect 11535 20100 11591 20102
rect 11615 20100 11671 20102
rect 11375 19066 11431 19068
rect 11455 19066 11511 19068
rect 11535 19066 11591 19068
rect 11615 19066 11671 19068
rect 11375 19014 11421 19066
rect 11421 19014 11431 19066
rect 11455 19014 11485 19066
rect 11485 19014 11497 19066
rect 11497 19014 11511 19066
rect 11535 19014 11549 19066
rect 11549 19014 11561 19066
rect 11561 19014 11591 19066
rect 11615 19014 11625 19066
rect 11625 19014 11671 19066
rect 11375 19012 11431 19014
rect 11455 19012 11511 19014
rect 11535 19012 11591 19014
rect 11615 19012 11671 19014
rect 11375 17978 11431 17980
rect 11455 17978 11511 17980
rect 11535 17978 11591 17980
rect 11615 17978 11671 17980
rect 11375 17926 11421 17978
rect 11421 17926 11431 17978
rect 11455 17926 11485 17978
rect 11485 17926 11497 17978
rect 11497 17926 11511 17978
rect 11535 17926 11549 17978
rect 11549 17926 11561 17978
rect 11561 17926 11591 17978
rect 11615 17926 11625 17978
rect 11625 17926 11671 17978
rect 11375 17924 11431 17926
rect 11455 17924 11511 17926
rect 11535 17924 11591 17926
rect 11615 17924 11671 17926
rect 11375 16890 11431 16892
rect 11455 16890 11511 16892
rect 11535 16890 11591 16892
rect 11615 16890 11671 16892
rect 11375 16838 11421 16890
rect 11421 16838 11431 16890
rect 11455 16838 11485 16890
rect 11485 16838 11497 16890
rect 11497 16838 11511 16890
rect 11535 16838 11549 16890
rect 11549 16838 11561 16890
rect 11561 16838 11591 16890
rect 11615 16838 11625 16890
rect 11625 16838 11671 16890
rect 11375 16836 11431 16838
rect 11455 16836 11511 16838
rect 11535 16836 11591 16838
rect 11615 16836 11671 16838
rect 11375 15802 11431 15804
rect 11455 15802 11511 15804
rect 11535 15802 11591 15804
rect 11615 15802 11671 15804
rect 11375 15750 11421 15802
rect 11421 15750 11431 15802
rect 11455 15750 11485 15802
rect 11485 15750 11497 15802
rect 11497 15750 11511 15802
rect 11535 15750 11549 15802
rect 11549 15750 11561 15802
rect 11561 15750 11591 15802
rect 11615 15750 11625 15802
rect 11625 15750 11671 15802
rect 11375 15748 11431 15750
rect 11455 15748 11511 15750
rect 11535 15748 11591 15750
rect 11615 15748 11671 15750
rect 11375 14714 11431 14716
rect 11455 14714 11511 14716
rect 11535 14714 11591 14716
rect 11615 14714 11671 14716
rect 11375 14662 11421 14714
rect 11421 14662 11431 14714
rect 11455 14662 11485 14714
rect 11485 14662 11497 14714
rect 11497 14662 11511 14714
rect 11535 14662 11549 14714
rect 11549 14662 11561 14714
rect 11561 14662 11591 14714
rect 11615 14662 11625 14714
rect 11625 14662 11671 14714
rect 11375 14660 11431 14662
rect 11455 14660 11511 14662
rect 11535 14660 11591 14662
rect 11615 14660 11671 14662
rect 11375 13626 11431 13628
rect 11455 13626 11511 13628
rect 11535 13626 11591 13628
rect 11615 13626 11671 13628
rect 11375 13574 11421 13626
rect 11421 13574 11431 13626
rect 11455 13574 11485 13626
rect 11485 13574 11497 13626
rect 11497 13574 11511 13626
rect 11535 13574 11549 13626
rect 11549 13574 11561 13626
rect 11561 13574 11591 13626
rect 11615 13574 11625 13626
rect 11625 13574 11671 13626
rect 11375 13572 11431 13574
rect 11455 13572 11511 13574
rect 11535 13572 11591 13574
rect 11615 13572 11671 13574
rect 11375 12538 11431 12540
rect 11455 12538 11511 12540
rect 11535 12538 11591 12540
rect 11615 12538 11671 12540
rect 11375 12486 11421 12538
rect 11421 12486 11431 12538
rect 11455 12486 11485 12538
rect 11485 12486 11497 12538
rect 11497 12486 11511 12538
rect 11535 12486 11549 12538
rect 11549 12486 11561 12538
rect 11561 12486 11591 12538
rect 11615 12486 11625 12538
rect 11625 12486 11671 12538
rect 11375 12484 11431 12486
rect 11455 12484 11511 12486
rect 11535 12484 11591 12486
rect 11615 12484 11671 12486
rect 11375 11450 11431 11452
rect 11455 11450 11511 11452
rect 11535 11450 11591 11452
rect 11615 11450 11671 11452
rect 11375 11398 11421 11450
rect 11421 11398 11431 11450
rect 11455 11398 11485 11450
rect 11485 11398 11497 11450
rect 11497 11398 11511 11450
rect 11535 11398 11549 11450
rect 11549 11398 11561 11450
rect 11561 11398 11591 11450
rect 11615 11398 11625 11450
rect 11625 11398 11671 11450
rect 11375 11396 11431 11398
rect 11455 11396 11511 11398
rect 11535 11396 11591 11398
rect 11615 11396 11671 11398
rect 11375 10362 11431 10364
rect 11455 10362 11511 10364
rect 11535 10362 11591 10364
rect 11615 10362 11671 10364
rect 11375 10310 11421 10362
rect 11421 10310 11431 10362
rect 11455 10310 11485 10362
rect 11485 10310 11497 10362
rect 11497 10310 11511 10362
rect 11535 10310 11549 10362
rect 11549 10310 11561 10362
rect 11561 10310 11591 10362
rect 11615 10310 11625 10362
rect 11625 10310 11671 10362
rect 11375 10308 11431 10310
rect 11455 10308 11511 10310
rect 11535 10308 11591 10310
rect 11615 10308 11671 10310
rect 11375 9274 11431 9276
rect 11455 9274 11511 9276
rect 11535 9274 11591 9276
rect 11615 9274 11671 9276
rect 11375 9222 11421 9274
rect 11421 9222 11431 9274
rect 11455 9222 11485 9274
rect 11485 9222 11497 9274
rect 11497 9222 11511 9274
rect 11535 9222 11549 9274
rect 11549 9222 11561 9274
rect 11561 9222 11591 9274
rect 11615 9222 11625 9274
rect 11625 9222 11671 9274
rect 11375 9220 11431 9222
rect 11455 9220 11511 9222
rect 11535 9220 11591 9222
rect 11615 9220 11671 9222
rect 11375 8186 11431 8188
rect 11455 8186 11511 8188
rect 11535 8186 11591 8188
rect 11615 8186 11671 8188
rect 11375 8134 11421 8186
rect 11421 8134 11431 8186
rect 11455 8134 11485 8186
rect 11485 8134 11497 8186
rect 11497 8134 11511 8186
rect 11535 8134 11549 8186
rect 11549 8134 11561 8186
rect 11561 8134 11591 8186
rect 11615 8134 11625 8186
rect 11625 8134 11671 8186
rect 11375 8132 11431 8134
rect 11455 8132 11511 8134
rect 11535 8132 11591 8134
rect 11615 8132 11671 8134
rect 11375 7098 11431 7100
rect 11455 7098 11511 7100
rect 11535 7098 11591 7100
rect 11615 7098 11671 7100
rect 11375 7046 11421 7098
rect 11421 7046 11431 7098
rect 11455 7046 11485 7098
rect 11485 7046 11497 7098
rect 11497 7046 11511 7098
rect 11535 7046 11549 7098
rect 11549 7046 11561 7098
rect 11561 7046 11591 7098
rect 11615 7046 11625 7098
rect 11625 7046 11671 7098
rect 11375 7044 11431 7046
rect 11455 7044 11511 7046
rect 11535 7044 11591 7046
rect 11615 7044 11671 7046
rect 11375 6010 11431 6012
rect 11455 6010 11511 6012
rect 11535 6010 11591 6012
rect 11615 6010 11671 6012
rect 11375 5958 11421 6010
rect 11421 5958 11431 6010
rect 11455 5958 11485 6010
rect 11485 5958 11497 6010
rect 11497 5958 11511 6010
rect 11535 5958 11549 6010
rect 11549 5958 11561 6010
rect 11561 5958 11591 6010
rect 11615 5958 11625 6010
rect 11625 5958 11671 6010
rect 11375 5956 11431 5958
rect 11455 5956 11511 5958
rect 11535 5956 11591 5958
rect 11615 5956 11671 5958
rect 11375 4922 11431 4924
rect 11455 4922 11511 4924
rect 11535 4922 11591 4924
rect 11615 4922 11671 4924
rect 11375 4870 11421 4922
rect 11421 4870 11431 4922
rect 11455 4870 11485 4922
rect 11485 4870 11497 4922
rect 11497 4870 11511 4922
rect 11535 4870 11549 4922
rect 11549 4870 11561 4922
rect 11561 4870 11591 4922
rect 11615 4870 11625 4922
rect 11625 4870 11671 4922
rect 11375 4868 11431 4870
rect 11455 4868 11511 4870
rect 11535 4868 11591 4870
rect 11615 4868 11671 4870
rect 11375 3834 11431 3836
rect 11455 3834 11511 3836
rect 11535 3834 11591 3836
rect 11615 3834 11671 3836
rect 11375 3782 11421 3834
rect 11421 3782 11431 3834
rect 11455 3782 11485 3834
rect 11485 3782 11497 3834
rect 11497 3782 11511 3834
rect 11535 3782 11549 3834
rect 11549 3782 11561 3834
rect 11561 3782 11591 3834
rect 11615 3782 11625 3834
rect 11625 3782 11671 3834
rect 11375 3780 11431 3782
rect 11455 3780 11511 3782
rect 11535 3780 11591 3782
rect 11615 3780 11671 3782
rect 14848 19610 14904 19612
rect 14928 19610 14984 19612
rect 15008 19610 15064 19612
rect 15088 19610 15144 19612
rect 14848 19558 14894 19610
rect 14894 19558 14904 19610
rect 14928 19558 14958 19610
rect 14958 19558 14970 19610
rect 14970 19558 14984 19610
rect 15008 19558 15022 19610
rect 15022 19558 15034 19610
rect 15034 19558 15064 19610
rect 15088 19558 15098 19610
rect 15098 19558 15144 19610
rect 14848 19556 14904 19558
rect 14928 19556 14984 19558
rect 15008 19556 15064 19558
rect 15088 19556 15144 19558
rect 14848 18522 14904 18524
rect 14928 18522 14984 18524
rect 15008 18522 15064 18524
rect 15088 18522 15144 18524
rect 14848 18470 14894 18522
rect 14894 18470 14904 18522
rect 14928 18470 14958 18522
rect 14958 18470 14970 18522
rect 14970 18470 14984 18522
rect 15008 18470 15022 18522
rect 15022 18470 15034 18522
rect 15034 18470 15064 18522
rect 15088 18470 15098 18522
rect 15098 18470 15144 18522
rect 14848 18468 14904 18470
rect 14928 18468 14984 18470
rect 15008 18468 15064 18470
rect 15088 18468 15144 18470
rect 14848 17434 14904 17436
rect 14928 17434 14984 17436
rect 15008 17434 15064 17436
rect 15088 17434 15144 17436
rect 14848 17382 14894 17434
rect 14894 17382 14904 17434
rect 14928 17382 14958 17434
rect 14958 17382 14970 17434
rect 14970 17382 14984 17434
rect 15008 17382 15022 17434
rect 15022 17382 15034 17434
rect 15034 17382 15064 17434
rect 15088 17382 15098 17434
rect 15098 17382 15144 17434
rect 14848 17380 14904 17382
rect 14928 17380 14984 17382
rect 15008 17380 15064 17382
rect 15088 17380 15144 17382
rect 11375 2746 11431 2748
rect 11455 2746 11511 2748
rect 11535 2746 11591 2748
rect 11615 2746 11671 2748
rect 11375 2694 11421 2746
rect 11421 2694 11431 2746
rect 11455 2694 11485 2746
rect 11485 2694 11497 2746
rect 11497 2694 11511 2746
rect 11535 2694 11549 2746
rect 11549 2694 11561 2746
rect 11561 2694 11591 2746
rect 11615 2694 11625 2746
rect 11625 2694 11671 2746
rect 11375 2692 11431 2694
rect 11455 2692 11511 2694
rect 11535 2692 11591 2694
rect 11615 2692 11671 2694
rect 18321 31034 18377 31036
rect 18401 31034 18457 31036
rect 18481 31034 18537 31036
rect 18561 31034 18617 31036
rect 18321 30982 18367 31034
rect 18367 30982 18377 31034
rect 18401 30982 18431 31034
rect 18431 30982 18443 31034
rect 18443 30982 18457 31034
rect 18481 30982 18495 31034
rect 18495 30982 18507 31034
rect 18507 30982 18537 31034
rect 18561 30982 18571 31034
rect 18571 30982 18617 31034
rect 18321 30980 18377 30982
rect 18401 30980 18457 30982
rect 18481 30980 18537 30982
rect 18561 30980 18617 30982
rect 18321 29946 18377 29948
rect 18401 29946 18457 29948
rect 18481 29946 18537 29948
rect 18561 29946 18617 29948
rect 18321 29894 18367 29946
rect 18367 29894 18377 29946
rect 18401 29894 18431 29946
rect 18431 29894 18443 29946
rect 18443 29894 18457 29946
rect 18481 29894 18495 29946
rect 18495 29894 18507 29946
rect 18507 29894 18537 29946
rect 18561 29894 18571 29946
rect 18571 29894 18617 29946
rect 18321 29892 18377 29894
rect 18401 29892 18457 29894
rect 18481 29892 18537 29894
rect 18561 29892 18617 29894
rect 18321 28858 18377 28860
rect 18401 28858 18457 28860
rect 18481 28858 18537 28860
rect 18561 28858 18617 28860
rect 18321 28806 18367 28858
rect 18367 28806 18377 28858
rect 18401 28806 18431 28858
rect 18431 28806 18443 28858
rect 18443 28806 18457 28858
rect 18481 28806 18495 28858
rect 18495 28806 18507 28858
rect 18507 28806 18537 28858
rect 18561 28806 18571 28858
rect 18571 28806 18617 28858
rect 18321 28804 18377 28806
rect 18401 28804 18457 28806
rect 18481 28804 18537 28806
rect 18561 28804 18617 28806
rect 18878 27940 18934 27976
rect 18878 27920 18880 27940
rect 18880 27920 18932 27940
rect 18932 27920 18934 27940
rect 18321 27770 18377 27772
rect 18401 27770 18457 27772
rect 18481 27770 18537 27772
rect 18561 27770 18617 27772
rect 18321 27718 18367 27770
rect 18367 27718 18377 27770
rect 18401 27718 18431 27770
rect 18431 27718 18443 27770
rect 18443 27718 18457 27770
rect 18481 27718 18495 27770
rect 18495 27718 18507 27770
rect 18507 27718 18537 27770
rect 18561 27718 18571 27770
rect 18571 27718 18617 27770
rect 18321 27716 18377 27718
rect 18401 27716 18457 27718
rect 18481 27716 18537 27718
rect 18561 27716 18617 27718
rect 18321 26682 18377 26684
rect 18401 26682 18457 26684
rect 18481 26682 18537 26684
rect 18561 26682 18617 26684
rect 18321 26630 18367 26682
rect 18367 26630 18377 26682
rect 18401 26630 18431 26682
rect 18431 26630 18443 26682
rect 18443 26630 18457 26682
rect 18481 26630 18495 26682
rect 18495 26630 18507 26682
rect 18507 26630 18537 26682
rect 18561 26630 18571 26682
rect 18571 26630 18617 26682
rect 18321 26628 18377 26630
rect 18401 26628 18457 26630
rect 18481 26628 18537 26630
rect 18561 26628 18617 26630
rect 14848 16346 14904 16348
rect 14928 16346 14984 16348
rect 15008 16346 15064 16348
rect 15088 16346 15144 16348
rect 14848 16294 14894 16346
rect 14894 16294 14904 16346
rect 14928 16294 14958 16346
rect 14958 16294 14970 16346
rect 14970 16294 14984 16346
rect 15008 16294 15022 16346
rect 15022 16294 15034 16346
rect 15034 16294 15064 16346
rect 15088 16294 15098 16346
rect 15098 16294 15144 16346
rect 14848 16292 14904 16294
rect 14928 16292 14984 16294
rect 15008 16292 15064 16294
rect 15088 16292 15144 16294
rect 14848 15258 14904 15260
rect 14928 15258 14984 15260
rect 15008 15258 15064 15260
rect 15088 15258 15144 15260
rect 14848 15206 14894 15258
rect 14894 15206 14904 15258
rect 14928 15206 14958 15258
rect 14958 15206 14970 15258
rect 14970 15206 14984 15258
rect 15008 15206 15022 15258
rect 15022 15206 15034 15258
rect 15034 15206 15064 15258
rect 15088 15206 15098 15258
rect 15098 15206 15144 15258
rect 14848 15204 14904 15206
rect 14928 15204 14984 15206
rect 15008 15204 15064 15206
rect 15088 15204 15144 15206
rect 14848 14170 14904 14172
rect 14928 14170 14984 14172
rect 15008 14170 15064 14172
rect 15088 14170 15144 14172
rect 14848 14118 14894 14170
rect 14894 14118 14904 14170
rect 14928 14118 14958 14170
rect 14958 14118 14970 14170
rect 14970 14118 14984 14170
rect 15008 14118 15022 14170
rect 15022 14118 15034 14170
rect 15034 14118 15064 14170
rect 15088 14118 15098 14170
rect 15098 14118 15144 14170
rect 14848 14116 14904 14118
rect 14928 14116 14984 14118
rect 15008 14116 15064 14118
rect 15088 14116 15144 14118
rect 14848 13082 14904 13084
rect 14928 13082 14984 13084
rect 15008 13082 15064 13084
rect 15088 13082 15144 13084
rect 14848 13030 14894 13082
rect 14894 13030 14904 13082
rect 14928 13030 14958 13082
rect 14958 13030 14970 13082
rect 14970 13030 14984 13082
rect 15008 13030 15022 13082
rect 15022 13030 15034 13082
rect 15034 13030 15064 13082
rect 15088 13030 15098 13082
rect 15098 13030 15144 13082
rect 14848 13028 14904 13030
rect 14928 13028 14984 13030
rect 15008 13028 15064 13030
rect 15088 13028 15144 13030
rect 18321 25594 18377 25596
rect 18401 25594 18457 25596
rect 18481 25594 18537 25596
rect 18561 25594 18617 25596
rect 18321 25542 18367 25594
rect 18367 25542 18377 25594
rect 18401 25542 18431 25594
rect 18431 25542 18443 25594
rect 18443 25542 18457 25594
rect 18481 25542 18495 25594
rect 18495 25542 18507 25594
rect 18507 25542 18537 25594
rect 18561 25542 18571 25594
rect 18571 25542 18617 25594
rect 18321 25540 18377 25542
rect 18401 25540 18457 25542
rect 18481 25540 18537 25542
rect 18561 25540 18617 25542
rect 18321 24506 18377 24508
rect 18401 24506 18457 24508
rect 18481 24506 18537 24508
rect 18561 24506 18617 24508
rect 18321 24454 18367 24506
rect 18367 24454 18377 24506
rect 18401 24454 18431 24506
rect 18431 24454 18443 24506
rect 18443 24454 18457 24506
rect 18481 24454 18495 24506
rect 18495 24454 18507 24506
rect 18507 24454 18537 24506
rect 18561 24454 18571 24506
rect 18571 24454 18617 24506
rect 18321 24452 18377 24454
rect 18401 24452 18457 24454
rect 18481 24452 18537 24454
rect 18561 24452 18617 24454
rect 18321 23418 18377 23420
rect 18401 23418 18457 23420
rect 18481 23418 18537 23420
rect 18561 23418 18617 23420
rect 18321 23366 18367 23418
rect 18367 23366 18377 23418
rect 18401 23366 18431 23418
rect 18431 23366 18443 23418
rect 18443 23366 18457 23418
rect 18481 23366 18495 23418
rect 18495 23366 18507 23418
rect 18507 23366 18537 23418
rect 18561 23366 18571 23418
rect 18571 23366 18617 23418
rect 18321 23364 18377 23366
rect 18401 23364 18457 23366
rect 18481 23364 18537 23366
rect 18561 23364 18617 23366
rect 14848 11994 14904 11996
rect 14928 11994 14984 11996
rect 15008 11994 15064 11996
rect 15088 11994 15144 11996
rect 14848 11942 14894 11994
rect 14894 11942 14904 11994
rect 14928 11942 14958 11994
rect 14958 11942 14970 11994
rect 14970 11942 14984 11994
rect 15008 11942 15022 11994
rect 15022 11942 15034 11994
rect 15034 11942 15064 11994
rect 15088 11942 15098 11994
rect 15098 11942 15144 11994
rect 14848 11940 14904 11942
rect 14928 11940 14984 11942
rect 15008 11940 15064 11942
rect 15088 11940 15144 11942
rect 14848 10906 14904 10908
rect 14928 10906 14984 10908
rect 15008 10906 15064 10908
rect 15088 10906 15144 10908
rect 14848 10854 14894 10906
rect 14894 10854 14904 10906
rect 14928 10854 14958 10906
rect 14958 10854 14970 10906
rect 14970 10854 14984 10906
rect 15008 10854 15022 10906
rect 15022 10854 15034 10906
rect 15034 10854 15064 10906
rect 15088 10854 15098 10906
rect 15098 10854 15144 10906
rect 14848 10852 14904 10854
rect 14928 10852 14984 10854
rect 15008 10852 15064 10854
rect 15088 10852 15144 10854
rect 14848 9818 14904 9820
rect 14928 9818 14984 9820
rect 15008 9818 15064 9820
rect 15088 9818 15144 9820
rect 14848 9766 14894 9818
rect 14894 9766 14904 9818
rect 14928 9766 14958 9818
rect 14958 9766 14970 9818
rect 14970 9766 14984 9818
rect 15008 9766 15022 9818
rect 15022 9766 15034 9818
rect 15034 9766 15064 9818
rect 15088 9766 15098 9818
rect 15098 9766 15144 9818
rect 14848 9764 14904 9766
rect 14928 9764 14984 9766
rect 15008 9764 15064 9766
rect 15088 9764 15144 9766
rect 14848 8730 14904 8732
rect 14928 8730 14984 8732
rect 15008 8730 15064 8732
rect 15088 8730 15144 8732
rect 14848 8678 14894 8730
rect 14894 8678 14904 8730
rect 14928 8678 14958 8730
rect 14958 8678 14970 8730
rect 14970 8678 14984 8730
rect 15008 8678 15022 8730
rect 15022 8678 15034 8730
rect 15034 8678 15064 8730
rect 15088 8678 15098 8730
rect 15098 8678 15144 8730
rect 14848 8676 14904 8678
rect 14928 8676 14984 8678
rect 15008 8676 15064 8678
rect 15088 8676 15144 8678
rect 14848 7642 14904 7644
rect 14928 7642 14984 7644
rect 15008 7642 15064 7644
rect 15088 7642 15144 7644
rect 14848 7590 14894 7642
rect 14894 7590 14904 7642
rect 14928 7590 14958 7642
rect 14958 7590 14970 7642
rect 14970 7590 14984 7642
rect 15008 7590 15022 7642
rect 15022 7590 15034 7642
rect 15034 7590 15064 7642
rect 15088 7590 15098 7642
rect 15098 7590 15144 7642
rect 14848 7588 14904 7590
rect 14928 7588 14984 7590
rect 15008 7588 15064 7590
rect 15088 7588 15144 7590
rect 14848 6554 14904 6556
rect 14928 6554 14984 6556
rect 15008 6554 15064 6556
rect 15088 6554 15144 6556
rect 14848 6502 14894 6554
rect 14894 6502 14904 6554
rect 14928 6502 14958 6554
rect 14958 6502 14970 6554
rect 14970 6502 14984 6554
rect 15008 6502 15022 6554
rect 15022 6502 15034 6554
rect 15034 6502 15064 6554
rect 15088 6502 15098 6554
rect 15098 6502 15144 6554
rect 14848 6500 14904 6502
rect 14928 6500 14984 6502
rect 15008 6500 15064 6502
rect 15088 6500 15144 6502
rect 14848 5466 14904 5468
rect 14928 5466 14984 5468
rect 15008 5466 15064 5468
rect 15088 5466 15144 5468
rect 14848 5414 14894 5466
rect 14894 5414 14904 5466
rect 14928 5414 14958 5466
rect 14958 5414 14970 5466
rect 14970 5414 14984 5466
rect 15008 5414 15022 5466
rect 15022 5414 15034 5466
rect 15034 5414 15064 5466
rect 15088 5414 15098 5466
rect 15098 5414 15144 5466
rect 14848 5412 14904 5414
rect 14928 5412 14984 5414
rect 15008 5412 15064 5414
rect 15088 5412 15144 5414
rect 14848 4378 14904 4380
rect 14928 4378 14984 4380
rect 15008 4378 15064 4380
rect 15088 4378 15144 4380
rect 14848 4326 14894 4378
rect 14894 4326 14904 4378
rect 14928 4326 14958 4378
rect 14958 4326 14970 4378
rect 14970 4326 14984 4378
rect 15008 4326 15022 4378
rect 15022 4326 15034 4378
rect 15034 4326 15064 4378
rect 15088 4326 15098 4378
rect 15098 4326 15144 4378
rect 14848 4324 14904 4326
rect 14928 4324 14984 4326
rect 15008 4324 15064 4326
rect 15088 4324 15144 4326
rect 14848 3290 14904 3292
rect 14928 3290 14984 3292
rect 15008 3290 15064 3292
rect 15088 3290 15144 3292
rect 14848 3238 14894 3290
rect 14894 3238 14904 3290
rect 14928 3238 14958 3290
rect 14958 3238 14970 3290
rect 14970 3238 14984 3290
rect 15008 3238 15022 3290
rect 15022 3238 15034 3290
rect 15034 3238 15064 3290
rect 15088 3238 15098 3290
rect 15098 3238 15144 3290
rect 14848 3236 14904 3238
rect 14928 3236 14984 3238
rect 15008 3236 15064 3238
rect 15088 3236 15144 3238
rect 14848 2202 14904 2204
rect 14928 2202 14984 2204
rect 15008 2202 15064 2204
rect 15088 2202 15144 2204
rect 14848 2150 14894 2202
rect 14894 2150 14904 2202
rect 14928 2150 14958 2202
rect 14958 2150 14970 2202
rect 14970 2150 14984 2202
rect 15008 2150 15022 2202
rect 15022 2150 15034 2202
rect 15034 2150 15064 2202
rect 15088 2150 15098 2202
rect 15098 2150 15144 2202
rect 14848 2148 14904 2150
rect 14928 2148 14984 2150
rect 15008 2148 15064 2150
rect 15088 2148 15144 2150
rect 18321 22330 18377 22332
rect 18401 22330 18457 22332
rect 18481 22330 18537 22332
rect 18561 22330 18617 22332
rect 18321 22278 18367 22330
rect 18367 22278 18377 22330
rect 18401 22278 18431 22330
rect 18431 22278 18443 22330
rect 18443 22278 18457 22330
rect 18481 22278 18495 22330
rect 18495 22278 18507 22330
rect 18507 22278 18537 22330
rect 18561 22278 18571 22330
rect 18571 22278 18617 22330
rect 18321 22276 18377 22278
rect 18401 22276 18457 22278
rect 18481 22276 18537 22278
rect 18561 22276 18617 22278
rect 18321 21242 18377 21244
rect 18401 21242 18457 21244
rect 18481 21242 18537 21244
rect 18561 21242 18617 21244
rect 18321 21190 18367 21242
rect 18367 21190 18377 21242
rect 18401 21190 18431 21242
rect 18431 21190 18443 21242
rect 18443 21190 18457 21242
rect 18481 21190 18495 21242
rect 18495 21190 18507 21242
rect 18507 21190 18537 21242
rect 18561 21190 18571 21242
rect 18571 21190 18617 21242
rect 18321 21188 18377 21190
rect 18401 21188 18457 21190
rect 18481 21188 18537 21190
rect 18561 21188 18617 21190
rect 18321 20154 18377 20156
rect 18401 20154 18457 20156
rect 18481 20154 18537 20156
rect 18561 20154 18617 20156
rect 18321 20102 18367 20154
rect 18367 20102 18377 20154
rect 18401 20102 18431 20154
rect 18431 20102 18443 20154
rect 18443 20102 18457 20154
rect 18481 20102 18495 20154
rect 18495 20102 18507 20154
rect 18507 20102 18537 20154
rect 18561 20102 18571 20154
rect 18571 20102 18617 20154
rect 18321 20100 18377 20102
rect 18401 20100 18457 20102
rect 18481 20100 18537 20102
rect 18561 20100 18617 20102
rect 18321 19066 18377 19068
rect 18401 19066 18457 19068
rect 18481 19066 18537 19068
rect 18561 19066 18617 19068
rect 18321 19014 18367 19066
rect 18367 19014 18377 19066
rect 18401 19014 18431 19066
rect 18431 19014 18443 19066
rect 18443 19014 18457 19066
rect 18481 19014 18495 19066
rect 18495 19014 18507 19066
rect 18507 19014 18537 19066
rect 18561 19014 18571 19066
rect 18571 19014 18617 19066
rect 18321 19012 18377 19014
rect 18401 19012 18457 19014
rect 18481 19012 18537 19014
rect 18561 19012 18617 19014
rect 18321 17978 18377 17980
rect 18401 17978 18457 17980
rect 18481 17978 18537 17980
rect 18561 17978 18617 17980
rect 18321 17926 18367 17978
rect 18367 17926 18377 17978
rect 18401 17926 18431 17978
rect 18431 17926 18443 17978
rect 18443 17926 18457 17978
rect 18481 17926 18495 17978
rect 18495 17926 18507 17978
rect 18507 17926 18537 17978
rect 18561 17926 18571 17978
rect 18571 17926 18617 17978
rect 18321 17924 18377 17926
rect 18401 17924 18457 17926
rect 18481 17924 18537 17926
rect 18561 17924 18617 17926
rect 18321 16890 18377 16892
rect 18401 16890 18457 16892
rect 18481 16890 18537 16892
rect 18561 16890 18617 16892
rect 18321 16838 18367 16890
rect 18367 16838 18377 16890
rect 18401 16838 18431 16890
rect 18431 16838 18443 16890
rect 18443 16838 18457 16890
rect 18481 16838 18495 16890
rect 18495 16838 18507 16890
rect 18507 16838 18537 16890
rect 18561 16838 18571 16890
rect 18571 16838 18617 16890
rect 18321 16836 18377 16838
rect 18401 16836 18457 16838
rect 18481 16836 18537 16838
rect 18561 16836 18617 16838
rect 18321 15802 18377 15804
rect 18401 15802 18457 15804
rect 18481 15802 18537 15804
rect 18561 15802 18617 15804
rect 18321 15750 18367 15802
rect 18367 15750 18377 15802
rect 18401 15750 18431 15802
rect 18431 15750 18443 15802
rect 18443 15750 18457 15802
rect 18481 15750 18495 15802
rect 18495 15750 18507 15802
rect 18507 15750 18537 15802
rect 18561 15750 18571 15802
rect 18571 15750 18617 15802
rect 18321 15748 18377 15750
rect 18401 15748 18457 15750
rect 18481 15748 18537 15750
rect 18561 15748 18617 15750
rect 18321 14714 18377 14716
rect 18401 14714 18457 14716
rect 18481 14714 18537 14716
rect 18561 14714 18617 14716
rect 18321 14662 18367 14714
rect 18367 14662 18377 14714
rect 18401 14662 18431 14714
rect 18431 14662 18443 14714
rect 18443 14662 18457 14714
rect 18481 14662 18495 14714
rect 18495 14662 18507 14714
rect 18507 14662 18537 14714
rect 18561 14662 18571 14714
rect 18571 14662 18617 14714
rect 18321 14660 18377 14662
rect 18401 14660 18457 14662
rect 18481 14660 18537 14662
rect 18561 14660 18617 14662
rect 18321 13626 18377 13628
rect 18401 13626 18457 13628
rect 18481 13626 18537 13628
rect 18561 13626 18617 13628
rect 18321 13574 18367 13626
rect 18367 13574 18377 13626
rect 18401 13574 18431 13626
rect 18431 13574 18443 13626
rect 18443 13574 18457 13626
rect 18481 13574 18495 13626
rect 18495 13574 18507 13626
rect 18507 13574 18537 13626
rect 18561 13574 18571 13626
rect 18571 13574 18617 13626
rect 18321 13572 18377 13574
rect 18401 13572 18457 13574
rect 18481 13572 18537 13574
rect 18561 13572 18617 13574
rect 18321 12538 18377 12540
rect 18401 12538 18457 12540
rect 18481 12538 18537 12540
rect 18561 12538 18617 12540
rect 18321 12486 18367 12538
rect 18367 12486 18377 12538
rect 18401 12486 18431 12538
rect 18431 12486 18443 12538
rect 18443 12486 18457 12538
rect 18481 12486 18495 12538
rect 18495 12486 18507 12538
rect 18507 12486 18537 12538
rect 18561 12486 18571 12538
rect 18571 12486 18617 12538
rect 18321 12484 18377 12486
rect 18401 12484 18457 12486
rect 18481 12484 18537 12486
rect 18561 12484 18617 12486
rect 18878 11892 18934 11928
rect 18878 11872 18880 11892
rect 18880 11872 18932 11892
rect 18932 11872 18934 11892
rect 18321 11450 18377 11452
rect 18401 11450 18457 11452
rect 18481 11450 18537 11452
rect 18561 11450 18617 11452
rect 18321 11398 18367 11450
rect 18367 11398 18377 11450
rect 18401 11398 18431 11450
rect 18431 11398 18443 11450
rect 18443 11398 18457 11450
rect 18481 11398 18495 11450
rect 18495 11398 18507 11450
rect 18507 11398 18537 11450
rect 18561 11398 18571 11450
rect 18571 11398 18617 11450
rect 18321 11396 18377 11398
rect 18401 11396 18457 11398
rect 18481 11396 18537 11398
rect 18561 11396 18617 11398
rect 21794 37018 21850 37020
rect 21874 37018 21930 37020
rect 21954 37018 22010 37020
rect 22034 37018 22090 37020
rect 21794 36966 21840 37018
rect 21840 36966 21850 37018
rect 21874 36966 21904 37018
rect 21904 36966 21916 37018
rect 21916 36966 21930 37018
rect 21954 36966 21968 37018
rect 21968 36966 21980 37018
rect 21980 36966 22010 37018
rect 22034 36966 22044 37018
rect 22044 36966 22090 37018
rect 21794 36964 21850 36966
rect 21874 36964 21930 36966
rect 21954 36964 22010 36966
rect 22034 36964 22090 36966
rect 21794 35930 21850 35932
rect 21874 35930 21930 35932
rect 21954 35930 22010 35932
rect 22034 35930 22090 35932
rect 21794 35878 21840 35930
rect 21840 35878 21850 35930
rect 21874 35878 21904 35930
rect 21904 35878 21916 35930
rect 21916 35878 21930 35930
rect 21954 35878 21968 35930
rect 21968 35878 21980 35930
rect 21980 35878 22010 35930
rect 22034 35878 22044 35930
rect 22044 35878 22090 35930
rect 21794 35876 21850 35878
rect 21874 35876 21930 35878
rect 21954 35876 22010 35878
rect 22034 35876 22090 35878
rect 26146 46960 26202 47016
rect 26054 46280 26110 46336
rect 25267 46266 25323 46268
rect 25347 46266 25403 46268
rect 25427 46266 25483 46268
rect 25507 46266 25563 46268
rect 25267 46214 25313 46266
rect 25313 46214 25323 46266
rect 25347 46214 25377 46266
rect 25377 46214 25389 46266
rect 25389 46214 25403 46266
rect 25427 46214 25441 46266
rect 25441 46214 25453 46266
rect 25453 46214 25483 46266
rect 25507 46214 25517 46266
rect 25517 46214 25563 46266
rect 25267 46212 25323 46214
rect 25347 46212 25403 46214
rect 25427 46212 25483 46214
rect 25507 46212 25563 46214
rect 25267 45178 25323 45180
rect 25347 45178 25403 45180
rect 25427 45178 25483 45180
rect 25507 45178 25563 45180
rect 25267 45126 25313 45178
rect 25313 45126 25323 45178
rect 25347 45126 25377 45178
rect 25377 45126 25389 45178
rect 25389 45126 25403 45178
rect 25427 45126 25441 45178
rect 25441 45126 25453 45178
rect 25453 45126 25483 45178
rect 25507 45126 25517 45178
rect 25517 45126 25563 45178
rect 25267 45124 25323 45126
rect 25347 45124 25403 45126
rect 25427 45124 25483 45126
rect 25507 45124 25563 45126
rect 25267 44090 25323 44092
rect 25347 44090 25403 44092
rect 25427 44090 25483 44092
rect 25507 44090 25563 44092
rect 25267 44038 25313 44090
rect 25313 44038 25323 44090
rect 25347 44038 25377 44090
rect 25377 44038 25389 44090
rect 25389 44038 25403 44090
rect 25427 44038 25441 44090
rect 25441 44038 25453 44090
rect 25453 44038 25483 44090
rect 25507 44038 25517 44090
rect 25517 44038 25563 44090
rect 25267 44036 25323 44038
rect 25347 44036 25403 44038
rect 25427 44036 25483 44038
rect 25507 44036 25563 44038
rect 25267 43002 25323 43004
rect 25347 43002 25403 43004
rect 25427 43002 25483 43004
rect 25507 43002 25563 43004
rect 25267 42950 25313 43002
rect 25313 42950 25323 43002
rect 25347 42950 25377 43002
rect 25377 42950 25389 43002
rect 25389 42950 25403 43002
rect 25427 42950 25441 43002
rect 25441 42950 25453 43002
rect 25453 42950 25483 43002
rect 25507 42950 25517 43002
rect 25517 42950 25563 43002
rect 25267 42948 25323 42950
rect 25347 42948 25403 42950
rect 25427 42948 25483 42950
rect 25507 42948 25563 42950
rect 25267 41914 25323 41916
rect 25347 41914 25403 41916
rect 25427 41914 25483 41916
rect 25507 41914 25563 41916
rect 25267 41862 25313 41914
rect 25313 41862 25323 41914
rect 25347 41862 25377 41914
rect 25377 41862 25389 41914
rect 25389 41862 25403 41914
rect 25427 41862 25441 41914
rect 25441 41862 25453 41914
rect 25453 41862 25483 41914
rect 25507 41862 25517 41914
rect 25517 41862 25563 41914
rect 25267 41860 25323 41862
rect 25347 41860 25403 41862
rect 25427 41860 25483 41862
rect 25507 41860 25563 41862
rect 25267 40826 25323 40828
rect 25347 40826 25403 40828
rect 25427 40826 25483 40828
rect 25507 40826 25563 40828
rect 25267 40774 25313 40826
rect 25313 40774 25323 40826
rect 25347 40774 25377 40826
rect 25377 40774 25389 40826
rect 25389 40774 25403 40826
rect 25427 40774 25441 40826
rect 25441 40774 25453 40826
rect 25453 40774 25483 40826
rect 25507 40774 25517 40826
rect 25517 40774 25563 40826
rect 25267 40772 25323 40774
rect 25347 40772 25403 40774
rect 25427 40772 25483 40774
rect 25507 40772 25563 40774
rect 25267 39738 25323 39740
rect 25347 39738 25403 39740
rect 25427 39738 25483 39740
rect 25507 39738 25563 39740
rect 25267 39686 25313 39738
rect 25313 39686 25323 39738
rect 25347 39686 25377 39738
rect 25377 39686 25389 39738
rect 25389 39686 25403 39738
rect 25427 39686 25441 39738
rect 25441 39686 25453 39738
rect 25453 39686 25483 39738
rect 25507 39686 25517 39738
rect 25517 39686 25563 39738
rect 25267 39684 25323 39686
rect 25347 39684 25403 39686
rect 25427 39684 25483 39686
rect 25507 39684 25563 39686
rect 25267 38650 25323 38652
rect 25347 38650 25403 38652
rect 25427 38650 25483 38652
rect 25507 38650 25563 38652
rect 25267 38598 25313 38650
rect 25313 38598 25323 38650
rect 25347 38598 25377 38650
rect 25377 38598 25389 38650
rect 25389 38598 25403 38650
rect 25427 38598 25441 38650
rect 25441 38598 25453 38650
rect 25453 38598 25483 38650
rect 25507 38598 25517 38650
rect 25517 38598 25563 38650
rect 25267 38596 25323 38598
rect 25347 38596 25403 38598
rect 25427 38596 25483 38598
rect 25507 38596 25563 38598
rect 25267 37562 25323 37564
rect 25347 37562 25403 37564
rect 25427 37562 25483 37564
rect 25507 37562 25563 37564
rect 25267 37510 25313 37562
rect 25313 37510 25323 37562
rect 25347 37510 25377 37562
rect 25377 37510 25389 37562
rect 25389 37510 25403 37562
rect 25427 37510 25441 37562
rect 25441 37510 25453 37562
rect 25453 37510 25483 37562
rect 25507 37510 25517 37562
rect 25517 37510 25563 37562
rect 25267 37508 25323 37510
rect 25347 37508 25403 37510
rect 25427 37508 25483 37510
rect 25507 37508 25563 37510
rect 21794 34842 21850 34844
rect 21874 34842 21930 34844
rect 21954 34842 22010 34844
rect 22034 34842 22090 34844
rect 21794 34790 21840 34842
rect 21840 34790 21850 34842
rect 21874 34790 21904 34842
rect 21904 34790 21916 34842
rect 21916 34790 21930 34842
rect 21954 34790 21968 34842
rect 21968 34790 21980 34842
rect 21980 34790 22010 34842
rect 22034 34790 22044 34842
rect 22044 34790 22090 34842
rect 21794 34788 21850 34790
rect 21874 34788 21930 34790
rect 21954 34788 22010 34790
rect 22034 34788 22090 34790
rect 21794 33754 21850 33756
rect 21874 33754 21930 33756
rect 21954 33754 22010 33756
rect 22034 33754 22090 33756
rect 21794 33702 21840 33754
rect 21840 33702 21850 33754
rect 21874 33702 21904 33754
rect 21904 33702 21916 33754
rect 21916 33702 21930 33754
rect 21954 33702 21968 33754
rect 21968 33702 21980 33754
rect 21980 33702 22010 33754
rect 22034 33702 22044 33754
rect 22044 33702 22090 33754
rect 21794 33700 21850 33702
rect 21874 33700 21930 33702
rect 21954 33700 22010 33702
rect 22034 33700 22090 33702
rect 21794 32666 21850 32668
rect 21874 32666 21930 32668
rect 21954 32666 22010 32668
rect 22034 32666 22090 32668
rect 21794 32614 21840 32666
rect 21840 32614 21850 32666
rect 21874 32614 21904 32666
rect 21904 32614 21916 32666
rect 21916 32614 21930 32666
rect 21954 32614 21968 32666
rect 21968 32614 21980 32666
rect 21980 32614 22010 32666
rect 22034 32614 22044 32666
rect 22044 32614 22090 32666
rect 21794 32612 21850 32614
rect 21874 32612 21930 32614
rect 21954 32612 22010 32614
rect 22034 32612 22090 32614
rect 21794 31578 21850 31580
rect 21874 31578 21930 31580
rect 21954 31578 22010 31580
rect 22034 31578 22090 31580
rect 21794 31526 21840 31578
rect 21840 31526 21850 31578
rect 21874 31526 21904 31578
rect 21904 31526 21916 31578
rect 21916 31526 21930 31578
rect 21954 31526 21968 31578
rect 21968 31526 21980 31578
rect 21980 31526 22010 31578
rect 22034 31526 22044 31578
rect 22044 31526 22090 31578
rect 21794 31524 21850 31526
rect 21874 31524 21930 31526
rect 21954 31524 22010 31526
rect 22034 31524 22090 31526
rect 21794 30490 21850 30492
rect 21874 30490 21930 30492
rect 21954 30490 22010 30492
rect 22034 30490 22090 30492
rect 21794 30438 21840 30490
rect 21840 30438 21850 30490
rect 21874 30438 21904 30490
rect 21904 30438 21916 30490
rect 21916 30438 21930 30490
rect 21954 30438 21968 30490
rect 21968 30438 21980 30490
rect 21980 30438 22010 30490
rect 22034 30438 22044 30490
rect 22044 30438 22090 30490
rect 21794 30436 21850 30438
rect 21874 30436 21930 30438
rect 21954 30436 22010 30438
rect 22034 30436 22090 30438
rect 21794 29402 21850 29404
rect 21874 29402 21930 29404
rect 21954 29402 22010 29404
rect 22034 29402 22090 29404
rect 21794 29350 21840 29402
rect 21840 29350 21850 29402
rect 21874 29350 21904 29402
rect 21904 29350 21916 29402
rect 21916 29350 21930 29402
rect 21954 29350 21968 29402
rect 21968 29350 21980 29402
rect 21980 29350 22010 29402
rect 22034 29350 22044 29402
rect 22044 29350 22090 29402
rect 21794 29348 21850 29350
rect 21874 29348 21930 29350
rect 21954 29348 22010 29350
rect 22034 29348 22090 29350
rect 21794 28314 21850 28316
rect 21874 28314 21930 28316
rect 21954 28314 22010 28316
rect 22034 28314 22090 28316
rect 21794 28262 21840 28314
rect 21840 28262 21850 28314
rect 21874 28262 21904 28314
rect 21904 28262 21916 28314
rect 21916 28262 21930 28314
rect 21954 28262 21968 28314
rect 21968 28262 21980 28314
rect 21980 28262 22010 28314
rect 22034 28262 22044 28314
rect 22044 28262 22090 28314
rect 21794 28260 21850 28262
rect 21874 28260 21930 28262
rect 21954 28260 22010 28262
rect 22034 28260 22090 28262
rect 21794 27226 21850 27228
rect 21874 27226 21930 27228
rect 21954 27226 22010 27228
rect 22034 27226 22090 27228
rect 21794 27174 21840 27226
rect 21840 27174 21850 27226
rect 21874 27174 21904 27226
rect 21904 27174 21916 27226
rect 21916 27174 21930 27226
rect 21954 27174 21968 27226
rect 21968 27174 21980 27226
rect 21980 27174 22010 27226
rect 22034 27174 22044 27226
rect 22044 27174 22090 27226
rect 21794 27172 21850 27174
rect 21874 27172 21930 27174
rect 21954 27172 22010 27174
rect 22034 27172 22090 27174
rect 21794 26138 21850 26140
rect 21874 26138 21930 26140
rect 21954 26138 22010 26140
rect 22034 26138 22090 26140
rect 21794 26086 21840 26138
rect 21840 26086 21850 26138
rect 21874 26086 21904 26138
rect 21904 26086 21916 26138
rect 21916 26086 21930 26138
rect 21954 26086 21968 26138
rect 21968 26086 21980 26138
rect 21980 26086 22010 26138
rect 22034 26086 22044 26138
rect 22044 26086 22090 26138
rect 21794 26084 21850 26086
rect 21874 26084 21930 26086
rect 21954 26084 22010 26086
rect 22034 26084 22090 26086
rect 21794 25050 21850 25052
rect 21874 25050 21930 25052
rect 21954 25050 22010 25052
rect 22034 25050 22090 25052
rect 21794 24998 21840 25050
rect 21840 24998 21850 25050
rect 21874 24998 21904 25050
rect 21904 24998 21916 25050
rect 21916 24998 21930 25050
rect 21954 24998 21968 25050
rect 21968 24998 21980 25050
rect 21980 24998 22010 25050
rect 22034 24998 22044 25050
rect 22044 24998 22090 25050
rect 21794 24996 21850 24998
rect 21874 24996 21930 24998
rect 21954 24996 22010 24998
rect 22034 24996 22090 24998
rect 21794 23962 21850 23964
rect 21874 23962 21930 23964
rect 21954 23962 22010 23964
rect 22034 23962 22090 23964
rect 21794 23910 21840 23962
rect 21840 23910 21850 23962
rect 21874 23910 21904 23962
rect 21904 23910 21916 23962
rect 21916 23910 21930 23962
rect 21954 23910 21968 23962
rect 21968 23910 21980 23962
rect 21980 23910 22010 23962
rect 22034 23910 22044 23962
rect 22044 23910 22090 23962
rect 21794 23908 21850 23910
rect 21874 23908 21930 23910
rect 21954 23908 22010 23910
rect 22034 23908 22090 23910
rect 21794 22874 21850 22876
rect 21874 22874 21930 22876
rect 21954 22874 22010 22876
rect 22034 22874 22090 22876
rect 21794 22822 21840 22874
rect 21840 22822 21850 22874
rect 21874 22822 21904 22874
rect 21904 22822 21916 22874
rect 21916 22822 21930 22874
rect 21954 22822 21968 22874
rect 21968 22822 21980 22874
rect 21980 22822 22010 22874
rect 22034 22822 22044 22874
rect 22044 22822 22090 22874
rect 21794 22820 21850 22822
rect 21874 22820 21930 22822
rect 21954 22820 22010 22822
rect 22034 22820 22090 22822
rect 21794 21786 21850 21788
rect 21874 21786 21930 21788
rect 21954 21786 22010 21788
rect 22034 21786 22090 21788
rect 21794 21734 21840 21786
rect 21840 21734 21850 21786
rect 21874 21734 21904 21786
rect 21904 21734 21916 21786
rect 21916 21734 21930 21786
rect 21954 21734 21968 21786
rect 21968 21734 21980 21786
rect 21980 21734 22010 21786
rect 22034 21734 22044 21786
rect 22044 21734 22090 21786
rect 21794 21732 21850 21734
rect 21874 21732 21930 21734
rect 21954 21732 22010 21734
rect 22034 21732 22090 21734
rect 18321 10362 18377 10364
rect 18401 10362 18457 10364
rect 18481 10362 18537 10364
rect 18561 10362 18617 10364
rect 18321 10310 18367 10362
rect 18367 10310 18377 10362
rect 18401 10310 18431 10362
rect 18431 10310 18443 10362
rect 18443 10310 18457 10362
rect 18481 10310 18495 10362
rect 18495 10310 18507 10362
rect 18507 10310 18537 10362
rect 18561 10310 18571 10362
rect 18571 10310 18617 10362
rect 18321 10308 18377 10310
rect 18401 10308 18457 10310
rect 18481 10308 18537 10310
rect 18561 10308 18617 10310
rect 21794 20698 21850 20700
rect 21874 20698 21930 20700
rect 21954 20698 22010 20700
rect 22034 20698 22090 20700
rect 21794 20646 21840 20698
rect 21840 20646 21850 20698
rect 21874 20646 21904 20698
rect 21904 20646 21916 20698
rect 21916 20646 21930 20698
rect 21954 20646 21968 20698
rect 21968 20646 21980 20698
rect 21980 20646 22010 20698
rect 22034 20646 22044 20698
rect 22044 20646 22090 20698
rect 21794 20644 21850 20646
rect 21874 20644 21930 20646
rect 21954 20644 22010 20646
rect 22034 20644 22090 20646
rect 21794 19610 21850 19612
rect 21874 19610 21930 19612
rect 21954 19610 22010 19612
rect 22034 19610 22090 19612
rect 21794 19558 21840 19610
rect 21840 19558 21850 19610
rect 21874 19558 21904 19610
rect 21904 19558 21916 19610
rect 21916 19558 21930 19610
rect 21954 19558 21968 19610
rect 21968 19558 21980 19610
rect 21980 19558 22010 19610
rect 22034 19558 22044 19610
rect 22044 19558 22090 19610
rect 21794 19556 21850 19558
rect 21874 19556 21930 19558
rect 21954 19556 22010 19558
rect 22034 19556 22090 19558
rect 21794 18522 21850 18524
rect 21874 18522 21930 18524
rect 21954 18522 22010 18524
rect 22034 18522 22090 18524
rect 21794 18470 21840 18522
rect 21840 18470 21850 18522
rect 21874 18470 21904 18522
rect 21904 18470 21916 18522
rect 21916 18470 21930 18522
rect 21954 18470 21968 18522
rect 21968 18470 21980 18522
rect 21980 18470 22010 18522
rect 22034 18470 22044 18522
rect 22044 18470 22090 18522
rect 21794 18468 21850 18470
rect 21874 18468 21930 18470
rect 21954 18468 22010 18470
rect 22034 18468 22090 18470
rect 21794 17434 21850 17436
rect 21874 17434 21930 17436
rect 21954 17434 22010 17436
rect 22034 17434 22090 17436
rect 21794 17382 21840 17434
rect 21840 17382 21850 17434
rect 21874 17382 21904 17434
rect 21904 17382 21916 17434
rect 21916 17382 21930 17434
rect 21954 17382 21968 17434
rect 21968 17382 21980 17434
rect 21980 17382 22010 17434
rect 22034 17382 22044 17434
rect 22044 17382 22090 17434
rect 21794 17380 21850 17382
rect 21874 17380 21930 17382
rect 21954 17380 22010 17382
rect 22034 17380 22090 17382
rect 21794 16346 21850 16348
rect 21874 16346 21930 16348
rect 21954 16346 22010 16348
rect 22034 16346 22090 16348
rect 21794 16294 21840 16346
rect 21840 16294 21850 16346
rect 21874 16294 21904 16346
rect 21904 16294 21916 16346
rect 21916 16294 21930 16346
rect 21954 16294 21968 16346
rect 21968 16294 21980 16346
rect 21980 16294 22010 16346
rect 22034 16294 22044 16346
rect 22044 16294 22090 16346
rect 21794 16292 21850 16294
rect 21874 16292 21930 16294
rect 21954 16292 22010 16294
rect 22034 16292 22090 16294
rect 21794 15258 21850 15260
rect 21874 15258 21930 15260
rect 21954 15258 22010 15260
rect 22034 15258 22090 15260
rect 21794 15206 21840 15258
rect 21840 15206 21850 15258
rect 21874 15206 21904 15258
rect 21904 15206 21916 15258
rect 21916 15206 21930 15258
rect 21954 15206 21968 15258
rect 21968 15206 21980 15258
rect 21980 15206 22010 15258
rect 22034 15206 22044 15258
rect 22044 15206 22090 15258
rect 21794 15204 21850 15206
rect 21874 15204 21930 15206
rect 21954 15204 22010 15206
rect 22034 15204 22090 15206
rect 21794 14170 21850 14172
rect 21874 14170 21930 14172
rect 21954 14170 22010 14172
rect 22034 14170 22090 14172
rect 21794 14118 21840 14170
rect 21840 14118 21850 14170
rect 21874 14118 21904 14170
rect 21904 14118 21916 14170
rect 21916 14118 21930 14170
rect 21954 14118 21968 14170
rect 21968 14118 21980 14170
rect 21980 14118 22010 14170
rect 22034 14118 22044 14170
rect 22044 14118 22090 14170
rect 21794 14116 21850 14118
rect 21874 14116 21930 14118
rect 21954 14116 22010 14118
rect 22034 14116 22090 14118
rect 21794 13082 21850 13084
rect 21874 13082 21930 13084
rect 21954 13082 22010 13084
rect 22034 13082 22090 13084
rect 21794 13030 21840 13082
rect 21840 13030 21850 13082
rect 21874 13030 21904 13082
rect 21904 13030 21916 13082
rect 21916 13030 21930 13082
rect 21954 13030 21968 13082
rect 21968 13030 21980 13082
rect 21980 13030 22010 13082
rect 22034 13030 22044 13082
rect 22044 13030 22090 13082
rect 21794 13028 21850 13030
rect 21874 13028 21930 13030
rect 21954 13028 22010 13030
rect 22034 13028 22090 13030
rect 25267 36474 25323 36476
rect 25347 36474 25403 36476
rect 25427 36474 25483 36476
rect 25507 36474 25563 36476
rect 25267 36422 25313 36474
rect 25313 36422 25323 36474
rect 25347 36422 25377 36474
rect 25377 36422 25389 36474
rect 25389 36422 25403 36474
rect 25427 36422 25441 36474
rect 25441 36422 25453 36474
rect 25453 36422 25483 36474
rect 25507 36422 25517 36474
rect 25517 36422 25563 36474
rect 25267 36420 25323 36422
rect 25347 36420 25403 36422
rect 25427 36420 25483 36422
rect 25507 36420 25563 36422
rect 25267 35386 25323 35388
rect 25347 35386 25403 35388
rect 25427 35386 25483 35388
rect 25507 35386 25563 35388
rect 25267 35334 25313 35386
rect 25313 35334 25323 35386
rect 25347 35334 25377 35386
rect 25377 35334 25389 35386
rect 25389 35334 25403 35386
rect 25427 35334 25441 35386
rect 25441 35334 25453 35386
rect 25453 35334 25483 35386
rect 25507 35334 25517 35386
rect 25517 35334 25563 35386
rect 25267 35332 25323 35334
rect 25347 35332 25403 35334
rect 25427 35332 25483 35334
rect 25507 35332 25563 35334
rect 26054 42880 26110 42936
rect 26146 41520 26202 41576
rect 26606 38392 26662 38448
rect 26146 36080 26202 36136
rect 25267 34298 25323 34300
rect 25347 34298 25403 34300
rect 25427 34298 25483 34300
rect 25507 34298 25563 34300
rect 25267 34246 25313 34298
rect 25313 34246 25323 34298
rect 25347 34246 25377 34298
rect 25377 34246 25389 34298
rect 25389 34246 25403 34298
rect 25427 34246 25441 34298
rect 25441 34246 25453 34298
rect 25453 34246 25483 34298
rect 25507 34246 25517 34298
rect 25517 34246 25563 34298
rect 25267 34244 25323 34246
rect 25347 34244 25403 34246
rect 25427 34244 25483 34246
rect 25507 34244 25563 34246
rect 25267 33210 25323 33212
rect 25347 33210 25403 33212
rect 25427 33210 25483 33212
rect 25507 33210 25563 33212
rect 25267 33158 25313 33210
rect 25313 33158 25323 33210
rect 25347 33158 25377 33210
rect 25377 33158 25389 33210
rect 25389 33158 25403 33210
rect 25427 33158 25441 33210
rect 25441 33158 25453 33210
rect 25453 33158 25483 33210
rect 25507 33158 25517 33210
rect 25517 33158 25563 33210
rect 25267 33156 25323 33158
rect 25347 33156 25403 33158
rect 25427 33156 25483 33158
rect 25507 33156 25563 33158
rect 25267 32122 25323 32124
rect 25347 32122 25403 32124
rect 25427 32122 25483 32124
rect 25507 32122 25563 32124
rect 25267 32070 25313 32122
rect 25313 32070 25323 32122
rect 25347 32070 25377 32122
rect 25377 32070 25389 32122
rect 25389 32070 25403 32122
rect 25427 32070 25441 32122
rect 25441 32070 25453 32122
rect 25453 32070 25483 32122
rect 25507 32070 25517 32122
rect 25517 32070 25563 32122
rect 25267 32068 25323 32070
rect 25347 32068 25403 32070
rect 25427 32068 25483 32070
rect 25507 32068 25563 32070
rect 25267 31034 25323 31036
rect 25347 31034 25403 31036
rect 25427 31034 25483 31036
rect 25507 31034 25563 31036
rect 25267 30982 25313 31034
rect 25313 30982 25323 31034
rect 25347 30982 25377 31034
rect 25377 30982 25389 31034
rect 25389 30982 25403 31034
rect 25427 30982 25441 31034
rect 25441 30982 25453 31034
rect 25453 30982 25483 31034
rect 25507 30982 25517 31034
rect 25517 30982 25563 31034
rect 25267 30980 25323 30982
rect 25347 30980 25403 30982
rect 25427 30980 25483 30982
rect 25507 30980 25563 30982
rect 25267 29946 25323 29948
rect 25347 29946 25403 29948
rect 25427 29946 25483 29948
rect 25507 29946 25563 29948
rect 25267 29894 25313 29946
rect 25313 29894 25323 29946
rect 25347 29894 25377 29946
rect 25377 29894 25389 29946
rect 25389 29894 25403 29946
rect 25427 29894 25441 29946
rect 25441 29894 25453 29946
rect 25453 29894 25483 29946
rect 25507 29894 25517 29946
rect 25517 29894 25563 29946
rect 25267 29892 25323 29894
rect 25347 29892 25403 29894
rect 25427 29892 25483 29894
rect 25507 29892 25563 29894
rect 26146 31320 26202 31376
rect 24766 29008 24822 29064
rect 25267 28858 25323 28860
rect 25347 28858 25403 28860
rect 25427 28858 25483 28860
rect 25507 28858 25563 28860
rect 25267 28806 25313 28858
rect 25313 28806 25323 28858
rect 25347 28806 25377 28858
rect 25377 28806 25389 28858
rect 25389 28806 25403 28858
rect 25427 28806 25441 28858
rect 25441 28806 25453 28858
rect 25453 28806 25483 28858
rect 25507 28806 25517 28858
rect 25517 28806 25563 28858
rect 25267 28804 25323 28806
rect 25347 28804 25403 28806
rect 25427 28804 25483 28806
rect 25507 28804 25563 28806
rect 25267 27770 25323 27772
rect 25347 27770 25403 27772
rect 25427 27770 25483 27772
rect 25507 27770 25563 27772
rect 25267 27718 25313 27770
rect 25313 27718 25323 27770
rect 25347 27718 25377 27770
rect 25377 27718 25389 27770
rect 25389 27718 25403 27770
rect 25427 27718 25441 27770
rect 25441 27718 25453 27770
rect 25453 27718 25483 27770
rect 25507 27718 25517 27770
rect 25517 27718 25563 27770
rect 25267 27716 25323 27718
rect 25347 27716 25403 27718
rect 25427 27716 25483 27718
rect 25507 27716 25563 27718
rect 25267 26682 25323 26684
rect 25347 26682 25403 26684
rect 25427 26682 25483 26684
rect 25507 26682 25563 26684
rect 25267 26630 25313 26682
rect 25313 26630 25323 26682
rect 25347 26630 25377 26682
rect 25377 26630 25389 26682
rect 25389 26630 25403 26682
rect 25427 26630 25441 26682
rect 25441 26630 25453 26682
rect 25453 26630 25483 26682
rect 25507 26630 25517 26682
rect 25517 26630 25563 26682
rect 25267 26628 25323 26630
rect 25347 26628 25403 26630
rect 25427 26628 25483 26630
rect 25507 26628 25563 26630
rect 25267 25594 25323 25596
rect 25347 25594 25403 25596
rect 25427 25594 25483 25596
rect 25507 25594 25563 25596
rect 25267 25542 25313 25594
rect 25313 25542 25323 25594
rect 25347 25542 25377 25594
rect 25377 25542 25389 25594
rect 25389 25542 25403 25594
rect 25427 25542 25441 25594
rect 25441 25542 25453 25594
rect 25453 25542 25483 25594
rect 25507 25542 25517 25594
rect 25517 25542 25563 25594
rect 25267 25540 25323 25542
rect 25347 25540 25403 25542
rect 25427 25540 25483 25542
rect 25507 25540 25563 25542
rect 25267 24506 25323 24508
rect 25347 24506 25403 24508
rect 25427 24506 25483 24508
rect 25507 24506 25563 24508
rect 25267 24454 25313 24506
rect 25313 24454 25323 24506
rect 25347 24454 25377 24506
rect 25377 24454 25389 24506
rect 25389 24454 25403 24506
rect 25427 24454 25441 24506
rect 25441 24454 25453 24506
rect 25453 24454 25483 24506
rect 25507 24454 25517 24506
rect 25517 24454 25563 24506
rect 25267 24452 25323 24454
rect 25347 24452 25403 24454
rect 25427 24452 25483 24454
rect 25507 24452 25563 24454
rect 25267 23418 25323 23420
rect 25347 23418 25403 23420
rect 25427 23418 25483 23420
rect 25507 23418 25563 23420
rect 25267 23366 25313 23418
rect 25313 23366 25323 23418
rect 25347 23366 25377 23418
rect 25377 23366 25389 23418
rect 25389 23366 25403 23418
rect 25427 23366 25441 23418
rect 25441 23366 25453 23418
rect 25453 23366 25483 23418
rect 25507 23366 25517 23418
rect 25517 23366 25563 23418
rect 25267 23364 25323 23366
rect 25347 23364 25403 23366
rect 25427 23364 25483 23366
rect 25507 23364 25563 23366
rect 25267 22330 25323 22332
rect 25347 22330 25403 22332
rect 25427 22330 25483 22332
rect 25507 22330 25563 22332
rect 25267 22278 25313 22330
rect 25313 22278 25323 22330
rect 25347 22278 25377 22330
rect 25377 22278 25389 22330
rect 25389 22278 25403 22330
rect 25427 22278 25441 22330
rect 25441 22278 25453 22330
rect 25453 22278 25483 22330
rect 25507 22278 25517 22330
rect 25517 22278 25563 22330
rect 25267 22276 25323 22278
rect 25347 22276 25403 22278
rect 25427 22276 25483 22278
rect 25507 22276 25563 22278
rect 25267 21242 25323 21244
rect 25347 21242 25403 21244
rect 25427 21242 25483 21244
rect 25507 21242 25563 21244
rect 25267 21190 25313 21242
rect 25313 21190 25323 21242
rect 25347 21190 25377 21242
rect 25377 21190 25389 21242
rect 25389 21190 25403 21242
rect 25427 21190 25441 21242
rect 25441 21190 25453 21242
rect 25453 21190 25483 21242
rect 25507 21190 25517 21242
rect 25517 21190 25563 21242
rect 25267 21188 25323 21190
rect 25347 21188 25403 21190
rect 25427 21188 25483 21190
rect 25507 21188 25563 21190
rect 26146 21392 26202 21448
rect 25267 20154 25323 20156
rect 25347 20154 25403 20156
rect 25427 20154 25483 20156
rect 25507 20154 25563 20156
rect 25267 20102 25313 20154
rect 25313 20102 25323 20154
rect 25347 20102 25377 20154
rect 25377 20102 25389 20154
rect 25389 20102 25403 20154
rect 25427 20102 25441 20154
rect 25441 20102 25453 20154
rect 25453 20102 25483 20154
rect 25507 20102 25517 20154
rect 25517 20102 25563 20154
rect 25267 20100 25323 20102
rect 25347 20100 25403 20102
rect 25427 20100 25483 20102
rect 25507 20100 25563 20102
rect 25267 19066 25323 19068
rect 25347 19066 25403 19068
rect 25427 19066 25483 19068
rect 25507 19066 25563 19068
rect 25267 19014 25313 19066
rect 25313 19014 25323 19066
rect 25347 19014 25377 19066
rect 25377 19014 25389 19066
rect 25389 19014 25403 19066
rect 25427 19014 25441 19066
rect 25441 19014 25453 19066
rect 25453 19014 25483 19066
rect 25507 19014 25517 19066
rect 25517 19014 25563 19066
rect 25267 19012 25323 19014
rect 25347 19012 25403 19014
rect 25427 19012 25483 19014
rect 25507 19012 25563 19014
rect 26606 29960 26662 30016
rect 27434 42200 27490 42256
rect 28630 47640 28686 47696
rect 28354 44940 28410 44976
rect 28354 44920 28356 44940
rect 28356 44920 28408 44940
rect 28408 44920 28410 44940
rect 27342 36780 27398 36816
rect 27342 36760 27344 36780
rect 27344 36760 27396 36780
rect 27396 36760 27398 36780
rect 27526 40840 27582 40896
rect 28740 46810 28796 46812
rect 28820 46810 28876 46812
rect 28900 46810 28956 46812
rect 28980 46810 29036 46812
rect 28740 46758 28786 46810
rect 28786 46758 28796 46810
rect 28820 46758 28850 46810
rect 28850 46758 28862 46810
rect 28862 46758 28876 46810
rect 28900 46758 28914 46810
rect 28914 46758 28926 46810
rect 28926 46758 28956 46810
rect 28980 46758 28990 46810
rect 28990 46758 29036 46810
rect 28740 46756 28796 46758
rect 28820 46756 28876 46758
rect 28900 46756 28956 46758
rect 28980 46756 29036 46758
rect 28740 45722 28796 45724
rect 28820 45722 28876 45724
rect 28900 45722 28956 45724
rect 28980 45722 29036 45724
rect 28740 45670 28786 45722
rect 28786 45670 28796 45722
rect 28820 45670 28850 45722
rect 28850 45670 28862 45722
rect 28862 45670 28876 45722
rect 28900 45670 28914 45722
rect 28914 45670 28926 45722
rect 28926 45670 28956 45722
rect 28980 45670 28990 45722
rect 28990 45670 29036 45722
rect 28740 45668 28796 45670
rect 28820 45668 28876 45670
rect 28900 45668 28956 45670
rect 28980 45668 29036 45670
rect 28740 44634 28796 44636
rect 28820 44634 28876 44636
rect 28900 44634 28956 44636
rect 28980 44634 29036 44636
rect 28740 44582 28786 44634
rect 28786 44582 28796 44634
rect 28820 44582 28850 44634
rect 28850 44582 28862 44634
rect 28862 44582 28876 44634
rect 28900 44582 28914 44634
rect 28914 44582 28926 44634
rect 28926 44582 28956 44634
rect 28980 44582 28990 44634
rect 28990 44582 29036 44634
rect 28740 44580 28796 44582
rect 28820 44580 28876 44582
rect 28900 44580 28956 44582
rect 28980 44580 29036 44582
rect 28740 43546 28796 43548
rect 28820 43546 28876 43548
rect 28900 43546 28956 43548
rect 28980 43546 29036 43548
rect 28740 43494 28786 43546
rect 28786 43494 28796 43546
rect 28820 43494 28850 43546
rect 28850 43494 28862 43546
rect 28862 43494 28876 43546
rect 28900 43494 28914 43546
rect 28914 43494 28926 43546
rect 28926 43494 28956 43546
rect 28980 43494 28990 43546
rect 28990 43494 29036 43546
rect 28740 43492 28796 43494
rect 28820 43492 28876 43494
rect 28900 43492 28956 43494
rect 28980 43492 29036 43494
rect 28740 42458 28796 42460
rect 28820 42458 28876 42460
rect 28900 42458 28956 42460
rect 28980 42458 29036 42460
rect 28740 42406 28786 42458
rect 28786 42406 28796 42458
rect 28820 42406 28850 42458
rect 28850 42406 28862 42458
rect 28862 42406 28876 42458
rect 28900 42406 28914 42458
rect 28914 42406 28926 42458
rect 28926 42406 28956 42458
rect 28980 42406 28990 42458
rect 28990 42406 29036 42458
rect 28740 42404 28796 42406
rect 28820 42404 28876 42406
rect 28900 42404 28956 42406
rect 28980 42404 29036 42406
rect 28740 41370 28796 41372
rect 28820 41370 28876 41372
rect 28900 41370 28956 41372
rect 28980 41370 29036 41372
rect 28740 41318 28786 41370
rect 28786 41318 28796 41370
rect 28820 41318 28850 41370
rect 28850 41318 28862 41370
rect 28862 41318 28876 41370
rect 28900 41318 28914 41370
rect 28914 41318 28926 41370
rect 28926 41318 28956 41370
rect 28980 41318 28990 41370
rect 28990 41318 29036 41370
rect 28740 41316 28796 41318
rect 28820 41316 28876 41318
rect 28900 41316 28956 41318
rect 28980 41316 29036 41318
rect 28740 40282 28796 40284
rect 28820 40282 28876 40284
rect 28900 40282 28956 40284
rect 28980 40282 29036 40284
rect 28740 40230 28786 40282
rect 28786 40230 28796 40282
rect 28820 40230 28850 40282
rect 28850 40230 28862 40282
rect 28862 40230 28876 40282
rect 28900 40230 28914 40282
rect 28914 40230 28926 40282
rect 28926 40230 28956 40282
rect 28980 40230 28990 40282
rect 28990 40230 29036 40282
rect 28740 40228 28796 40230
rect 28820 40228 28876 40230
rect 28900 40228 28956 40230
rect 28980 40228 29036 40230
rect 29918 40160 29974 40216
rect 28630 39480 28686 39536
rect 28740 39194 28796 39196
rect 28820 39194 28876 39196
rect 28900 39194 28956 39196
rect 28980 39194 29036 39196
rect 28740 39142 28786 39194
rect 28786 39142 28796 39194
rect 28820 39142 28850 39194
rect 28850 39142 28862 39194
rect 28862 39142 28876 39194
rect 28900 39142 28914 39194
rect 28914 39142 28926 39194
rect 28926 39142 28956 39194
rect 28980 39142 28990 39194
rect 28990 39142 29036 39194
rect 28740 39140 28796 39142
rect 28820 39140 28876 39142
rect 28900 39140 28956 39142
rect 28980 39140 29036 39142
rect 28740 38106 28796 38108
rect 28820 38106 28876 38108
rect 28900 38106 28956 38108
rect 28980 38106 29036 38108
rect 28740 38054 28786 38106
rect 28786 38054 28796 38106
rect 28820 38054 28850 38106
rect 28850 38054 28862 38106
rect 28862 38054 28876 38106
rect 28900 38054 28914 38106
rect 28914 38054 28926 38106
rect 28926 38054 28956 38106
rect 28980 38054 28990 38106
rect 28990 38054 29036 38106
rect 28740 38052 28796 38054
rect 28820 38052 28876 38054
rect 28900 38052 28956 38054
rect 28980 38052 29036 38054
rect 27526 34040 27582 34096
rect 27434 32272 27490 32328
rect 25267 17978 25323 17980
rect 25347 17978 25403 17980
rect 25427 17978 25483 17980
rect 25507 17978 25563 17980
rect 25267 17926 25313 17978
rect 25313 17926 25323 17978
rect 25347 17926 25377 17978
rect 25377 17926 25389 17978
rect 25389 17926 25403 17978
rect 25427 17926 25441 17978
rect 25441 17926 25453 17978
rect 25453 17926 25483 17978
rect 25507 17926 25517 17978
rect 25517 17926 25563 17978
rect 25267 17924 25323 17926
rect 25347 17924 25403 17926
rect 25427 17924 25483 17926
rect 25507 17924 25563 17926
rect 25267 16890 25323 16892
rect 25347 16890 25403 16892
rect 25427 16890 25483 16892
rect 25507 16890 25563 16892
rect 25267 16838 25313 16890
rect 25313 16838 25323 16890
rect 25347 16838 25377 16890
rect 25377 16838 25389 16890
rect 25389 16838 25403 16890
rect 25427 16838 25441 16890
rect 25441 16838 25453 16890
rect 25453 16838 25483 16890
rect 25507 16838 25517 16890
rect 25517 16838 25563 16890
rect 25267 16836 25323 16838
rect 25347 16836 25403 16838
rect 25427 16836 25483 16838
rect 25507 16836 25563 16838
rect 25267 15802 25323 15804
rect 25347 15802 25403 15804
rect 25427 15802 25483 15804
rect 25507 15802 25563 15804
rect 25267 15750 25313 15802
rect 25313 15750 25323 15802
rect 25347 15750 25377 15802
rect 25377 15750 25389 15802
rect 25389 15750 25403 15802
rect 25427 15750 25441 15802
rect 25441 15750 25453 15802
rect 25453 15750 25483 15802
rect 25507 15750 25517 15802
rect 25517 15750 25563 15802
rect 25267 15748 25323 15750
rect 25347 15748 25403 15750
rect 25427 15748 25483 15750
rect 25507 15748 25563 15750
rect 25502 15000 25558 15056
rect 25267 14714 25323 14716
rect 25347 14714 25403 14716
rect 25427 14714 25483 14716
rect 25507 14714 25563 14716
rect 25267 14662 25313 14714
rect 25313 14662 25323 14714
rect 25347 14662 25377 14714
rect 25377 14662 25389 14714
rect 25389 14662 25403 14714
rect 25427 14662 25441 14714
rect 25441 14662 25453 14714
rect 25453 14662 25483 14714
rect 25507 14662 25517 14714
rect 25517 14662 25563 14714
rect 25267 14660 25323 14662
rect 25347 14660 25403 14662
rect 25427 14660 25483 14662
rect 25507 14660 25563 14662
rect 25267 13626 25323 13628
rect 25347 13626 25403 13628
rect 25427 13626 25483 13628
rect 25507 13626 25563 13628
rect 25267 13574 25313 13626
rect 25313 13574 25323 13626
rect 25347 13574 25377 13626
rect 25377 13574 25389 13626
rect 25389 13574 25403 13626
rect 25427 13574 25441 13626
rect 25441 13574 25453 13626
rect 25453 13574 25483 13626
rect 25507 13574 25517 13626
rect 25517 13574 25563 13626
rect 25267 13572 25323 13574
rect 25347 13572 25403 13574
rect 25427 13572 25483 13574
rect 25507 13572 25563 13574
rect 25267 12538 25323 12540
rect 25347 12538 25403 12540
rect 25427 12538 25483 12540
rect 25507 12538 25563 12540
rect 25267 12486 25313 12538
rect 25313 12486 25323 12538
rect 25347 12486 25377 12538
rect 25377 12486 25389 12538
rect 25389 12486 25403 12538
rect 25427 12486 25441 12538
rect 25441 12486 25453 12538
rect 25453 12486 25483 12538
rect 25507 12486 25517 12538
rect 25517 12486 25563 12538
rect 25267 12484 25323 12486
rect 25347 12484 25403 12486
rect 25427 12484 25483 12486
rect 25507 12484 25563 12486
rect 21794 11994 21850 11996
rect 21874 11994 21930 11996
rect 21954 11994 22010 11996
rect 22034 11994 22090 11996
rect 21794 11942 21840 11994
rect 21840 11942 21850 11994
rect 21874 11942 21904 11994
rect 21904 11942 21916 11994
rect 21916 11942 21930 11994
rect 21954 11942 21968 11994
rect 21968 11942 21980 11994
rect 21980 11942 22010 11994
rect 22034 11942 22044 11994
rect 22044 11942 22090 11994
rect 21794 11940 21850 11942
rect 21874 11940 21930 11942
rect 21954 11940 22010 11942
rect 22034 11940 22090 11942
rect 25267 11450 25323 11452
rect 25347 11450 25403 11452
rect 25427 11450 25483 11452
rect 25507 11450 25563 11452
rect 25267 11398 25313 11450
rect 25313 11398 25323 11450
rect 25347 11398 25377 11450
rect 25377 11398 25389 11450
rect 25389 11398 25403 11450
rect 25427 11398 25441 11450
rect 25441 11398 25453 11450
rect 25453 11398 25483 11450
rect 25507 11398 25517 11450
rect 25517 11398 25563 11450
rect 25267 11396 25323 11398
rect 25347 11396 25403 11398
rect 25427 11396 25483 11398
rect 25507 11396 25563 11398
rect 21794 10906 21850 10908
rect 21874 10906 21930 10908
rect 21954 10906 22010 10908
rect 22034 10906 22090 10908
rect 21794 10854 21840 10906
rect 21840 10854 21850 10906
rect 21874 10854 21904 10906
rect 21904 10854 21916 10906
rect 21916 10854 21930 10906
rect 21954 10854 21968 10906
rect 21968 10854 21980 10906
rect 21980 10854 22010 10906
rect 22034 10854 22044 10906
rect 22044 10854 22090 10906
rect 21794 10852 21850 10854
rect 21874 10852 21930 10854
rect 21954 10852 22010 10854
rect 22034 10852 22090 10854
rect 25267 10362 25323 10364
rect 25347 10362 25403 10364
rect 25427 10362 25483 10364
rect 25507 10362 25563 10364
rect 25267 10310 25313 10362
rect 25313 10310 25323 10362
rect 25347 10310 25377 10362
rect 25377 10310 25389 10362
rect 25389 10310 25403 10362
rect 25427 10310 25441 10362
rect 25441 10310 25453 10362
rect 25453 10310 25483 10362
rect 25507 10310 25517 10362
rect 25517 10310 25563 10362
rect 25267 10308 25323 10310
rect 25347 10308 25403 10310
rect 25427 10308 25483 10310
rect 25507 10308 25563 10310
rect 21794 9818 21850 9820
rect 21874 9818 21930 9820
rect 21954 9818 22010 9820
rect 22034 9818 22090 9820
rect 21794 9766 21840 9818
rect 21840 9766 21850 9818
rect 21874 9766 21904 9818
rect 21904 9766 21916 9818
rect 21916 9766 21930 9818
rect 21954 9766 21968 9818
rect 21968 9766 21980 9818
rect 21980 9766 22010 9818
rect 22034 9766 22044 9818
rect 22044 9766 22090 9818
rect 21794 9764 21850 9766
rect 21874 9764 21930 9766
rect 21954 9764 22010 9766
rect 22034 9764 22090 9766
rect 18321 9274 18377 9276
rect 18401 9274 18457 9276
rect 18481 9274 18537 9276
rect 18561 9274 18617 9276
rect 18321 9222 18367 9274
rect 18367 9222 18377 9274
rect 18401 9222 18431 9274
rect 18431 9222 18443 9274
rect 18443 9222 18457 9274
rect 18481 9222 18495 9274
rect 18495 9222 18507 9274
rect 18507 9222 18537 9274
rect 18561 9222 18571 9274
rect 18571 9222 18617 9274
rect 18321 9220 18377 9222
rect 18401 9220 18457 9222
rect 18481 9220 18537 9222
rect 18561 9220 18617 9222
rect 18321 8186 18377 8188
rect 18401 8186 18457 8188
rect 18481 8186 18537 8188
rect 18561 8186 18617 8188
rect 18321 8134 18367 8186
rect 18367 8134 18377 8186
rect 18401 8134 18431 8186
rect 18431 8134 18443 8186
rect 18443 8134 18457 8186
rect 18481 8134 18495 8186
rect 18495 8134 18507 8186
rect 18507 8134 18537 8186
rect 18561 8134 18571 8186
rect 18571 8134 18617 8186
rect 18321 8132 18377 8134
rect 18401 8132 18457 8134
rect 18481 8132 18537 8134
rect 18561 8132 18617 8134
rect 18321 7098 18377 7100
rect 18401 7098 18457 7100
rect 18481 7098 18537 7100
rect 18561 7098 18617 7100
rect 18321 7046 18367 7098
rect 18367 7046 18377 7098
rect 18401 7046 18431 7098
rect 18431 7046 18443 7098
rect 18443 7046 18457 7098
rect 18481 7046 18495 7098
rect 18495 7046 18507 7098
rect 18507 7046 18537 7098
rect 18561 7046 18571 7098
rect 18571 7046 18617 7098
rect 18321 7044 18377 7046
rect 18401 7044 18457 7046
rect 18481 7044 18537 7046
rect 18561 7044 18617 7046
rect 18321 6010 18377 6012
rect 18401 6010 18457 6012
rect 18481 6010 18537 6012
rect 18561 6010 18617 6012
rect 18321 5958 18367 6010
rect 18367 5958 18377 6010
rect 18401 5958 18431 6010
rect 18431 5958 18443 6010
rect 18443 5958 18457 6010
rect 18481 5958 18495 6010
rect 18495 5958 18507 6010
rect 18507 5958 18537 6010
rect 18561 5958 18571 6010
rect 18571 5958 18617 6010
rect 18321 5956 18377 5958
rect 18401 5956 18457 5958
rect 18481 5956 18537 5958
rect 18561 5956 18617 5958
rect 18321 4922 18377 4924
rect 18401 4922 18457 4924
rect 18481 4922 18537 4924
rect 18561 4922 18617 4924
rect 18321 4870 18367 4922
rect 18367 4870 18377 4922
rect 18401 4870 18431 4922
rect 18431 4870 18443 4922
rect 18443 4870 18457 4922
rect 18481 4870 18495 4922
rect 18495 4870 18507 4922
rect 18507 4870 18537 4922
rect 18561 4870 18571 4922
rect 18571 4870 18617 4922
rect 18321 4868 18377 4870
rect 18401 4868 18457 4870
rect 18481 4868 18537 4870
rect 18561 4868 18617 4870
rect 25267 9274 25323 9276
rect 25347 9274 25403 9276
rect 25427 9274 25483 9276
rect 25507 9274 25563 9276
rect 25267 9222 25313 9274
rect 25313 9222 25323 9274
rect 25347 9222 25377 9274
rect 25377 9222 25389 9274
rect 25389 9222 25403 9274
rect 25427 9222 25441 9274
rect 25441 9222 25453 9274
rect 25453 9222 25483 9274
rect 25507 9222 25517 9274
rect 25517 9222 25563 9274
rect 25267 9220 25323 9222
rect 25347 9220 25403 9222
rect 25427 9220 25483 9222
rect 25507 9220 25563 9222
rect 21794 8730 21850 8732
rect 21874 8730 21930 8732
rect 21954 8730 22010 8732
rect 22034 8730 22090 8732
rect 21794 8678 21840 8730
rect 21840 8678 21850 8730
rect 21874 8678 21904 8730
rect 21904 8678 21916 8730
rect 21916 8678 21930 8730
rect 21954 8678 21968 8730
rect 21968 8678 21980 8730
rect 21980 8678 22010 8730
rect 22034 8678 22044 8730
rect 22044 8678 22090 8730
rect 21794 8676 21850 8678
rect 21874 8676 21930 8678
rect 21954 8676 22010 8678
rect 22034 8676 22090 8678
rect 26146 8200 26202 8256
rect 25267 8186 25323 8188
rect 25347 8186 25403 8188
rect 25427 8186 25483 8188
rect 25507 8186 25563 8188
rect 25267 8134 25313 8186
rect 25313 8134 25323 8186
rect 25347 8134 25377 8186
rect 25377 8134 25389 8186
rect 25389 8134 25403 8186
rect 25427 8134 25441 8186
rect 25441 8134 25453 8186
rect 25453 8134 25483 8186
rect 25507 8134 25517 8186
rect 25517 8134 25563 8186
rect 25267 8132 25323 8134
rect 25347 8132 25403 8134
rect 25427 8132 25483 8134
rect 25507 8132 25563 8134
rect 21794 7642 21850 7644
rect 21874 7642 21930 7644
rect 21954 7642 22010 7644
rect 22034 7642 22090 7644
rect 21794 7590 21840 7642
rect 21840 7590 21850 7642
rect 21874 7590 21904 7642
rect 21904 7590 21916 7642
rect 21916 7590 21930 7642
rect 21954 7590 21968 7642
rect 21968 7590 21980 7642
rect 21980 7590 22010 7642
rect 22034 7590 22044 7642
rect 22044 7590 22090 7642
rect 21794 7588 21850 7590
rect 21874 7588 21930 7590
rect 21954 7588 22010 7590
rect 22034 7588 22090 7590
rect 25267 7098 25323 7100
rect 25347 7098 25403 7100
rect 25427 7098 25483 7100
rect 25507 7098 25563 7100
rect 25267 7046 25313 7098
rect 25313 7046 25323 7098
rect 25347 7046 25377 7098
rect 25377 7046 25389 7098
rect 25389 7046 25403 7098
rect 25427 7046 25441 7098
rect 25441 7046 25453 7098
rect 25453 7046 25483 7098
rect 25507 7046 25517 7098
rect 25517 7046 25563 7098
rect 25267 7044 25323 7046
rect 25347 7044 25403 7046
rect 25427 7044 25483 7046
rect 25507 7044 25563 7046
rect 21794 6554 21850 6556
rect 21874 6554 21930 6556
rect 21954 6554 22010 6556
rect 22034 6554 22090 6556
rect 21794 6502 21840 6554
rect 21840 6502 21850 6554
rect 21874 6502 21904 6554
rect 21904 6502 21916 6554
rect 21916 6502 21930 6554
rect 21954 6502 21968 6554
rect 21968 6502 21980 6554
rect 21980 6502 22010 6554
rect 22034 6502 22044 6554
rect 22044 6502 22090 6554
rect 21794 6500 21850 6502
rect 21874 6500 21930 6502
rect 21954 6500 22010 6502
rect 22034 6500 22090 6502
rect 25267 6010 25323 6012
rect 25347 6010 25403 6012
rect 25427 6010 25483 6012
rect 25507 6010 25563 6012
rect 25267 5958 25313 6010
rect 25313 5958 25323 6010
rect 25347 5958 25377 6010
rect 25377 5958 25389 6010
rect 25389 5958 25403 6010
rect 25427 5958 25441 6010
rect 25441 5958 25453 6010
rect 25453 5958 25483 6010
rect 25507 5958 25517 6010
rect 25517 5958 25563 6010
rect 25267 5956 25323 5958
rect 25347 5956 25403 5958
rect 25427 5956 25483 5958
rect 25507 5956 25563 5958
rect 21794 5466 21850 5468
rect 21874 5466 21930 5468
rect 21954 5466 22010 5468
rect 22034 5466 22090 5468
rect 21794 5414 21840 5466
rect 21840 5414 21850 5466
rect 21874 5414 21904 5466
rect 21904 5414 21916 5466
rect 21916 5414 21930 5466
rect 21954 5414 21968 5466
rect 21968 5414 21980 5466
rect 21980 5414 22010 5466
rect 22034 5414 22044 5466
rect 22044 5414 22090 5466
rect 21794 5412 21850 5414
rect 21874 5412 21930 5414
rect 21954 5412 22010 5414
rect 22034 5412 22090 5414
rect 25267 4922 25323 4924
rect 25347 4922 25403 4924
rect 25427 4922 25483 4924
rect 25507 4922 25563 4924
rect 25267 4870 25313 4922
rect 25313 4870 25323 4922
rect 25347 4870 25377 4922
rect 25377 4870 25389 4922
rect 25389 4870 25403 4922
rect 25427 4870 25441 4922
rect 25441 4870 25453 4922
rect 25453 4870 25483 4922
rect 25507 4870 25517 4922
rect 25517 4870 25563 4922
rect 25267 4868 25323 4870
rect 25347 4868 25403 4870
rect 25427 4868 25483 4870
rect 25507 4868 25563 4870
rect 18321 3834 18377 3836
rect 18401 3834 18457 3836
rect 18481 3834 18537 3836
rect 18561 3834 18617 3836
rect 18321 3782 18367 3834
rect 18367 3782 18377 3834
rect 18401 3782 18431 3834
rect 18431 3782 18443 3834
rect 18443 3782 18457 3834
rect 18481 3782 18495 3834
rect 18495 3782 18507 3834
rect 18507 3782 18537 3834
rect 18561 3782 18571 3834
rect 18571 3782 18617 3834
rect 18321 3780 18377 3782
rect 18401 3780 18457 3782
rect 18481 3780 18537 3782
rect 18561 3780 18617 3782
rect 18321 2746 18377 2748
rect 18401 2746 18457 2748
rect 18481 2746 18537 2748
rect 18561 2746 18617 2748
rect 18321 2694 18367 2746
rect 18367 2694 18377 2746
rect 18401 2694 18431 2746
rect 18431 2694 18443 2746
rect 18443 2694 18457 2746
rect 18481 2694 18495 2746
rect 18495 2694 18507 2746
rect 18507 2694 18537 2746
rect 18561 2694 18571 2746
rect 18571 2694 18617 2746
rect 18321 2692 18377 2694
rect 18401 2692 18457 2694
rect 18481 2692 18537 2694
rect 18561 2692 18617 2694
rect 21794 4378 21850 4380
rect 21874 4378 21930 4380
rect 21954 4378 22010 4380
rect 22034 4378 22090 4380
rect 21794 4326 21840 4378
rect 21840 4326 21850 4378
rect 21874 4326 21904 4378
rect 21904 4326 21916 4378
rect 21916 4326 21930 4378
rect 21954 4326 21968 4378
rect 21968 4326 21980 4378
rect 21980 4326 22010 4378
rect 22034 4326 22044 4378
rect 22044 4326 22090 4378
rect 21794 4324 21850 4326
rect 21874 4324 21930 4326
rect 21954 4324 22010 4326
rect 22034 4324 22090 4326
rect 25267 3834 25323 3836
rect 25347 3834 25403 3836
rect 25427 3834 25483 3836
rect 25507 3834 25563 3836
rect 25267 3782 25313 3834
rect 25313 3782 25323 3834
rect 25347 3782 25377 3834
rect 25377 3782 25389 3834
rect 25389 3782 25403 3834
rect 25427 3782 25441 3834
rect 25441 3782 25453 3834
rect 25453 3782 25483 3834
rect 25507 3782 25517 3834
rect 25517 3782 25563 3834
rect 25267 3780 25323 3782
rect 25347 3780 25403 3782
rect 25427 3780 25483 3782
rect 25507 3780 25563 3782
rect 27526 30640 27582 30696
rect 27526 28600 27582 28656
rect 27526 27532 27582 27568
rect 27526 27512 27528 27532
rect 27528 27512 27580 27532
rect 27580 27512 27582 27532
rect 27526 25200 27582 25256
rect 27526 21120 27582 21176
rect 27526 20440 27582 20496
rect 27526 14320 27582 14376
rect 27526 10240 27582 10296
rect 21794 3290 21850 3292
rect 21874 3290 21930 3292
rect 21954 3290 22010 3292
rect 22034 3290 22090 3292
rect 21794 3238 21840 3290
rect 21840 3238 21850 3290
rect 21874 3238 21904 3290
rect 21904 3238 21916 3290
rect 21916 3238 21930 3290
rect 21954 3238 21968 3290
rect 21968 3238 21980 3290
rect 21980 3238 22010 3290
rect 22034 3238 22044 3290
rect 22044 3238 22090 3290
rect 21794 3236 21850 3238
rect 21874 3236 21930 3238
rect 21954 3236 22010 3238
rect 22034 3236 22090 3238
rect 26146 3440 26202 3496
rect 21794 2202 21850 2204
rect 21874 2202 21930 2204
rect 21954 2202 22010 2204
rect 22034 2202 22090 2204
rect 21794 2150 21840 2202
rect 21840 2150 21850 2202
rect 21874 2150 21904 2202
rect 21904 2150 21916 2202
rect 21916 2150 21930 2202
rect 21954 2150 21968 2202
rect 21968 2150 21980 2202
rect 21980 2150 22010 2202
rect 22034 2150 22044 2202
rect 22044 2150 22090 2202
rect 21794 2148 21850 2150
rect 21874 2148 21930 2150
rect 21954 2148 22010 2150
rect 22034 2148 22090 2150
rect 26146 2760 26202 2816
rect 25267 2746 25323 2748
rect 25347 2746 25403 2748
rect 25427 2746 25483 2748
rect 25507 2746 25563 2748
rect 25267 2694 25313 2746
rect 25313 2694 25323 2746
rect 25347 2694 25377 2746
rect 25377 2694 25389 2746
rect 25389 2694 25403 2746
rect 25427 2694 25441 2746
rect 25441 2694 25453 2746
rect 25453 2694 25483 2746
rect 25507 2694 25517 2746
rect 25517 2694 25563 2746
rect 25267 2692 25323 2694
rect 25347 2692 25403 2694
rect 25427 2692 25483 2694
rect 25507 2692 25563 2694
rect 27526 5208 27582 5264
rect 27434 2488 27490 2544
rect 28740 37018 28796 37020
rect 28820 37018 28876 37020
rect 28900 37018 28956 37020
rect 28980 37018 29036 37020
rect 28740 36966 28786 37018
rect 28786 36966 28796 37018
rect 28820 36966 28850 37018
rect 28850 36966 28862 37018
rect 28862 36966 28876 37018
rect 28900 36966 28914 37018
rect 28914 36966 28926 37018
rect 28926 36966 28956 37018
rect 28980 36966 28990 37018
rect 28990 36966 29036 37018
rect 28740 36964 28796 36966
rect 28820 36964 28876 36966
rect 28900 36964 28956 36966
rect 28980 36964 29036 36966
rect 28740 35930 28796 35932
rect 28820 35930 28876 35932
rect 28900 35930 28956 35932
rect 28980 35930 29036 35932
rect 28740 35878 28786 35930
rect 28786 35878 28796 35930
rect 28820 35878 28850 35930
rect 28850 35878 28862 35930
rect 28862 35878 28876 35930
rect 28900 35878 28914 35930
rect 28914 35878 28926 35930
rect 28926 35878 28956 35930
rect 28980 35878 28990 35930
rect 28990 35878 29036 35930
rect 28740 35876 28796 35878
rect 28820 35876 28876 35878
rect 28900 35876 28956 35878
rect 28980 35876 29036 35878
rect 28740 34842 28796 34844
rect 28820 34842 28876 34844
rect 28900 34842 28956 34844
rect 28980 34842 29036 34844
rect 28740 34790 28786 34842
rect 28786 34790 28796 34842
rect 28820 34790 28850 34842
rect 28850 34790 28862 34842
rect 28862 34790 28876 34842
rect 28900 34790 28914 34842
rect 28914 34790 28926 34842
rect 28926 34790 28956 34842
rect 28980 34790 28990 34842
rect 28990 34790 29036 34842
rect 28740 34788 28796 34790
rect 28820 34788 28876 34790
rect 28900 34788 28956 34790
rect 28980 34788 29036 34790
rect 28740 33754 28796 33756
rect 28820 33754 28876 33756
rect 28900 33754 28956 33756
rect 28980 33754 29036 33756
rect 28740 33702 28786 33754
rect 28786 33702 28796 33754
rect 28820 33702 28850 33754
rect 28850 33702 28862 33754
rect 28862 33702 28876 33754
rect 28900 33702 28914 33754
rect 28914 33702 28926 33754
rect 28926 33702 28956 33754
rect 28980 33702 28990 33754
rect 28990 33702 29036 33754
rect 28740 33700 28796 33702
rect 28820 33700 28876 33702
rect 28900 33700 28956 33702
rect 28980 33700 29036 33702
rect 28740 32666 28796 32668
rect 28820 32666 28876 32668
rect 28900 32666 28956 32668
rect 28980 32666 29036 32668
rect 28740 32614 28786 32666
rect 28786 32614 28796 32666
rect 28820 32614 28850 32666
rect 28850 32614 28862 32666
rect 28862 32614 28876 32666
rect 28900 32614 28914 32666
rect 28914 32614 28926 32666
rect 28926 32614 28956 32666
rect 28980 32614 28990 32666
rect 28990 32614 29036 32666
rect 28740 32612 28796 32614
rect 28820 32612 28876 32614
rect 28900 32612 28956 32614
rect 28980 32612 29036 32614
rect 28354 32000 28410 32056
rect 28740 31578 28796 31580
rect 28820 31578 28876 31580
rect 28900 31578 28956 31580
rect 28980 31578 29036 31580
rect 28740 31526 28786 31578
rect 28786 31526 28796 31578
rect 28820 31526 28850 31578
rect 28850 31526 28862 31578
rect 28862 31526 28876 31578
rect 28900 31526 28914 31578
rect 28914 31526 28926 31578
rect 28926 31526 28956 31578
rect 28980 31526 28990 31578
rect 28990 31526 29036 31578
rect 28740 31524 28796 31526
rect 28820 31524 28876 31526
rect 28900 31524 28956 31526
rect 28980 31524 29036 31526
rect 28740 30490 28796 30492
rect 28820 30490 28876 30492
rect 28900 30490 28956 30492
rect 28980 30490 29036 30492
rect 28740 30438 28786 30490
rect 28786 30438 28796 30490
rect 28820 30438 28850 30490
rect 28850 30438 28862 30490
rect 28862 30438 28876 30490
rect 28900 30438 28914 30490
rect 28914 30438 28926 30490
rect 28926 30438 28956 30490
rect 28980 30438 28990 30490
rect 28990 30438 29036 30490
rect 28740 30436 28796 30438
rect 28820 30436 28876 30438
rect 28900 30436 28956 30438
rect 28980 30436 29036 30438
rect 28740 29402 28796 29404
rect 28820 29402 28876 29404
rect 28900 29402 28956 29404
rect 28980 29402 29036 29404
rect 28740 29350 28786 29402
rect 28786 29350 28796 29402
rect 28820 29350 28850 29402
rect 28850 29350 28862 29402
rect 28862 29350 28876 29402
rect 28900 29350 28914 29402
rect 28914 29350 28926 29402
rect 28926 29350 28956 29402
rect 28980 29350 28990 29402
rect 28990 29350 29036 29402
rect 28740 29348 28796 29350
rect 28820 29348 28876 29350
rect 28900 29348 28956 29350
rect 28980 29348 29036 29350
rect 28740 28314 28796 28316
rect 28820 28314 28876 28316
rect 28900 28314 28956 28316
rect 28980 28314 29036 28316
rect 28740 28262 28786 28314
rect 28786 28262 28796 28314
rect 28820 28262 28850 28314
rect 28850 28262 28862 28314
rect 28862 28262 28876 28314
rect 28900 28262 28914 28314
rect 28914 28262 28926 28314
rect 28926 28262 28956 28314
rect 28980 28262 28990 28314
rect 28990 28262 29036 28314
rect 28740 28260 28796 28262
rect 28820 28260 28876 28262
rect 28900 28260 28956 28262
rect 28980 28260 29036 28262
rect 28740 27226 28796 27228
rect 28820 27226 28876 27228
rect 28900 27226 28956 27228
rect 28980 27226 29036 27228
rect 28740 27174 28786 27226
rect 28786 27174 28796 27226
rect 28820 27174 28850 27226
rect 28850 27174 28862 27226
rect 28862 27174 28876 27226
rect 28900 27174 28914 27226
rect 28914 27174 28926 27226
rect 28926 27174 28956 27226
rect 28980 27174 28990 27226
rect 28990 27174 29036 27226
rect 28740 27172 28796 27174
rect 28820 27172 28876 27174
rect 28900 27172 28956 27174
rect 28980 27172 29036 27174
rect 28354 26560 28410 26616
rect 28740 26138 28796 26140
rect 28820 26138 28876 26140
rect 28900 26138 28956 26140
rect 28980 26138 29036 26140
rect 28740 26086 28786 26138
rect 28786 26086 28796 26138
rect 28820 26086 28850 26138
rect 28850 26086 28862 26138
rect 28862 26086 28876 26138
rect 28900 26086 28914 26138
rect 28914 26086 28926 26138
rect 28926 26086 28956 26138
rect 28980 26086 28990 26138
rect 28990 26086 29036 26138
rect 28740 26084 28796 26086
rect 28820 26084 28876 26086
rect 28900 26084 28956 26086
rect 28980 26084 29036 26086
rect 28740 25050 28796 25052
rect 28820 25050 28876 25052
rect 28900 25050 28956 25052
rect 28980 25050 29036 25052
rect 28740 24998 28786 25050
rect 28786 24998 28796 25050
rect 28820 24998 28850 25050
rect 28850 24998 28862 25050
rect 28862 24998 28876 25050
rect 28900 24998 28914 25050
rect 28914 24998 28926 25050
rect 28926 24998 28956 25050
rect 28980 24998 28990 25050
rect 28990 24998 29036 25050
rect 28740 24996 28796 24998
rect 28820 24996 28876 24998
rect 28900 24996 28956 24998
rect 28980 24996 29036 24998
rect 28354 24520 28410 24576
rect 28740 23962 28796 23964
rect 28820 23962 28876 23964
rect 28900 23962 28956 23964
rect 28980 23962 29036 23964
rect 28740 23910 28786 23962
rect 28786 23910 28796 23962
rect 28820 23910 28850 23962
rect 28850 23910 28862 23962
rect 28862 23910 28876 23962
rect 28900 23910 28914 23962
rect 28914 23910 28926 23962
rect 28926 23910 28956 23962
rect 28980 23910 28990 23962
rect 28990 23910 29036 23962
rect 28740 23908 28796 23910
rect 28820 23908 28876 23910
rect 28900 23908 28956 23910
rect 28980 23908 29036 23910
rect 29918 23840 29974 23896
rect 28740 22874 28796 22876
rect 28820 22874 28876 22876
rect 28900 22874 28956 22876
rect 28980 22874 29036 22876
rect 28740 22822 28786 22874
rect 28786 22822 28796 22874
rect 28820 22822 28850 22874
rect 28850 22822 28862 22874
rect 28862 22822 28876 22874
rect 28900 22822 28914 22874
rect 28914 22822 28926 22874
rect 28926 22822 28956 22874
rect 28980 22822 28990 22874
rect 28990 22822 29036 22874
rect 28740 22820 28796 22822
rect 28820 22820 28876 22822
rect 28900 22820 28956 22822
rect 28980 22820 29036 22822
rect 28740 21786 28796 21788
rect 28820 21786 28876 21788
rect 28900 21786 28956 21788
rect 28980 21786 29036 21788
rect 28740 21734 28786 21786
rect 28786 21734 28796 21786
rect 28820 21734 28850 21786
rect 28850 21734 28862 21786
rect 28862 21734 28876 21786
rect 28900 21734 28914 21786
rect 28914 21734 28926 21786
rect 28926 21734 28956 21786
rect 28980 21734 28990 21786
rect 28990 21734 29036 21786
rect 28740 21732 28796 21734
rect 28820 21732 28876 21734
rect 28900 21732 28956 21734
rect 28980 21732 29036 21734
rect 28740 20698 28796 20700
rect 28820 20698 28876 20700
rect 28900 20698 28956 20700
rect 28980 20698 29036 20700
rect 28740 20646 28786 20698
rect 28786 20646 28796 20698
rect 28820 20646 28850 20698
rect 28850 20646 28862 20698
rect 28862 20646 28876 20698
rect 28900 20646 28914 20698
rect 28914 20646 28926 20698
rect 28926 20646 28956 20698
rect 28980 20646 28990 20698
rect 28990 20646 29036 20698
rect 28740 20644 28796 20646
rect 28820 20644 28876 20646
rect 28900 20644 28956 20646
rect 28980 20644 29036 20646
rect 28630 19760 28686 19816
rect 28740 19610 28796 19612
rect 28820 19610 28876 19612
rect 28900 19610 28956 19612
rect 28980 19610 29036 19612
rect 28740 19558 28786 19610
rect 28786 19558 28796 19610
rect 28820 19558 28850 19610
rect 28850 19558 28862 19610
rect 28862 19558 28876 19610
rect 28900 19558 28914 19610
rect 28914 19558 28926 19610
rect 28926 19558 28956 19610
rect 28980 19558 28990 19610
rect 28990 19558 29036 19610
rect 28740 19556 28796 19558
rect 28820 19556 28876 19558
rect 28900 19556 28956 19558
rect 28980 19556 29036 19558
rect 28740 18522 28796 18524
rect 28820 18522 28876 18524
rect 28900 18522 28956 18524
rect 28980 18522 29036 18524
rect 28740 18470 28786 18522
rect 28786 18470 28796 18522
rect 28820 18470 28850 18522
rect 28850 18470 28862 18522
rect 28862 18470 28876 18522
rect 28900 18470 28914 18522
rect 28914 18470 28926 18522
rect 28926 18470 28956 18522
rect 28980 18470 28990 18522
rect 28990 18470 29036 18522
rect 28740 18468 28796 18470
rect 28820 18468 28876 18470
rect 28900 18468 28956 18470
rect 28980 18468 29036 18470
rect 28740 17434 28796 17436
rect 28820 17434 28876 17436
rect 28900 17434 28956 17436
rect 28980 17434 29036 17436
rect 28740 17382 28786 17434
rect 28786 17382 28796 17434
rect 28820 17382 28850 17434
rect 28850 17382 28862 17434
rect 28862 17382 28876 17434
rect 28900 17382 28914 17434
rect 28914 17382 28926 17434
rect 28926 17382 28956 17434
rect 28980 17382 28990 17434
rect 28990 17382 29036 17434
rect 28740 17380 28796 17382
rect 28820 17380 28876 17382
rect 28900 17380 28956 17382
rect 28980 17380 29036 17382
rect 29918 16360 29974 16416
rect 28740 16346 28796 16348
rect 28820 16346 28876 16348
rect 28900 16346 28956 16348
rect 28980 16346 29036 16348
rect 28740 16294 28786 16346
rect 28786 16294 28796 16346
rect 28820 16294 28850 16346
rect 28850 16294 28862 16346
rect 28862 16294 28876 16346
rect 28900 16294 28914 16346
rect 28914 16294 28926 16346
rect 28926 16294 28956 16346
rect 28980 16294 28990 16346
rect 28990 16294 29036 16346
rect 28740 16292 28796 16294
rect 28820 16292 28876 16294
rect 28900 16292 28956 16294
rect 28980 16292 29036 16294
rect 28630 15680 28686 15736
rect 28740 15258 28796 15260
rect 28820 15258 28876 15260
rect 28900 15258 28956 15260
rect 28980 15258 29036 15260
rect 28740 15206 28786 15258
rect 28786 15206 28796 15258
rect 28820 15206 28850 15258
rect 28850 15206 28862 15258
rect 28862 15206 28876 15258
rect 28900 15206 28914 15258
rect 28914 15206 28926 15258
rect 28926 15206 28956 15258
rect 28980 15206 28990 15258
rect 28990 15206 29036 15258
rect 28740 15204 28796 15206
rect 28820 15204 28876 15206
rect 28900 15204 28956 15206
rect 28980 15204 29036 15206
rect 28740 14170 28796 14172
rect 28820 14170 28876 14172
rect 28900 14170 28956 14172
rect 28980 14170 29036 14172
rect 28740 14118 28786 14170
rect 28786 14118 28796 14170
rect 28820 14118 28850 14170
rect 28850 14118 28862 14170
rect 28862 14118 28876 14170
rect 28900 14118 28914 14170
rect 28914 14118 28926 14170
rect 28926 14118 28956 14170
rect 28980 14118 28990 14170
rect 28990 14118 29036 14170
rect 28740 14116 28796 14118
rect 28820 14116 28876 14118
rect 28900 14116 28956 14118
rect 28980 14116 29036 14118
rect 28740 13082 28796 13084
rect 28820 13082 28876 13084
rect 28900 13082 28956 13084
rect 28980 13082 29036 13084
rect 28740 13030 28786 13082
rect 28786 13030 28796 13082
rect 28820 13030 28850 13082
rect 28850 13030 28862 13082
rect 28862 13030 28876 13082
rect 28900 13030 28914 13082
rect 28914 13030 28926 13082
rect 28926 13030 28956 13082
rect 28980 13030 28990 13082
rect 28990 13030 29036 13082
rect 28740 13028 28796 13030
rect 28820 13028 28876 13030
rect 28900 13028 28956 13030
rect 28980 13028 29036 13030
rect 28354 12300 28410 12336
rect 28354 12280 28356 12300
rect 28356 12280 28408 12300
rect 28408 12280 28410 12300
rect 28740 11994 28796 11996
rect 28820 11994 28876 11996
rect 28900 11994 28956 11996
rect 28980 11994 29036 11996
rect 28740 11942 28786 11994
rect 28786 11942 28796 11994
rect 28820 11942 28850 11994
rect 28850 11942 28862 11994
rect 28862 11942 28876 11994
rect 28900 11942 28914 11994
rect 28914 11942 28926 11994
rect 28926 11942 28956 11994
rect 28980 11942 28990 11994
rect 28990 11942 29036 11994
rect 28740 11940 28796 11942
rect 28820 11940 28876 11942
rect 28900 11940 28956 11942
rect 28980 11940 29036 11942
rect 29918 10920 29974 10976
rect 28740 10906 28796 10908
rect 28820 10906 28876 10908
rect 28900 10906 28956 10908
rect 28980 10906 29036 10908
rect 28740 10854 28786 10906
rect 28786 10854 28796 10906
rect 28820 10854 28850 10906
rect 28850 10854 28862 10906
rect 28862 10854 28876 10906
rect 28900 10854 28914 10906
rect 28914 10854 28926 10906
rect 28926 10854 28956 10906
rect 28980 10854 28990 10906
rect 28990 10854 29036 10906
rect 28740 10852 28796 10854
rect 28820 10852 28876 10854
rect 28900 10852 28956 10854
rect 28980 10852 29036 10854
rect 28740 9818 28796 9820
rect 28820 9818 28876 9820
rect 28900 9818 28956 9820
rect 28980 9818 29036 9820
rect 28740 9766 28786 9818
rect 28786 9766 28796 9818
rect 28820 9766 28850 9818
rect 28850 9766 28862 9818
rect 28862 9766 28876 9818
rect 28900 9766 28914 9818
rect 28914 9766 28926 9818
rect 28926 9766 28956 9818
rect 28980 9766 28990 9818
rect 28990 9766 29036 9818
rect 28740 9764 28796 9766
rect 28820 9764 28876 9766
rect 28900 9764 28956 9766
rect 28980 9764 29036 9766
rect 28354 8916 28356 8936
rect 28356 8916 28408 8936
rect 28408 8916 28410 8936
rect 28354 8880 28410 8916
rect 28740 8730 28796 8732
rect 28820 8730 28876 8732
rect 28900 8730 28956 8732
rect 28980 8730 29036 8732
rect 28740 8678 28786 8730
rect 28786 8678 28796 8730
rect 28820 8678 28850 8730
rect 28850 8678 28862 8730
rect 28862 8678 28876 8730
rect 28900 8678 28914 8730
rect 28914 8678 28926 8730
rect 28926 8678 28956 8730
rect 28980 8678 28990 8730
rect 28990 8678 29036 8730
rect 28740 8676 28796 8678
rect 28820 8676 28876 8678
rect 28900 8676 28956 8678
rect 28980 8676 29036 8678
rect 28740 7642 28796 7644
rect 28820 7642 28876 7644
rect 28900 7642 28956 7644
rect 28980 7642 29036 7644
rect 28740 7590 28786 7642
rect 28786 7590 28796 7642
rect 28820 7590 28850 7642
rect 28850 7590 28862 7642
rect 28862 7590 28876 7642
rect 28900 7590 28914 7642
rect 28914 7590 28926 7642
rect 28926 7590 28956 7642
rect 28980 7590 28990 7642
rect 28990 7590 29036 7642
rect 28740 7588 28796 7590
rect 28820 7588 28876 7590
rect 28900 7588 28956 7590
rect 28980 7588 29036 7590
rect 29918 7520 29974 7576
rect 28354 6860 28410 6896
rect 28354 6840 28356 6860
rect 28356 6840 28408 6860
rect 28408 6840 28410 6860
rect 28740 6554 28796 6556
rect 28820 6554 28876 6556
rect 28900 6554 28956 6556
rect 28980 6554 29036 6556
rect 28740 6502 28786 6554
rect 28786 6502 28796 6554
rect 28820 6502 28850 6554
rect 28850 6502 28862 6554
rect 28862 6502 28876 6554
rect 28900 6502 28914 6554
rect 28914 6502 28926 6554
rect 28926 6502 28956 6554
rect 28980 6502 28990 6554
rect 28990 6502 29036 6554
rect 28740 6500 28796 6502
rect 28820 6500 28876 6502
rect 28900 6500 28956 6502
rect 28980 6500 29036 6502
rect 28740 5466 28796 5468
rect 28820 5466 28876 5468
rect 28900 5466 28956 5468
rect 28980 5466 29036 5468
rect 28740 5414 28786 5466
rect 28786 5414 28796 5466
rect 28820 5414 28850 5466
rect 28850 5414 28862 5466
rect 28862 5414 28876 5466
rect 28900 5414 28914 5466
rect 28914 5414 28926 5466
rect 28926 5414 28956 5466
rect 28980 5414 28990 5466
rect 28990 5414 29036 5466
rect 28740 5412 28796 5414
rect 28820 5412 28876 5414
rect 28900 5412 28956 5414
rect 28980 5412 29036 5414
rect 28740 4378 28796 4380
rect 28820 4378 28876 4380
rect 28900 4378 28956 4380
rect 28980 4378 29036 4380
rect 28740 4326 28786 4378
rect 28786 4326 28796 4378
rect 28820 4326 28850 4378
rect 28850 4326 28862 4378
rect 28862 4326 28876 4378
rect 28900 4326 28914 4378
rect 28914 4326 28926 4378
rect 28926 4326 28956 4378
rect 28980 4326 28990 4378
rect 28990 4326 29036 4378
rect 28740 4324 28796 4326
rect 28820 4324 28876 4326
rect 28900 4324 28956 4326
rect 28980 4324 29036 4326
rect 28740 3290 28796 3292
rect 28820 3290 28876 3292
rect 28900 3290 28956 3292
rect 28980 3290 29036 3292
rect 28740 3238 28786 3290
rect 28786 3238 28796 3290
rect 28820 3238 28850 3290
rect 28850 3238 28862 3290
rect 28862 3238 28876 3290
rect 28900 3238 28914 3290
rect 28914 3238 28926 3290
rect 28926 3238 28956 3290
rect 28980 3238 28990 3290
rect 28990 3238 29036 3290
rect 28740 3236 28796 3238
rect 28820 3236 28876 3238
rect 28900 3236 28956 3238
rect 28980 3236 29036 3238
rect 28740 2202 28796 2204
rect 28820 2202 28876 2204
rect 28900 2202 28956 2204
rect 28980 2202 29036 2204
rect 28740 2150 28786 2202
rect 28786 2150 28796 2202
rect 28820 2150 28850 2202
rect 28850 2150 28862 2202
rect 28862 2150 28876 2202
rect 28900 2150 28914 2202
rect 28914 2150 28926 2202
rect 28926 2150 28956 2202
rect 28980 2150 28990 2202
rect 28990 2150 29036 2202
rect 28740 2148 28796 2150
rect 28820 2148 28876 2150
rect 28900 2148 28956 2150
rect 28980 2148 29036 2150
rect 27526 1400 27582 1456
<< metal3 >>
rect 200 49738 800 49828
rect 2957 49738 3023 49741
rect 200 49736 3023 49738
rect 200 49680 2962 49736
rect 3018 49680 3023 49736
rect 200 49678 3023 49680
rect 200 49588 800 49678
rect 2957 49675 3023 49678
rect 26601 49058 26667 49061
rect 29200 49058 29800 49148
rect 26601 49056 29800 49058
rect 26601 49000 26606 49056
rect 26662 49000 29800 49056
rect 26601 48998 29800 49000
rect 26601 48995 26667 48998
rect 29200 48908 29800 48998
rect 200 48228 800 48468
rect 29200 48228 29800 48468
rect 200 47548 800 47788
rect 28625 47698 28691 47701
rect 29200 47698 29800 47788
rect 28625 47696 29800 47698
rect 28625 47640 28630 47696
rect 28686 47640 29800 47696
rect 28625 47638 29800 47640
rect 28625 47635 28691 47638
rect 29200 47548 29800 47638
rect 4419 47360 4735 47361
rect 4419 47296 4425 47360
rect 4489 47296 4505 47360
rect 4569 47296 4585 47360
rect 4649 47296 4665 47360
rect 4729 47296 4735 47360
rect 4419 47295 4735 47296
rect 11365 47360 11681 47361
rect 11365 47296 11371 47360
rect 11435 47296 11451 47360
rect 11515 47296 11531 47360
rect 11595 47296 11611 47360
rect 11675 47296 11681 47360
rect 11365 47295 11681 47296
rect 18311 47360 18627 47361
rect 18311 47296 18317 47360
rect 18381 47296 18397 47360
rect 18461 47296 18477 47360
rect 18541 47296 18557 47360
rect 18621 47296 18627 47360
rect 18311 47295 18627 47296
rect 25257 47360 25573 47361
rect 25257 47296 25263 47360
rect 25327 47296 25343 47360
rect 25407 47296 25423 47360
rect 25487 47296 25503 47360
rect 25567 47296 25573 47360
rect 25257 47295 25573 47296
rect 200 46868 800 47108
rect 26141 47018 26207 47021
rect 29200 47018 29800 47108
rect 26141 47016 29800 47018
rect 26141 46960 26146 47016
rect 26202 46960 29800 47016
rect 26141 46958 29800 46960
rect 26141 46955 26207 46958
rect 29200 46868 29800 46958
rect 7892 46816 8208 46817
rect 7892 46752 7898 46816
rect 7962 46752 7978 46816
rect 8042 46752 8058 46816
rect 8122 46752 8138 46816
rect 8202 46752 8208 46816
rect 7892 46751 8208 46752
rect 14838 46816 15154 46817
rect 14838 46752 14844 46816
rect 14908 46752 14924 46816
rect 14988 46752 15004 46816
rect 15068 46752 15084 46816
rect 15148 46752 15154 46816
rect 14838 46751 15154 46752
rect 21784 46816 22100 46817
rect 21784 46752 21790 46816
rect 21854 46752 21870 46816
rect 21934 46752 21950 46816
rect 22014 46752 22030 46816
rect 22094 46752 22100 46816
rect 21784 46751 22100 46752
rect 28730 46816 29046 46817
rect 28730 46752 28736 46816
rect 28800 46752 28816 46816
rect 28880 46752 28896 46816
rect 28960 46752 28976 46816
rect 29040 46752 29046 46816
rect 28730 46751 29046 46752
rect 200 46188 800 46428
rect 26049 46338 26115 46341
rect 29200 46338 29800 46428
rect 26049 46336 29800 46338
rect 26049 46280 26054 46336
rect 26110 46280 29800 46336
rect 26049 46278 29800 46280
rect 26049 46275 26115 46278
rect 4419 46272 4735 46273
rect 4419 46208 4425 46272
rect 4489 46208 4505 46272
rect 4569 46208 4585 46272
rect 4649 46208 4665 46272
rect 4729 46208 4735 46272
rect 4419 46207 4735 46208
rect 11365 46272 11681 46273
rect 11365 46208 11371 46272
rect 11435 46208 11451 46272
rect 11515 46208 11531 46272
rect 11595 46208 11611 46272
rect 11675 46208 11681 46272
rect 11365 46207 11681 46208
rect 18311 46272 18627 46273
rect 18311 46208 18317 46272
rect 18381 46208 18397 46272
rect 18461 46208 18477 46272
rect 18541 46208 18557 46272
rect 18621 46208 18627 46272
rect 18311 46207 18627 46208
rect 25257 46272 25573 46273
rect 25257 46208 25263 46272
rect 25327 46208 25343 46272
rect 25407 46208 25423 46272
rect 25487 46208 25503 46272
rect 25567 46208 25573 46272
rect 25257 46207 25573 46208
rect 29200 46188 29800 46278
rect 200 45508 800 45748
rect 7892 45728 8208 45729
rect 7892 45664 7898 45728
rect 7962 45664 7978 45728
rect 8042 45664 8058 45728
rect 8122 45664 8138 45728
rect 8202 45664 8208 45728
rect 7892 45663 8208 45664
rect 14838 45728 15154 45729
rect 14838 45664 14844 45728
rect 14908 45664 14924 45728
rect 14988 45664 15004 45728
rect 15068 45664 15084 45728
rect 15148 45664 15154 45728
rect 14838 45663 15154 45664
rect 21784 45728 22100 45729
rect 21784 45664 21790 45728
rect 21854 45664 21870 45728
rect 21934 45664 21950 45728
rect 22014 45664 22030 45728
rect 22094 45664 22100 45728
rect 21784 45663 22100 45664
rect 28730 45728 29046 45729
rect 28730 45664 28736 45728
rect 28800 45664 28816 45728
rect 28880 45664 28896 45728
rect 28960 45664 28976 45728
rect 29040 45664 29046 45728
rect 28730 45663 29046 45664
rect 29200 45508 29800 45748
rect 4419 45184 4735 45185
rect 4419 45120 4425 45184
rect 4489 45120 4505 45184
rect 4569 45120 4585 45184
rect 4649 45120 4665 45184
rect 4729 45120 4735 45184
rect 4419 45119 4735 45120
rect 11365 45184 11681 45185
rect 11365 45120 11371 45184
rect 11435 45120 11451 45184
rect 11515 45120 11531 45184
rect 11595 45120 11611 45184
rect 11675 45120 11681 45184
rect 11365 45119 11681 45120
rect 18311 45184 18627 45185
rect 18311 45120 18317 45184
rect 18381 45120 18397 45184
rect 18461 45120 18477 45184
rect 18541 45120 18557 45184
rect 18621 45120 18627 45184
rect 18311 45119 18627 45120
rect 25257 45184 25573 45185
rect 25257 45120 25263 45184
rect 25327 45120 25343 45184
rect 25407 45120 25423 45184
rect 25487 45120 25503 45184
rect 25567 45120 25573 45184
rect 25257 45119 25573 45120
rect 200 44978 800 45068
rect 4245 44978 4311 44981
rect 200 44976 4311 44978
rect 200 44920 4250 44976
rect 4306 44920 4311 44976
rect 200 44918 4311 44920
rect 200 44828 800 44918
rect 4245 44915 4311 44918
rect 28349 44978 28415 44981
rect 29200 44978 29800 45068
rect 28349 44976 29800 44978
rect 28349 44920 28354 44976
rect 28410 44920 29800 44976
rect 28349 44918 29800 44920
rect 28349 44915 28415 44918
rect 29200 44828 29800 44918
rect 7892 44640 8208 44641
rect 7892 44576 7898 44640
rect 7962 44576 7978 44640
rect 8042 44576 8058 44640
rect 8122 44576 8138 44640
rect 8202 44576 8208 44640
rect 7892 44575 8208 44576
rect 14838 44640 15154 44641
rect 14838 44576 14844 44640
rect 14908 44576 14924 44640
rect 14988 44576 15004 44640
rect 15068 44576 15084 44640
rect 15148 44576 15154 44640
rect 14838 44575 15154 44576
rect 21784 44640 22100 44641
rect 21784 44576 21790 44640
rect 21854 44576 21870 44640
rect 21934 44576 21950 44640
rect 22014 44576 22030 44640
rect 22094 44576 22100 44640
rect 21784 44575 22100 44576
rect 28730 44640 29046 44641
rect 28730 44576 28736 44640
rect 28800 44576 28816 44640
rect 28880 44576 28896 44640
rect 28960 44576 28976 44640
rect 29040 44576 29046 44640
rect 28730 44575 29046 44576
rect 200 44298 800 44388
rect 3601 44298 3667 44301
rect 200 44296 3667 44298
rect 200 44240 3606 44296
rect 3662 44240 3667 44296
rect 200 44238 3667 44240
rect 200 44148 800 44238
rect 3601 44235 3667 44238
rect 4419 44096 4735 44097
rect 4419 44032 4425 44096
rect 4489 44032 4505 44096
rect 4569 44032 4585 44096
rect 4649 44032 4665 44096
rect 4729 44032 4735 44096
rect 4419 44031 4735 44032
rect 11365 44096 11681 44097
rect 11365 44032 11371 44096
rect 11435 44032 11451 44096
rect 11515 44032 11531 44096
rect 11595 44032 11611 44096
rect 11675 44032 11681 44096
rect 11365 44031 11681 44032
rect 18311 44096 18627 44097
rect 18311 44032 18317 44096
rect 18381 44032 18397 44096
rect 18461 44032 18477 44096
rect 18541 44032 18557 44096
rect 18621 44032 18627 44096
rect 18311 44031 18627 44032
rect 25257 44096 25573 44097
rect 25257 44032 25263 44096
rect 25327 44032 25343 44096
rect 25407 44032 25423 44096
rect 25487 44032 25503 44096
rect 25567 44032 25573 44096
rect 25257 44031 25573 44032
rect 7892 43552 8208 43553
rect 7892 43488 7898 43552
rect 7962 43488 7978 43552
rect 8042 43488 8058 43552
rect 8122 43488 8138 43552
rect 8202 43488 8208 43552
rect 7892 43487 8208 43488
rect 14838 43552 15154 43553
rect 14838 43488 14844 43552
rect 14908 43488 14924 43552
rect 14988 43488 15004 43552
rect 15068 43488 15084 43552
rect 15148 43488 15154 43552
rect 14838 43487 15154 43488
rect 21784 43552 22100 43553
rect 21784 43488 21790 43552
rect 21854 43488 21870 43552
rect 21934 43488 21950 43552
rect 22014 43488 22030 43552
rect 22094 43488 22100 43552
rect 21784 43487 22100 43488
rect 28730 43552 29046 43553
rect 28730 43488 28736 43552
rect 28800 43488 28816 43552
rect 28880 43488 28896 43552
rect 28960 43488 28976 43552
rect 29040 43488 29046 43552
rect 28730 43487 29046 43488
rect 29200 43468 29800 43708
rect 200 42788 800 43028
rect 4419 43008 4735 43009
rect 4419 42944 4425 43008
rect 4489 42944 4505 43008
rect 4569 42944 4585 43008
rect 4649 42944 4665 43008
rect 4729 42944 4735 43008
rect 4419 42943 4735 42944
rect 11365 43008 11681 43009
rect 11365 42944 11371 43008
rect 11435 42944 11451 43008
rect 11515 42944 11531 43008
rect 11595 42944 11611 43008
rect 11675 42944 11681 43008
rect 11365 42943 11681 42944
rect 18311 43008 18627 43009
rect 18311 42944 18317 43008
rect 18381 42944 18397 43008
rect 18461 42944 18477 43008
rect 18541 42944 18557 43008
rect 18621 42944 18627 43008
rect 18311 42943 18627 42944
rect 25257 43008 25573 43009
rect 25257 42944 25263 43008
rect 25327 42944 25343 43008
rect 25407 42944 25423 43008
rect 25487 42944 25503 43008
rect 25567 42944 25573 43008
rect 25257 42943 25573 42944
rect 26049 42938 26115 42941
rect 29200 42938 29800 43028
rect 26049 42936 29800 42938
rect 26049 42880 26054 42936
rect 26110 42880 29800 42936
rect 26049 42878 29800 42880
rect 26049 42875 26115 42878
rect 29200 42788 29800 42878
rect 7892 42464 8208 42465
rect 7892 42400 7898 42464
rect 7962 42400 7978 42464
rect 8042 42400 8058 42464
rect 8122 42400 8138 42464
rect 8202 42400 8208 42464
rect 7892 42399 8208 42400
rect 14838 42464 15154 42465
rect 14838 42400 14844 42464
rect 14908 42400 14924 42464
rect 14988 42400 15004 42464
rect 15068 42400 15084 42464
rect 15148 42400 15154 42464
rect 14838 42399 15154 42400
rect 21784 42464 22100 42465
rect 21784 42400 21790 42464
rect 21854 42400 21870 42464
rect 21934 42400 21950 42464
rect 22014 42400 22030 42464
rect 22094 42400 22100 42464
rect 21784 42399 22100 42400
rect 28730 42464 29046 42465
rect 28730 42400 28736 42464
rect 28800 42400 28816 42464
rect 28880 42400 28896 42464
rect 28960 42400 28976 42464
rect 29040 42400 29046 42464
rect 28730 42399 29046 42400
rect 200 42258 800 42348
rect 1577 42258 1643 42261
rect 200 42256 1643 42258
rect 200 42200 1582 42256
rect 1638 42200 1643 42256
rect 200 42198 1643 42200
rect 200 42108 800 42198
rect 1577 42195 1643 42198
rect 27429 42258 27495 42261
rect 29200 42258 29800 42348
rect 27429 42256 29800 42258
rect 27429 42200 27434 42256
rect 27490 42200 29800 42256
rect 27429 42198 29800 42200
rect 27429 42195 27495 42198
rect 29200 42108 29800 42198
rect 4419 41920 4735 41921
rect 4419 41856 4425 41920
rect 4489 41856 4505 41920
rect 4569 41856 4585 41920
rect 4649 41856 4665 41920
rect 4729 41856 4735 41920
rect 4419 41855 4735 41856
rect 11365 41920 11681 41921
rect 11365 41856 11371 41920
rect 11435 41856 11451 41920
rect 11515 41856 11531 41920
rect 11595 41856 11611 41920
rect 11675 41856 11681 41920
rect 11365 41855 11681 41856
rect 18311 41920 18627 41921
rect 18311 41856 18317 41920
rect 18381 41856 18397 41920
rect 18461 41856 18477 41920
rect 18541 41856 18557 41920
rect 18621 41856 18627 41920
rect 18311 41855 18627 41856
rect 25257 41920 25573 41921
rect 25257 41856 25263 41920
rect 25327 41856 25343 41920
rect 25407 41856 25423 41920
rect 25487 41856 25503 41920
rect 25567 41856 25573 41920
rect 25257 41855 25573 41856
rect 200 41578 800 41668
rect 2773 41578 2839 41581
rect 200 41576 2839 41578
rect 200 41520 2778 41576
rect 2834 41520 2839 41576
rect 200 41518 2839 41520
rect 200 41428 800 41518
rect 2773 41515 2839 41518
rect 26141 41578 26207 41581
rect 29200 41578 29800 41668
rect 26141 41576 29800 41578
rect 26141 41520 26146 41576
rect 26202 41520 29800 41576
rect 26141 41518 29800 41520
rect 26141 41515 26207 41518
rect 29200 41428 29800 41518
rect 7892 41376 8208 41377
rect 7892 41312 7898 41376
rect 7962 41312 7978 41376
rect 8042 41312 8058 41376
rect 8122 41312 8138 41376
rect 8202 41312 8208 41376
rect 7892 41311 8208 41312
rect 14838 41376 15154 41377
rect 14838 41312 14844 41376
rect 14908 41312 14924 41376
rect 14988 41312 15004 41376
rect 15068 41312 15084 41376
rect 15148 41312 15154 41376
rect 14838 41311 15154 41312
rect 21784 41376 22100 41377
rect 21784 41312 21790 41376
rect 21854 41312 21870 41376
rect 21934 41312 21950 41376
rect 22014 41312 22030 41376
rect 22094 41312 22100 41376
rect 21784 41311 22100 41312
rect 28730 41376 29046 41377
rect 28730 41312 28736 41376
rect 28800 41312 28816 41376
rect 28880 41312 28896 41376
rect 28960 41312 28976 41376
rect 29040 41312 29046 41376
rect 28730 41311 29046 41312
rect 200 40748 800 40988
rect 27521 40898 27587 40901
rect 29200 40898 29800 40988
rect 27521 40896 29800 40898
rect 27521 40840 27526 40896
rect 27582 40840 29800 40896
rect 27521 40838 29800 40840
rect 27521 40835 27587 40838
rect 4419 40832 4735 40833
rect 4419 40768 4425 40832
rect 4489 40768 4505 40832
rect 4569 40768 4585 40832
rect 4649 40768 4665 40832
rect 4729 40768 4735 40832
rect 4419 40767 4735 40768
rect 11365 40832 11681 40833
rect 11365 40768 11371 40832
rect 11435 40768 11451 40832
rect 11515 40768 11531 40832
rect 11595 40768 11611 40832
rect 11675 40768 11681 40832
rect 11365 40767 11681 40768
rect 18311 40832 18627 40833
rect 18311 40768 18317 40832
rect 18381 40768 18397 40832
rect 18461 40768 18477 40832
rect 18541 40768 18557 40832
rect 18621 40768 18627 40832
rect 18311 40767 18627 40768
rect 25257 40832 25573 40833
rect 25257 40768 25263 40832
rect 25327 40768 25343 40832
rect 25407 40768 25423 40832
rect 25487 40768 25503 40832
rect 25567 40768 25573 40832
rect 25257 40767 25573 40768
rect 29200 40748 29800 40838
rect 200 40068 800 40308
rect 7892 40288 8208 40289
rect 7892 40224 7898 40288
rect 7962 40224 7978 40288
rect 8042 40224 8058 40288
rect 8122 40224 8138 40288
rect 8202 40224 8208 40288
rect 7892 40223 8208 40224
rect 14838 40288 15154 40289
rect 14838 40224 14844 40288
rect 14908 40224 14924 40288
rect 14988 40224 15004 40288
rect 15068 40224 15084 40288
rect 15148 40224 15154 40288
rect 14838 40223 15154 40224
rect 21784 40288 22100 40289
rect 21784 40224 21790 40288
rect 21854 40224 21870 40288
rect 21934 40224 21950 40288
rect 22014 40224 22030 40288
rect 22094 40224 22100 40288
rect 21784 40223 22100 40224
rect 28730 40288 29046 40289
rect 28730 40224 28736 40288
rect 28800 40224 28816 40288
rect 28880 40224 28896 40288
rect 28960 40224 28976 40288
rect 29040 40224 29046 40288
rect 28730 40223 29046 40224
rect 29200 40218 29800 40308
rect 29913 40218 29979 40221
rect 29200 40216 29979 40218
rect 29200 40160 29918 40216
rect 29974 40160 29979 40216
rect 29200 40158 29979 40160
rect 29200 40068 29800 40158
rect 29913 40155 29979 40158
rect 4419 39744 4735 39745
rect 4419 39680 4425 39744
rect 4489 39680 4505 39744
rect 4569 39680 4585 39744
rect 4649 39680 4665 39744
rect 4729 39680 4735 39744
rect 4419 39679 4735 39680
rect 11365 39744 11681 39745
rect 11365 39680 11371 39744
rect 11435 39680 11451 39744
rect 11515 39680 11531 39744
rect 11595 39680 11611 39744
rect 11675 39680 11681 39744
rect 11365 39679 11681 39680
rect 18311 39744 18627 39745
rect 18311 39680 18317 39744
rect 18381 39680 18397 39744
rect 18461 39680 18477 39744
rect 18541 39680 18557 39744
rect 18621 39680 18627 39744
rect 18311 39679 18627 39680
rect 25257 39744 25573 39745
rect 25257 39680 25263 39744
rect 25327 39680 25343 39744
rect 25407 39680 25423 39744
rect 25487 39680 25503 39744
rect 25567 39680 25573 39744
rect 25257 39679 25573 39680
rect 200 39388 800 39628
rect 28625 39538 28691 39541
rect 29200 39538 29800 39628
rect 28625 39536 29800 39538
rect 28625 39480 28630 39536
rect 28686 39480 29800 39536
rect 28625 39478 29800 39480
rect 28625 39475 28691 39478
rect 29200 39388 29800 39478
rect 7892 39200 8208 39201
rect 7892 39136 7898 39200
rect 7962 39136 7978 39200
rect 8042 39136 8058 39200
rect 8122 39136 8138 39200
rect 8202 39136 8208 39200
rect 7892 39135 8208 39136
rect 14838 39200 15154 39201
rect 14838 39136 14844 39200
rect 14908 39136 14924 39200
rect 14988 39136 15004 39200
rect 15068 39136 15084 39200
rect 15148 39136 15154 39200
rect 14838 39135 15154 39136
rect 21784 39200 22100 39201
rect 21784 39136 21790 39200
rect 21854 39136 21870 39200
rect 21934 39136 21950 39200
rect 22014 39136 22030 39200
rect 22094 39136 22100 39200
rect 21784 39135 22100 39136
rect 28730 39200 29046 39201
rect 28730 39136 28736 39200
rect 28800 39136 28816 39200
rect 28880 39136 28896 39200
rect 28960 39136 28976 39200
rect 29040 39136 29046 39200
rect 28730 39135 29046 39136
rect 200 38858 800 38948
rect 2773 38858 2839 38861
rect 200 38856 2839 38858
rect 200 38800 2778 38856
rect 2834 38800 2839 38856
rect 200 38798 2839 38800
rect 200 38708 800 38798
rect 2773 38795 2839 38798
rect 4419 38656 4735 38657
rect 4419 38592 4425 38656
rect 4489 38592 4505 38656
rect 4569 38592 4585 38656
rect 4649 38592 4665 38656
rect 4729 38592 4735 38656
rect 4419 38591 4735 38592
rect 11365 38656 11681 38657
rect 11365 38592 11371 38656
rect 11435 38592 11451 38656
rect 11515 38592 11531 38656
rect 11595 38592 11611 38656
rect 11675 38592 11681 38656
rect 11365 38591 11681 38592
rect 18311 38656 18627 38657
rect 18311 38592 18317 38656
rect 18381 38592 18397 38656
rect 18461 38592 18477 38656
rect 18541 38592 18557 38656
rect 18621 38592 18627 38656
rect 18311 38591 18627 38592
rect 25257 38656 25573 38657
rect 25257 38592 25263 38656
rect 25327 38592 25343 38656
rect 25407 38592 25423 38656
rect 25487 38592 25503 38656
rect 25567 38592 25573 38656
rect 25257 38591 25573 38592
rect 19517 38450 19583 38453
rect 20621 38450 20687 38453
rect 26601 38450 26667 38453
rect 19517 38448 26667 38450
rect 19517 38392 19522 38448
rect 19578 38392 20626 38448
rect 20682 38392 26606 38448
rect 26662 38392 26667 38448
rect 19517 38390 26667 38392
rect 19517 38387 19583 38390
rect 20621 38387 20687 38390
rect 26601 38387 26667 38390
rect 7892 38112 8208 38113
rect 7892 38048 7898 38112
rect 7962 38048 7978 38112
rect 8042 38048 8058 38112
rect 8122 38048 8138 38112
rect 8202 38048 8208 38112
rect 7892 38047 8208 38048
rect 14838 38112 15154 38113
rect 14838 38048 14844 38112
rect 14908 38048 14924 38112
rect 14988 38048 15004 38112
rect 15068 38048 15084 38112
rect 15148 38048 15154 38112
rect 14838 38047 15154 38048
rect 21784 38112 22100 38113
rect 21784 38048 21790 38112
rect 21854 38048 21870 38112
rect 21934 38048 21950 38112
rect 22014 38048 22030 38112
rect 22094 38048 22100 38112
rect 21784 38047 22100 38048
rect 28730 38112 29046 38113
rect 28730 38048 28736 38112
rect 28800 38048 28816 38112
rect 28880 38048 28896 38112
rect 28960 38048 28976 38112
rect 29040 38048 29046 38112
rect 28730 38047 29046 38048
rect 29200 38028 29800 38268
rect 200 37498 800 37588
rect 4419 37568 4735 37569
rect 4419 37504 4425 37568
rect 4489 37504 4505 37568
rect 4569 37504 4585 37568
rect 4649 37504 4665 37568
rect 4729 37504 4735 37568
rect 4419 37503 4735 37504
rect 11365 37568 11681 37569
rect 11365 37504 11371 37568
rect 11435 37504 11451 37568
rect 11515 37504 11531 37568
rect 11595 37504 11611 37568
rect 11675 37504 11681 37568
rect 11365 37503 11681 37504
rect 18311 37568 18627 37569
rect 18311 37504 18317 37568
rect 18381 37504 18397 37568
rect 18461 37504 18477 37568
rect 18541 37504 18557 37568
rect 18621 37504 18627 37568
rect 18311 37503 18627 37504
rect 25257 37568 25573 37569
rect 25257 37504 25263 37568
rect 25327 37504 25343 37568
rect 25407 37504 25423 37568
rect 25487 37504 25503 37568
rect 25567 37504 25573 37568
rect 25257 37503 25573 37504
rect 1669 37498 1735 37501
rect 200 37496 1735 37498
rect 200 37440 1674 37496
rect 1730 37440 1735 37496
rect 200 37438 1735 37440
rect 200 37348 800 37438
rect 1669 37435 1735 37438
rect 29200 37348 29800 37588
rect 7892 37024 8208 37025
rect 7892 36960 7898 37024
rect 7962 36960 7978 37024
rect 8042 36960 8058 37024
rect 8122 36960 8138 37024
rect 8202 36960 8208 37024
rect 7892 36959 8208 36960
rect 14838 37024 15154 37025
rect 14838 36960 14844 37024
rect 14908 36960 14924 37024
rect 14988 36960 15004 37024
rect 15068 36960 15084 37024
rect 15148 36960 15154 37024
rect 14838 36959 15154 36960
rect 21784 37024 22100 37025
rect 21784 36960 21790 37024
rect 21854 36960 21870 37024
rect 21934 36960 21950 37024
rect 22014 36960 22030 37024
rect 22094 36960 22100 37024
rect 21784 36959 22100 36960
rect 28730 37024 29046 37025
rect 28730 36960 28736 37024
rect 28800 36960 28816 37024
rect 28880 36960 28896 37024
rect 28960 36960 28976 37024
rect 29040 36960 29046 37024
rect 28730 36959 29046 36960
rect 200 36818 800 36908
rect 2865 36818 2931 36821
rect 200 36816 2931 36818
rect 200 36760 2870 36816
rect 2926 36760 2931 36816
rect 200 36758 2931 36760
rect 200 36668 800 36758
rect 2865 36755 2931 36758
rect 27337 36818 27403 36821
rect 29200 36818 29800 36908
rect 27337 36816 29800 36818
rect 27337 36760 27342 36816
rect 27398 36760 29800 36816
rect 27337 36758 29800 36760
rect 27337 36755 27403 36758
rect 29200 36668 29800 36758
rect 4419 36480 4735 36481
rect 4419 36416 4425 36480
rect 4489 36416 4505 36480
rect 4569 36416 4585 36480
rect 4649 36416 4665 36480
rect 4729 36416 4735 36480
rect 4419 36415 4735 36416
rect 11365 36480 11681 36481
rect 11365 36416 11371 36480
rect 11435 36416 11451 36480
rect 11515 36416 11531 36480
rect 11595 36416 11611 36480
rect 11675 36416 11681 36480
rect 11365 36415 11681 36416
rect 18311 36480 18627 36481
rect 18311 36416 18317 36480
rect 18381 36416 18397 36480
rect 18461 36416 18477 36480
rect 18541 36416 18557 36480
rect 18621 36416 18627 36480
rect 18311 36415 18627 36416
rect 25257 36480 25573 36481
rect 25257 36416 25263 36480
rect 25327 36416 25343 36480
rect 25407 36416 25423 36480
rect 25487 36416 25503 36480
rect 25567 36416 25573 36480
rect 25257 36415 25573 36416
rect 200 36138 800 36228
rect 1669 36138 1735 36141
rect 200 36136 1735 36138
rect 200 36080 1674 36136
rect 1730 36080 1735 36136
rect 200 36078 1735 36080
rect 200 35988 800 36078
rect 1669 36075 1735 36078
rect 26141 36138 26207 36141
rect 29200 36138 29800 36228
rect 26141 36136 29800 36138
rect 26141 36080 26146 36136
rect 26202 36080 29800 36136
rect 26141 36078 29800 36080
rect 26141 36075 26207 36078
rect 29200 35988 29800 36078
rect 7892 35936 8208 35937
rect 7892 35872 7898 35936
rect 7962 35872 7978 35936
rect 8042 35872 8058 35936
rect 8122 35872 8138 35936
rect 8202 35872 8208 35936
rect 7892 35871 8208 35872
rect 14838 35936 15154 35937
rect 14838 35872 14844 35936
rect 14908 35872 14924 35936
rect 14988 35872 15004 35936
rect 15068 35872 15084 35936
rect 15148 35872 15154 35936
rect 14838 35871 15154 35872
rect 21784 35936 22100 35937
rect 21784 35872 21790 35936
rect 21854 35872 21870 35936
rect 21934 35872 21950 35936
rect 22014 35872 22030 35936
rect 22094 35872 22100 35936
rect 21784 35871 22100 35872
rect 28730 35936 29046 35937
rect 28730 35872 28736 35936
rect 28800 35872 28816 35936
rect 28880 35872 28896 35936
rect 28960 35872 28976 35936
rect 29040 35872 29046 35936
rect 28730 35871 29046 35872
rect 200 35308 800 35548
rect 4419 35392 4735 35393
rect 4419 35328 4425 35392
rect 4489 35328 4505 35392
rect 4569 35328 4585 35392
rect 4649 35328 4665 35392
rect 4729 35328 4735 35392
rect 4419 35327 4735 35328
rect 11365 35392 11681 35393
rect 11365 35328 11371 35392
rect 11435 35328 11451 35392
rect 11515 35328 11531 35392
rect 11595 35328 11611 35392
rect 11675 35328 11681 35392
rect 11365 35327 11681 35328
rect 18311 35392 18627 35393
rect 18311 35328 18317 35392
rect 18381 35328 18397 35392
rect 18461 35328 18477 35392
rect 18541 35328 18557 35392
rect 18621 35328 18627 35392
rect 18311 35327 18627 35328
rect 25257 35392 25573 35393
rect 25257 35328 25263 35392
rect 25327 35328 25343 35392
rect 25407 35328 25423 35392
rect 25487 35328 25503 35392
rect 25567 35328 25573 35392
rect 25257 35327 25573 35328
rect 29200 35308 29800 35548
rect 200 34778 800 34868
rect 7892 34848 8208 34849
rect 7892 34784 7898 34848
rect 7962 34784 7978 34848
rect 8042 34784 8058 34848
rect 8122 34784 8138 34848
rect 8202 34784 8208 34848
rect 7892 34783 8208 34784
rect 14838 34848 15154 34849
rect 14838 34784 14844 34848
rect 14908 34784 14924 34848
rect 14988 34784 15004 34848
rect 15068 34784 15084 34848
rect 15148 34784 15154 34848
rect 14838 34783 15154 34784
rect 21784 34848 22100 34849
rect 21784 34784 21790 34848
rect 21854 34784 21870 34848
rect 21934 34784 21950 34848
rect 22014 34784 22030 34848
rect 22094 34784 22100 34848
rect 21784 34783 22100 34784
rect 28730 34848 29046 34849
rect 28730 34784 28736 34848
rect 28800 34784 28816 34848
rect 28880 34784 28896 34848
rect 28960 34784 28976 34848
rect 29040 34784 29046 34848
rect 28730 34783 29046 34784
rect 2773 34778 2839 34781
rect 200 34776 2839 34778
rect 200 34720 2778 34776
rect 2834 34720 2839 34776
rect 200 34718 2839 34720
rect 200 34628 800 34718
rect 2773 34715 2839 34718
rect 29200 34628 29800 34868
rect 4419 34304 4735 34305
rect 4419 34240 4425 34304
rect 4489 34240 4505 34304
rect 4569 34240 4585 34304
rect 4649 34240 4665 34304
rect 4729 34240 4735 34304
rect 4419 34239 4735 34240
rect 11365 34304 11681 34305
rect 11365 34240 11371 34304
rect 11435 34240 11451 34304
rect 11515 34240 11531 34304
rect 11595 34240 11611 34304
rect 11675 34240 11681 34304
rect 11365 34239 11681 34240
rect 18311 34304 18627 34305
rect 18311 34240 18317 34304
rect 18381 34240 18397 34304
rect 18461 34240 18477 34304
rect 18541 34240 18557 34304
rect 18621 34240 18627 34304
rect 18311 34239 18627 34240
rect 25257 34304 25573 34305
rect 25257 34240 25263 34304
rect 25327 34240 25343 34304
rect 25407 34240 25423 34304
rect 25487 34240 25503 34304
rect 25567 34240 25573 34304
rect 25257 34239 25573 34240
rect 200 33948 800 34188
rect 27521 34098 27587 34101
rect 29200 34098 29800 34188
rect 27521 34096 29800 34098
rect 27521 34040 27526 34096
rect 27582 34040 29800 34096
rect 27521 34038 29800 34040
rect 27521 34035 27587 34038
rect 29200 33948 29800 34038
rect 7892 33760 8208 33761
rect 7892 33696 7898 33760
rect 7962 33696 7978 33760
rect 8042 33696 8058 33760
rect 8122 33696 8138 33760
rect 8202 33696 8208 33760
rect 7892 33695 8208 33696
rect 14838 33760 15154 33761
rect 14838 33696 14844 33760
rect 14908 33696 14924 33760
rect 14988 33696 15004 33760
rect 15068 33696 15084 33760
rect 15148 33696 15154 33760
rect 14838 33695 15154 33696
rect 21784 33760 22100 33761
rect 21784 33696 21790 33760
rect 21854 33696 21870 33760
rect 21934 33696 21950 33760
rect 22014 33696 22030 33760
rect 22094 33696 22100 33760
rect 21784 33695 22100 33696
rect 28730 33760 29046 33761
rect 28730 33696 28736 33760
rect 28800 33696 28816 33760
rect 28880 33696 28896 33760
rect 28960 33696 28976 33760
rect 29040 33696 29046 33760
rect 28730 33695 29046 33696
rect 200 33418 800 33508
rect 3509 33418 3575 33421
rect 200 33416 3575 33418
rect 200 33360 3514 33416
rect 3570 33360 3575 33416
rect 200 33358 3575 33360
rect 200 33268 800 33358
rect 3509 33355 3575 33358
rect 4419 33216 4735 33217
rect 4419 33152 4425 33216
rect 4489 33152 4505 33216
rect 4569 33152 4585 33216
rect 4649 33152 4665 33216
rect 4729 33152 4735 33216
rect 4419 33151 4735 33152
rect 11365 33216 11681 33217
rect 11365 33152 11371 33216
rect 11435 33152 11451 33216
rect 11515 33152 11531 33216
rect 11595 33152 11611 33216
rect 11675 33152 11681 33216
rect 11365 33151 11681 33152
rect 18311 33216 18627 33217
rect 18311 33152 18317 33216
rect 18381 33152 18397 33216
rect 18461 33152 18477 33216
rect 18541 33152 18557 33216
rect 18621 33152 18627 33216
rect 18311 33151 18627 33152
rect 25257 33216 25573 33217
rect 25257 33152 25263 33216
rect 25327 33152 25343 33216
rect 25407 33152 25423 33216
rect 25487 33152 25503 33216
rect 25567 33152 25573 33216
rect 25257 33151 25573 33152
rect 29200 32738 29800 32828
rect 29200 32678 29930 32738
rect 7892 32672 8208 32673
rect 7892 32608 7898 32672
rect 7962 32608 7978 32672
rect 8042 32608 8058 32672
rect 8122 32608 8138 32672
rect 8202 32608 8208 32672
rect 7892 32607 8208 32608
rect 14838 32672 15154 32673
rect 14838 32608 14844 32672
rect 14908 32608 14924 32672
rect 14988 32608 15004 32672
rect 15068 32608 15084 32672
rect 15148 32608 15154 32672
rect 14838 32607 15154 32608
rect 21784 32672 22100 32673
rect 21784 32608 21790 32672
rect 21854 32608 21870 32672
rect 21934 32608 21950 32672
rect 22014 32608 22030 32672
rect 22094 32608 22100 32672
rect 21784 32607 22100 32608
rect 28730 32672 29046 32673
rect 28730 32608 28736 32672
rect 28800 32608 28816 32672
rect 28880 32608 28896 32672
rect 28960 32608 28976 32672
rect 29040 32608 29046 32672
rect 28730 32607 29046 32608
rect 29200 32602 29800 32678
rect 29870 32602 29930 32678
rect 29200 32588 29930 32602
rect 29318 32542 29930 32588
rect 27429 32330 27495 32333
rect 29318 32330 29378 32542
rect 27429 32328 29378 32330
rect 27429 32272 27434 32328
rect 27490 32272 29378 32328
rect 27429 32270 29378 32272
rect 27429 32267 27495 32270
rect 200 32058 800 32148
rect 4419 32128 4735 32129
rect 4419 32064 4425 32128
rect 4489 32064 4505 32128
rect 4569 32064 4585 32128
rect 4649 32064 4665 32128
rect 4729 32064 4735 32128
rect 4419 32063 4735 32064
rect 11365 32128 11681 32129
rect 11365 32064 11371 32128
rect 11435 32064 11451 32128
rect 11515 32064 11531 32128
rect 11595 32064 11611 32128
rect 11675 32064 11681 32128
rect 11365 32063 11681 32064
rect 18311 32128 18627 32129
rect 18311 32064 18317 32128
rect 18381 32064 18397 32128
rect 18461 32064 18477 32128
rect 18541 32064 18557 32128
rect 18621 32064 18627 32128
rect 18311 32063 18627 32064
rect 25257 32128 25573 32129
rect 25257 32064 25263 32128
rect 25327 32064 25343 32128
rect 25407 32064 25423 32128
rect 25487 32064 25503 32128
rect 25567 32064 25573 32128
rect 25257 32063 25573 32064
rect 2773 32058 2839 32061
rect 200 32056 2839 32058
rect 200 32000 2778 32056
rect 2834 32000 2839 32056
rect 200 31998 2839 32000
rect 200 31908 800 31998
rect 2773 31995 2839 31998
rect 28349 32058 28415 32061
rect 29200 32058 29800 32148
rect 28349 32056 29800 32058
rect 28349 32000 28354 32056
rect 28410 32000 29800 32056
rect 28349 31998 29800 32000
rect 28349 31995 28415 31998
rect 29200 31908 29800 31998
rect 7892 31584 8208 31585
rect 7892 31520 7898 31584
rect 7962 31520 7978 31584
rect 8042 31520 8058 31584
rect 8122 31520 8138 31584
rect 8202 31520 8208 31584
rect 7892 31519 8208 31520
rect 14838 31584 15154 31585
rect 14838 31520 14844 31584
rect 14908 31520 14924 31584
rect 14988 31520 15004 31584
rect 15068 31520 15084 31584
rect 15148 31520 15154 31584
rect 14838 31519 15154 31520
rect 21784 31584 22100 31585
rect 21784 31520 21790 31584
rect 21854 31520 21870 31584
rect 21934 31520 21950 31584
rect 22014 31520 22030 31584
rect 22094 31520 22100 31584
rect 21784 31519 22100 31520
rect 28730 31584 29046 31585
rect 28730 31520 28736 31584
rect 28800 31520 28816 31584
rect 28880 31520 28896 31584
rect 28960 31520 28976 31584
rect 29040 31520 29046 31584
rect 28730 31519 29046 31520
rect 200 31228 800 31468
rect 26141 31378 26207 31381
rect 29200 31378 29800 31468
rect 26141 31376 29800 31378
rect 26141 31320 26146 31376
rect 26202 31320 29800 31376
rect 26141 31318 29800 31320
rect 26141 31315 26207 31318
rect 29200 31228 29800 31318
rect 4419 31040 4735 31041
rect 4419 30976 4425 31040
rect 4489 30976 4505 31040
rect 4569 30976 4585 31040
rect 4649 30976 4665 31040
rect 4729 30976 4735 31040
rect 4419 30975 4735 30976
rect 11365 31040 11681 31041
rect 11365 30976 11371 31040
rect 11435 30976 11451 31040
rect 11515 30976 11531 31040
rect 11595 30976 11611 31040
rect 11675 30976 11681 31040
rect 11365 30975 11681 30976
rect 18311 31040 18627 31041
rect 18311 30976 18317 31040
rect 18381 30976 18397 31040
rect 18461 30976 18477 31040
rect 18541 30976 18557 31040
rect 18621 30976 18627 31040
rect 18311 30975 18627 30976
rect 25257 31040 25573 31041
rect 25257 30976 25263 31040
rect 25327 30976 25343 31040
rect 25407 30976 25423 31040
rect 25487 30976 25503 31040
rect 25567 30976 25573 31040
rect 25257 30975 25573 30976
rect 200 30548 800 30788
rect 27521 30698 27587 30701
rect 29200 30698 29800 30788
rect 27521 30696 29800 30698
rect 27521 30640 27526 30696
rect 27582 30640 29800 30696
rect 27521 30638 29800 30640
rect 27521 30635 27587 30638
rect 29200 30548 29800 30638
rect 7892 30496 8208 30497
rect 7892 30432 7898 30496
rect 7962 30432 7978 30496
rect 8042 30432 8058 30496
rect 8122 30432 8138 30496
rect 8202 30432 8208 30496
rect 7892 30431 8208 30432
rect 14838 30496 15154 30497
rect 14838 30432 14844 30496
rect 14908 30432 14924 30496
rect 14988 30432 15004 30496
rect 15068 30432 15084 30496
rect 15148 30432 15154 30496
rect 14838 30431 15154 30432
rect 21784 30496 22100 30497
rect 21784 30432 21790 30496
rect 21854 30432 21870 30496
rect 21934 30432 21950 30496
rect 22014 30432 22030 30496
rect 22094 30432 22100 30496
rect 21784 30431 22100 30432
rect 28730 30496 29046 30497
rect 28730 30432 28736 30496
rect 28800 30432 28816 30496
rect 28880 30432 28896 30496
rect 28960 30432 28976 30496
rect 29040 30432 29046 30496
rect 28730 30431 29046 30432
rect 200 30018 800 30108
rect 1577 30018 1643 30021
rect 200 30016 1643 30018
rect 200 29960 1582 30016
rect 1638 29960 1643 30016
rect 200 29958 1643 29960
rect 200 29868 800 29958
rect 1577 29955 1643 29958
rect 26601 30018 26667 30021
rect 29200 30018 29800 30108
rect 26601 30016 29800 30018
rect 26601 29960 26606 30016
rect 26662 29960 29800 30016
rect 26601 29958 29800 29960
rect 26601 29955 26667 29958
rect 4419 29952 4735 29953
rect 4419 29888 4425 29952
rect 4489 29888 4505 29952
rect 4569 29888 4585 29952
rect 4649 29888 4665 29952
rect 4729 29888 4735 29952
rect 4419 29887 4735 29888
rect 11365 29952 11681 29953
rect 11365 29888 11371 29952
rect 11435 29888 11451 29952
rect 11515 29888 11531 29952
rect 11595 29888 11611 29952
rect 11675 29888 11681 29952
rect 11365 29887 11681 29888
rect 18311 29952 18627 29953
rect 18311 29888 18317 29952
rect 18381 29888 18397 29952
rect 18461 29888 18477 29952
rect 18541 29888 18557 29952
rect 18621 29888 18627 29952
rect 18311 29887 18627 29888
rect 25257 29952 25573 29953
rect 25257 29888 25263 29952
rect 25327 29888 25343 29952
rect 25407 29888 25423 29952
rect 25487 29888 25503 29952
rect 25567 29888 25573 29952
rect 25257 29887 25573 29888
rect 29200 29868 29800 29958
rect 200 29188 800 29428
rect 7892 29408 8208 29409
rect 7892 29344 7898 29408
rect 7962 29344 7978 29408
rect 8042 29344 8058 29408
rect 8122 29344 8138 29408
rect 8202 29344 8208 29408
rect 7892 29343 8208 29344
rect 14838 29408 15154 29409
rect 14838 29344 14844 29408
rect 14908 29344 14924 29408
rect 14988 29344 15004 29408
rect 15068 29344 15084 29408
rect 15148 29344 15154 29408
rect 14838 29343 15154 29344
rect 21784 29408 22100 29409
rect 21784 29344 21790 29408
rect 21854 29344 21870 29408
rect 21934 29344 21950 29408
rect 22014 29344 22030 29408
rect 22094 29344 22100 29408
rect 21784 29343 22100 29344
rect 28730 29408 29046 29409
rect 28730 29344 28736 29408
rect 28800 29344 28816 29408
rect 28880 29344 28896 29408
rect 28960 29344 28976 29408
rect 29040 29344 29046 29408
rect 28730 29343 29046 29344
rect 29200 29338 29800 29428
rect 29200 29278 29930 29338
rect 29200 29202 29800 29278
rect 29870 29202 29930 29278
rect 29200 29188 29930 29202
rect 29318 29142 29930 29188
rect 24761 29066 24827 29069
rect 29318 29066 29378 29142
rect 24761 29064 29378 29066
rect 24761 29008 24766 29064
rect 24822 29008 29378 29064
rect 24761 29006 29378 29008
rect 24761 29003 24827 29006
rect 4419 28864 4735 28865
rect 4419 28800 4425 28864
rect 4489 28800 4505 28864
rect 4569 28800 4585 28864
rect 4649 28800 4665 28864
rect 4729 28800 4735 28864
rect 4419 28799 4735 28800
rect 11365 28864 11681 28865
rect 11365 28800 11371 28864
rect 11435 28800 11451 28864
rect 11515 28800 11531 28864
rect 11595 28800 11611 28864
rect 11675 28800 11681 28864
rect 11365 28799 11681 28800
rect 18311 28864 18627 28865
rect 18311 28800 18317 28864
rect 18381 28800 18397 28864
rect 18461 28800 18477 28864
rect 18541 28800 18557 28864
rect 18621 28800 18627 28864
rect 18311 28799 18627 28800
rect 25257 28864 25573 28865
rect 25257 28800 25263 28864
rect 25327 28800 25343 28864
rect 25407 28800 25423 28864
rect 25487 28800 25503 28864
rect 25567 28800 25573 28864
rect 25257 28799 25573 28800
rect 200 28508 800 28748
rect 27521 28658 27587 28661
rect 29200 28658 29800 28748
rect 27521 28656 29800 28658
rect 27521 28600 27526 28656
rect 27582 28600 29800 28656
rect 27521 28598 29800 28600
rect 27521 28595 27587 28598
rect 29200 28508 29800 28598
rect 7892 28320 8208 28321
rect 7892 28256 7898 28320
rect 7962 28256 7978 28320
rect 8042 28256 8058 28320
rect 8122 28256 8138 28320
rect 8202 28256 8208 28320
rect 7892 28255 8208 28256
rect 14838 28320 15154 28321
rect 14838 28256 14844 28320
rect 14908 28256 14924 28320
rect 14988 28256 15004 28320
rect 15068 28256 15084 28320
rect 15148 28256 15154 28320
rect 14838 28255 15154 28256
rect 21784 28320 22100 28321
rect 21784 28256 21790 28320
rect 21854 28256 21870 28320
rect 21934 28256 21950 28320
rect 22014 28256 22030 28320
rect 22094 28256 22100 28320
rect 21784 28255 22100 28256
rect 28730 28320 29046 28321
rect 28730 28256 28736 28320
rect 28800 28256 28816 28320
rect 28880 28256 28896 28320
rect 28960 28256 28976 28320
rect 29040 28256 29046 28320
rect 28730 28255 29046 28256
rect 200 27978 800 28068
rect 1577 27978 1643 27981
rect 18873 27980 18939 27981
rect 200 27976 1643 27978
rect 200 27920 1582 27976
rect 1638 27920 1643 27976
rect 200 27918 1643 27920
rect 200 27828 800 27918
rect 1577 27915 1643 27918
rect 18822 27916 18828 27980
rect 18892 27978 18939 27980
rect 18892 27976 18984 27978
rect 18934 27920 18984 27976
rect 18892 27918 18984 27920
rect 18892 27916 18939 27918
rect 18873 27915 18939 27916
rect 4419 27776 4735 27777
rect 4419 27712 4425 27776
rect 4489 27712 4505 27776
rect 4569 27712 4585 27776
rect 4649 27712 4665 27776
rect 4729 27712 4735 27776
rect 4419 27711 4735 27712
rect 11365 27776 11681 27777
rect 11365 27712 11371 27776
rect 11435 27712 11451 27776
rect 11515 27712 11531 27776
rect 11595 27712 11611 27776
rect 11675 27712 11681 27776
rect 11365 27711 11681 27712
rect 18311 27776 18627 27777
rect 18311 27712 18317 27776
rect 18381 27712 18397 27776
rect 18461 27712 18477 27776
rect 18541 27712 18557 27776
rect 18621 27712 18627 27776
rect 18311 27711 18627 27712
rect 25257 27776 25573 27777
rect 25257 27712 25263 27776
rect 25327 27712 25343 27776
rect 25407 27712 25423 27776
rect 25487 27712 25503 27776
rect 25567 27712 25573 27776
rect 25257 27711 25573 27712
rect 27521 27570 27587 27573
rect 27521 27568 29378 27570
rect 27521 27512 27526 27568
rect 27582 27512 29378 27568
rect 27521 27510 29378 27512
rect 27521 27507 27587 27510
rect 29318 27434 29378 27510
rect 29318 27388 29930 27434
rect 29200 27374 29930 27388
rect 29200 27298 29800 27374
rect 29870 27298 29930 27374
rect 29200 27238 29930 27298
rect 7892 27232 8208 27233
rect 7892 27168 7898 27232
rect 7962 27168 7978 27232
rect 8042 27168 8058 27232
rect 8122 27168 8138 27232
rect 8202 27168 8208 27232
rect 7892 27167 8208 27168
rect 14838 27232 15154 27233
rect 14838 27168 14844 27232
rect 14908 27168 14924 27232
rect 14988 27168 15004 27232
rect 15068 27168 15084 27232
rect 15148 27168 15154 27232
rect 14838 27167 15154 27168
rect 21784 27232 22100 27233
rect 21784 27168 21790 27232
rect 21854 27168 21870 27232
rect 21934 27168 21950 27232
rect 22014 27168 22030 27232
rect 22094 27168 22100 27232
rect 21784 27167 22100 27168
rect 28730 27232 29046 27233
rect 28730 27168 28736 27232
rect 28800 27168 28816 27232
rect 28880 27168 28896 27232
rect 28960 27168 28976 27232
rect 29040 27168 29046 27232
rect 28730 27167 29046 27168
rect 29200 27148 29800 27238
rect 200 26468 800 26708
rect 4419 26688 4735 26689
rect 4419 26624 4425 26688
rect 4489 26624 4505 26688
rect 4569 26624 4585 26688
rect 4649 26624 4665 26688
rect 4729 26624 4735 26688
rect 4419 26623 4735 26624
rect 11365 26688 11681 26689
rect 11365 26624 11371 26688
rect 11435 26624 11451 26688
rect 11515 26624 11531 26688
rect 11595 26624 11611 26688
rect 11675 26624 11681 26688
rect 11365 26623 11681 26624
rect 18311 26688 18627 26689
rect 18311 26624 18317 26688
rect 18381 26624 18397 26688
rect 18461 26624 18477 26688
rect 18541 26624 18557 26688
rect 18621 26624 18627 26688
rect 18311 26623 18627 26624
rect 25257 26688 25573 26689
rect 25257 26624 25263 26688
rect 25327 26624 25343 26688
rect 25407 26624 25423 26688
rect 25487 26624 25503 26688
rect 25567 26624 25573 26688
rect 25257 26623 25573 26624
rect 28349 26618 28415 26621
rect 29200 26618 29800 26708
rect 28349 26616 29800 26618
rect 28349 26560 28354 26616
rect 28410 26560 29800 26616
rect 28349 26558 29800 26560
rect 28349 26555 28415 26558
rect 29200 26468 29800 26558
rect 7892 26144 8208 26145
rect 7892 26080 7898 26144
rect 7962 26080 7978 26144
rect 8042 26080 8058 26144
rect 8122 26080 8138 26144
rect 8202 26080 8208 26144
rect 7892 26079 8208 26080
rect 14838 26144 15154 26145
rect 14838 26080 14844 26144
rect 14908 26080 14924 26144
rect 14988 26080 15004 26144
rect 15068 26080 15084 26144
rect 15148 26080 15154 26144
rect 14838 26079 15154 26080
rect 21784 26144 22100 26145
rect 21784 26080 21790 26144
rect 21854 26080 21870 26144
rect 21934 26080 21950 26144
rect 22014 26080 22030 26144
rect 22094 26080 22100 26144
rect 21784 26079 22100 26080
rect 28730 26144 29046 26145
rect 28730 26080 28736 26144
rect 28800 26080 28816 26144
rect 28880 26080 28896 26144
rect 28960 26080 28976 26144
rect 29040 26080 29046 26144
rect 28730 26079 29046 26080
rect 200 25938 800 26028
rect 2773 25938 2839 25941
rect 200 25936 2839 25938
rect 200 25880 2778 25936
rect 2834 25880 2839 25936
rect 200 25878 2839 25880
rect 200 25788 800 25878
rect 2773 25875 2839 25878
rect 29200 25788 29800 26028
rect 4419 25600 4735 25601
rect 4419 25536 4425 25600
rect 4489 25536 4505 25600
rect 4569 25536 4585 25600
rect 4649 25536 4665 25600
rect 4729 25536 4735 25600
rect 4419 25535 4735 25536
rect 11365 25600 11681 25601
rect 11365 25536 11371 25600
rect 11435 25536 11451 25600
rect 11515 25536 11531 25600
rect 11595 25536 11611 25600
rect 11675 25536 11681 25600
rect 11365 25535 11681 25536
rect 18311 25600 18627 25601
rect 18311 25536 18317 25600
rect 18381 25536 18397 25600
rect 18461 25536 18477 25600
rect 18541 25536 18557 25600
rect 18621 25536 18627 25600
rect 18311 25535 18627 25536
rect 25257 25600 25573 25601
rect 25257 25536 25263 25600
rect 25327 25536 25343 25600
rect 25407 25536 25423 25600
rect 25487 25536 25503 25600
rect 25567 25536 25573 25600
rect 25257 25535 25573 25536
rect 200 25258 800 25348
rect 1577 25258 1643 25261
rect 200 25256 1643 25258
rect 200 25200 1582 25256
rect 1638 25200 1643 25256
rect 200 25198 1643 25200
rect 200 25108 800 25198
rect 1577 25195 1643 25198
rect 27521 25258 27587 25261
rect 29200 25258 29800 25348
rect 27521 25256 29800 25258
rect 27521 25200 27526 25256
rect 27582 25200 29800 25256
rect 27521 25198 29800 25200
rect 27521 25195 27587 25198
rect 29200 25108 29800 25198
rect 7892 25056 8208 25057
rect 7892 24992 7898 25056
rect 7962 24992 7978 25056
rect 8042 24992 8058 25056
rect 8122 24992 8138 25056
rect 8202 24992 8208 25056
rect 7892 24991 8208 24992
rect 14838 25056 15154 25057
rect 14838 24992 14844 25056
rect 14908 24992 14924 25056
rect 14988 24992 15004 25056
rect 15068 24992 15084 25056
rect 15148 24992 15154 25056
rect 14838 24991 15154 24992
rect 21784 25056 22100 25057
rect 21784 24992 21790 25056
rect 21854 24992 21870 25056
rect 21934 24992 21950 25056
rect 22014 24992 22030 25056
rect 22094 24992 22100 25056
rect 21784 24991 22100 24992
rect 28730 25056 29046 25057
rect 28730 24992 28736 25056
rect 28800 24992 28816 25056
rect 28880 24992 28896 25056
rect 28960 24992 28976 25056
rect 29040 24992 29046 25056
rect 28730 24991 29046 24992
rect 200 24428 800 24668
rect 28349 24578 28415 24581
rect 29200 24578 29800 24668
rect 28349 24576 29800 24578
rect 28349 24520 28354 24576
rect 28410 24520 29800 24576
rect 28349 24518 29800 24520
rect 28349 24515 28415 24518
rect 4419 24512 4735 24513
rect 4419 24448 4425 24512
rect 4489 24448 4505 24512
rect 4569 24448 4585 24512
rect 4649 24448 4665 24512
rect 4729 24448 4735 24512
rect 4419 24447 4735 24448
rect 11365 24512 11681 24513
rect 11365 24448 11371 24512
rect 11435 24448 11451 24512
rect 11515 24448 11531 24512
rect 11595 24448 11611 24512
rect 11675 24448 11681 24512
rect 11365 24447 11681 24448
rect 18311 24512 18627 24513
rect 18311 24448 18317 24512
rect 18381 24448 18397 24512
rect 18461 24448 18477 24512
rect 18541 24448 18557 24512
rect 18621 24448 18627 24512
rect 18311 24447 18627 24448
rect 25257 24512 25573 24513
rect 25257 24448 25263 24512
rect 25327 24448 25343 24512
rect 25407 24448 25423 24512
rect 25487 24448 25503 24512
rect 25567 24448 25573 24512
rect 25257 24447 25573 24448
rect 29200 24428 29800 24518
rect 200 23748 800 23988
rect 7892 23968 8208 23969
rect 7892 23904 7898 23968
rect 7962 23904 7978 23968
rect 8042 23904 8058 23968
rect 8122 23904 8138 23968
rect 8202 23904 8208 23968
rect 7892 23903 8208 23904
rect 14838 23968 15154 23969
rect 14838 23904 14844 23968
rect 14908 23904 14924 23968
rect 14988 23904 15004 23968
rect 15068 23904 15084 23968
rect 15148 23904 15154 23968
rect 14838 23903 15154 23904
rect 21784 23968 22100 23969
rect 21784 23904 21790 23968
rect 21854 23904 21870 23968
rect 21934 23904 21950 23968
rect 22014 23904 22030 23968
rect 22094 23904 22100 23968
rect 21784 23903 22100 23904
rect 28730 23968 29046 23969
rect 28730 23904 28736 23968
rect 28800 23904 28816 23968
rect 28880 23904 28896 23968
rect 28960 23904 28976 23968
rect 29040 23904 29046 23968
rect 28730 23903 29046 23904
rect 29200 23898 29800 23988
rect 29913 23898 29979 23901
rect 29200 23896 29979 23898
rect 29200 23840 29918 23896
rect 29974 23840 29979 23896
rect 29200 23838 29979 23840
rect 29200 23748 29800 23838
rect 29913 23835 29979 23838
rect 4419 23424 4735 23425
rect 4419 23360 4425 23424
rect 4489 23360 4505 23424
rect 4569 23360 4585 23424
rect 4649 23360 4665 23424
rect 4729 23360 4735 23424
rect 4419 23359 4735 23360
rect 11365 23424 11681 23425
rect 11365 23360 11371 23424
rect 11435 23360 11451 23424
rect 11515 23360 11531 23424
rect 11595 23360 11611 23424
rect 11675 23360 11681 23424
rect 11365 23359 11681 23360
rect 18311 23424 18627 23425
rect 18311 23360 18317 23424
rect 18381 23360 18397 23424
rect 18461 23360 18477 23424
rect 18541 23360 18557 23424
rect 18621 23360 18627 23424
rect 18311 23359 18627 23360
rect 25257 23424 25573 23425
rect 25257 23360 25263 23424
rect 25327 23360 25343 23424
rect 25407 23360 25423 23424
rect 25487 23360 25503 23424
rect 25567 23360 25573 23424
rect 25257 23359 25573 23360
rect 200 23068 800 23308
rect 29200 23068 29800 23308
rect 7892 22880 8208 22881
rect 7892 22816 7898 22880
rect 7962 22816 7978 22880
rect 8042 22816 8058 22880
rect 8122 22816 8138 22880
rect 8202 22816 8208 22880
rect 7892 22815 8208 22816
rect 14838 22880 15154 22881
rect 14838 22816 14844 22880
rect 14908 22816 14924 22880
rect 14988 22816 15004 22880
rect 15068 22816 15084 22880
rect 15148 22816 15154 22880
rect 14838 22815 15154 22816
rect 21784 22880 22100 22881
rect 21784 22816 21790 22880
rect 21854 22816 21870 22880
rect 21934 22816 21950 22880
rect 22014 22816 22030 22880
rect 22094 22816 22100 22880
rect 21784 22815 22100 22816
rect 28730 22880 29046 22881
rect 28730 22816 28736 22880
rect 28800 22816 28816 22880
rect 28880 22816 28896 22880
rect 28960 22816 28976 22880
rect 29040 22816 29046 22880
rect 28730 22815 29046 22816
rect 200 22388 800 22628
rect 4419 22336 4735 22337
rect 4419 22272 4425 22336
rect 4489 22272 4505 22336
rect 4569 22272 4585 22336
rect 4649 22272 4665 22336
rect 4729 22272 4735 22336
rect 4419 22271 4735 22272
rect 11365 22336 11681 22337
rect 11365 22272 11371 22336
rect 11435 22272 11451 22336
rect 11515 22272 11531 22336
rect 11595 22272 11611 22336
rect 11675 22272 11681 22336
rect 11365 22271 11681 22272
rect 18311 22336 18627 22337
rect 18311 22272 18317 22336
rect 18381 22272 18397 22336
rect 18461 22272 18477 22336
rect 18541 22272 18557 22336
rect 18621 22272 18627 22336
rect 18311 22271 18627 22272
rect 25257 22336 25573 22337
rect 25257 22272 25263 22336
rect 25327 22272 25343 22336
rect 25407 22272 25423 22336
rect 25487 22272 25503 22336
rect 25567 22272 25573 22336
rect 25257 22271 25573 22272
rect 29200 21858 29800 21948
rect 29200 21798 29930 21858
rect 7892 21792 8208 21793
rect 7892 21728 7898 21792
rect 7962 21728 7978 21792
rect 8042 21728 8058 21792
rect 8122 21728 8138 21792
rect 8202 21728 8208 21792
rect 7892 21727 8208 21728
rect 14838 21792 15154 21793
rect 14838 21728 14844 21792
rect 14908 21728 14924 21792
rect 14988 21728 15004 21792
rect 15068 21728 15084 21792
rect 15148 21728 15154 21792
rect 14838 21727 15154 21728
rect 21784 21792 22100 21793
rect 21784 21728 21790 21792
rect 21854 21728 21870 21792
rect 21934 21728 21950 21792
rect 22014 21728 22030 21792
rect 22094 21728 22100 21792
rect 21784 21727 22100 21728
rect 28730 21792 29046 21793
rect 28730 21728 28736 21792
rect 28800 21728 28816 21792
rect 28880 21728 28896 21792
rect 28960 21728 28976 21792
rect 29040 21728 29046 21792
rect 28730 21727 29046 21728
rect 29200 21722 29800 21798
rect 29870 21722 29930 21798
rect 29200 21708 29930 21722
rect 29318 21662 29930 21708
rect 26141 21450 26207 21453
rect 29318 21450 29378 21662
rect 26141 21448 29378 21450
rect 26141 21392 26146 21448
rect 26202 21392 29378 21448
rect 26141 21390 29378 21392
rect 26141 21387 26207 21390
rect 200 21028 800 21268
rect 4419 21248 4735 21249
rect 4419 21184 4425 21248
rect 4489 21184 4505 21248
rect 4569 21184 4585 21248
rect 4649 21184 4665 21248
rect 4729 21184 4735 21248
rect 4419 21183 4735 21184
rect 11365 21248 11681 21249
rect 11365 21184 11371 21248
rect 11435 21184 11451 21248
rect 11515 21184 11531 21248
rect 11595 21184 11611 21248
rect 11675 21184 11681 21248
rect 11365 21183 11681 21184
rect 18311 21248 18627 21249
rect 18311 21184 18317 21248
rect 18381 21184 18397 21248
rect 18461 21184 18477 21248
rect 18541 21184 18557 21248
rect 18621 21184 18627 21248
rect 18311 21183 18627 21184
rect 25257 21248 25573 21249
rect 25257 21184 25263 21248
rect 25327 21184 25343 21248
rect 25407 21184 25423 21248
rect 25487 21184 25503 21248
rect 25567 21184 25573 21248
rect 25257 21183 25573 21184
rect 27521 21178 27587 21181
rect 29200 21178 29800 21268
rect 27521 21176 29800 21178
rect 27521 21120 27526 21176
rect 27582 21120 29800 21176
rect 27521 21118 29800 21120
rect 27521 21115 27587 21118
rect 29200 21028 29800 21118
rect 7892 20704 8208 20705
rect 7892 20640 7898 20704
rect 7962 20640 7978 20704
rect 8042 20640 8058 20704
rect 8122 20640 8138 20704
rect 8202 20640 8208 20704
rect 7892 20639 8208 20640
rect 14838 20704 15154 20705
rect 14838 20640 14844 20704
rect 14908 20640 14924 20704
rect 14988 20640 15004 20704
rect 15068 20640 15084 20704
rect 15148 20640 15154 20704
rect 14838 20639 15154 20640
rect 21784 20704 22100 20705
rect 21784 20640 21790 20704
rect 21854 20640 21870 20704
rect 21934 20640 21950 20704
rect 22014 20640 22030 20704
rect 22094 20640 22100 20704
rect 21784 20639 22100 20640
rect 28730 20704 29046 20705
rect 28730 20640 28736 20704
rect 28800 20640 28816 20704
rect 28880 20640 28896 20704
rect 28960 20640 28976 20704
rect 29040 20640 29046 20704
rect 28730 20639 29046 20640
rect 200 20348 800 20588
rect 27521 20498 27587 20501
rect 29200 20498 29800 20588
rect 27521 20496 29800 20498
rect 27521 20440 27526 20496
rect 27582 20440 29800 20496
rect 27521 20438 29800 20440
rect 27521 20435 27587 20438
rect 29200 20348 29800 20438
rect 4419 20160 4735 20161
rect 4419 20096 4425 20160
rect 4489 20096 4505 20160
rect 4569 20096 4585 20160
rect 4649 20096 4665 20160
rect 4729 20096 4735 20160
rect 4419 20095 4735 20096
rect 11365 20160 11681 20161
rect 11365 20096 11371 20160
rect 11435 20096 11451 20160
rect 11515 20096 11531 20160
rect 11595 20096 11611 20160
rect 11675 20096 11681 20160
rect 11365 20095 11681 20096
rect 18311 20160 18627 20161
rect 18311 20096 18317 20160
rect 18381 20096 18397 20160
rect 18461 20096 18477 20160
rect 18541 20096 18557 20160
rect 18621 20096 18627 20160
rect 18311 20095 18627 20096
rect 25257 20160 25573 20161
rect 25257 20096 25263 20160
rect 25327 20096 25343 20160
rect 25407 20096 25423 20160
rect 25487 20096 25503 20160
rect 25567 20096 25573 20160
rect 25257 20095 25573 20096
rect 200 19818 800 19908
rect 2773 19818 2839 19821
rect 200 19816 2839 19818
rect 200 19760 2778 19816
rect 2834 19760 2839 19816
rect 200 19758 2839 19760
rect 200 19668 800 19758
rect 2773 19755 2839 19758
rect 28625 19818 28691 19821
rect 29200 19818 29800 19908
rect 28625 19816 29800 19818
rect 28625 19760 28630 19816
rect 28686 19760 29800 19816
rect 28625 19758 29800 19760
rect 28625 19755 28691 19758
rect 29200 19668 29800 19758
rect 7892 19616 8208 19617
rect 7892 19552 7898 19616
rect 7962 19552 7978 19616
rect 8042 19552 8058 19616
rect 8122 19552 8138 19616
rect 8202 19552 8208 19616
rect 7892 19551 8208 19552
rect 14838 19616 15154 19617
rect 14838 19552 14844 19616
rect 14908 19552 14924 19616
rect 14988 19552 15004 19616
rect 15068 19552 15084 19616
rect 15148 19552 15154 19616
rect 14838 19551 15154 19552
rect 21784 19616 22100 19617
rect 21784 19552 21790 19616
rect 21854 19552 21870 19616
rect 21934 19552 21950 19616
rect 22014 19552 22030 19616
rect 22094 19552 22100 19616
rect 21784 19551 22100 19552
rect 28730 19616 29046 19617
rect 28730 19552 28736 19616
rect 28800 19552 28816 19616
rect 28880 19552 28896 19616
rect 28960 19552 28976 19616
rect 29040 19552 29046 19616
rect 28730 19551 29046 19552
rect 200 19138 800 19228
rect 2129 19138 2195 19141
rect 200 19136 2195 19138
rect 200 19080 2134 19136
rect 2190 19080 2195 19136
rect 200 19078 2195 19080
rect 200 18988 800 19078
rect 2129 19075 2195 19078
rect 4419 19072 4735 19073
rect 4419 19008 4425 19072
rect 4489 19008 4505 19072
rect 4569 19008 4585 19072
rect 4649 19008 4665 19072
rect 4729 19008 4735 19072
rect 4419 19007 4735 19008
rect 11365 19072 11681 19073
rect 11365 19008 11371 19072
rect 11435 19008 11451 19072
rect 11515 19008 11531 19072
rect 11595 19008 11611 19072
rect 11675 19008 11681 19072
rect 11365 19007 11681 19008
rect 18311 19072 18627 19073
rect 18311 19008 18317 19072
rect 18381 19008 18397 19072
rect 18461 19008 18477 19072
rect 18541 19008 18557 19072
rect 18621 19008 18627 19072
rect 18311 19007 18627 19008
rect 25257 19072 25573 19073
rect 25257 19008 25263 19072
rect 25327 19008 25343 19072
rect 25407 19008 25423 19072
rect 25487 19008 25503 19072
rect 25567 19008 25573 19072
rect 25257 19007 25573 19008
rect 29200 18988 29800 19228
rect 200 18458 800 18548
rect 7892 18528 8208 18529
rect 7892 18464 7898 18528
rect 7962 18464 7978 18528
rect 8042 18464 8058 18528
rect 8122 18464 8138 18528
rect 8202 18464 8208 18528
rect 7892 18463 8208 18464
rect 14838 18528 15154 18529
rect 14838 18464 14844 18528
rect 14908 18464 14924 18528
rect 14988 18464 15004 18528
rect 15068 18464 15084 18528
rect 15148 18464 15154 18528
rect 14838 18463 15154 18464
rect 21784 18528 22100 18529
rect 21784 18464 21790 18528
rect 21854 18464 21870 18528
rect 21934 18464 21950 18528
rect 22014 18464 22030 18528
rect 22094 18464 22100 18528
rect 21784 18463 22100 18464
rect 28730 18528 29046 18529
rect 28730 18464 28736 18528
rect 28800 18464 28816 18528
rect 28880 18464 28896 18528
rect 28960 18464 28976 18528
rect 29040 18464 29046 18528
rect 28730 18463 29046 18464
rect 1577 18458 1643 18461
rect 200 18456 1643 18458
rect 200 18400 1582 18456
rect 1638 18400 1643 18456
rect 200 18398 1643 18400
rect 200 18308 800 18398
rect 1577 18395 1643 18398
rect 29200 18308 29800 18548
rect 4419 17984 4735 17985
rect 4419 17920 4425 17984
rect 4489 17920 4505 17984
rect 4569 17920 4585 17984
rect 4649 17920 4665 17984
rect 4729 17920 4735 17984
rect 4419 17919 4735 17920
rect 11365 17984 11681 17985
rect 11365 17920 11371 17984
rect 11435 17920 11451 17984
rect 11515 17920 11531 17984
rect 11595 17920 11611 17984
rect 11675 17920 11681 17984
rect 11365 17919 11681 17920
rect 18311 17984 18627 17985
rect 18311 17920 18317 17984
rect 18381 17920 18397 17984
rect 18461 17920 18477 17984
rect 18541 17920 18557 17984
rect 18621 17920 18627 17984
rect 18311 17919 18627 17920
rect 25257 17984 25573 17985
rect 25257 17920 25263 17984
rect 25327 17920 25343 17984
rect 25407 17920 25423 17984
rect 25487 17920 25503 17984
rect 25567 17920 25573 17984
rect 25257 17919 25573 17920
rect 200 17778 800 17868
rect 2773 17778 2839 17781
rect 200 17776 2839 17778
rect 200 17720 2778 17776
rect 2834 17720 2839 17776
rect 200 17718 2839 17720
rect 200 17628 800 17718
rect 2773 17715 2839 17718
rect 29200 17628 29800 17868
rect 7892 17440 8208 17441
rect 7892 17376 7898 17440
rect 7962 17376 7978 17440
rect 8042 17376 8058 17440
rect 8122 17376 8138 17440
rect 8202 17376 8208 17440
rect 7892 17375 8208 17376
rect 14838 17440 15154 17441
rect 14838 17376 14844 17440
rect 14908 17376 14924 17440
rect 14988 17376 15004 17440
rect 15068 17376 15084 17440
rect 15148 17376 15154 17440
rect 14838 17375 15154 17376
rect 21784 17440 22100 17441
rect 21784 17376 21790 17440
rect 21854 17376 21870 17440
rect 21934 17376 21950 17440
rect 22014 17376 22030 17440
rect 22094 17376 22100 17440
rect 21784 17375 22100 17376
rect 28730 17440 29046 17441
rect 28730 17376 28736 17440
rect 28800 17376 28816 17440
rect 28880 17376 28896 17440
rect 28960 17376 28976 17440
rect 29040 17376 29046 17440
rect 28730 17375 29046 17376
rect 200 16948 800 17188
rect 4419 16896 4735 16897
rect 4419 16832 4425 16896
rect 4489 16832 4505 16896
rect 4569 16832 4585 16896
rect 4649 16832 4665 16896
rect 4729 16832 4735 16896
rect 4419 16831 4735 16832
rect 11365 16896 11681 16897
rect 11365 16832 11371 16896
rect 11435 16832 11451 16896
rect 11515 16832 11531 16896
rect 11595 16832 11611 16896
rect 11675 16832 11681 16896
rect 11365 16831 11681 16832
rect 18311 16896 18627 16897
rect 18311 16832 18317 16896
rect 18381 16832 18397 16896
rect 18461 16832 18477 16896
rect 18541 16832 18557 16896
rect 18621 16832 18627 16896
rect 18311 16831 18627 16832
rect 25257 16896 25573 16897
rect 25257 16832 25263 16896
rect 25327 16832 25343 16896
rect 25407 16832 25423 16896
rect 25487 16832 25503 16896
rect 25567 16832 25573 16896
rect 25257 16831 25573 16832
rect 29200 16418 29800 16508
rect 29913 16418 29979 16421
rect 29200 16416 29979 16418
rect 29200 16360 29918 16416
rect 29974 16360 29979 16416
rect 29200 16358 29979 16360
rect 7892 16352 8208 16353
rect 7892 16288 7898 16352
rect 7962 16288 7978 16352
rect 8042 16288 8058 16352
rect 8122 16288 8138 16352
rect 8202 16288 8208 16352
rect 7892 16287 8208 16288
rect 14838 16352 15154 16353
rect 14838 16288 14844 16352
rect 14908 16288 14924 16352
rect 14988 16288 15004 16352
rect 15068 16288 15084 16352
rect 15148 16288 15154 16352
rect 14838 16287 15154 16288
rect 21784 16352 22100 16353
rect 21784 16288 21790 16352
rect 21854 16288 21870 16352
rect 21934 16288 21950 16352
rect 22014 16288 22030 16352
rect 22094 16288 22100 16352
rect 21784 16287 22100 16288
rect 28730 16352 29046 16353
rect 28730 16288 28736 16352
rect 28800 16288 28816 16352
rect 28880 16288 28896 16352
rect 28960 16288 28976 16352
rect 29040 16288 29046 16352
rect 28730 16287 29046 16288
rect 29200 16268 29800 16358
rect 29913 16355 29979 16358
rect 200 15738 800 15828
rect 4419 15808 4735 15809
rect 4419 15744 4425 15808
rect 4489 15744 4505 15808
rect 4569 15744 4585 15808
rect 4649 15744 4665 15808
rect 4729 15744 4735 15808
rect 4419 15743 4735 15744
rect 11365 15808 11681 15809
rect 11365 15744 11371 15808
rect 11435 15744 11451 15808
rect 11515 15744 11531 15808
rect 11595 15744 11611 15808
rect 11675 15744 11681 15808
rect 11365 15743 11681 15744
rect 18311 15808 18627 15809
rect 18311 15744 18317 15808
rect 18381 15744 18397 15808
rect 18461 15744 18477 15808
rect 18541 15744 18557 15808
rect 18621 15744 18627 15808
rect 18311 15743 18627 15744
rect 25257 15808 25573 15809
rect 25257 15744 25263 15808
rect 25327 15744 25343 15808
rect 25407 15744 25423 15808
rect 25487 15744 25503 15808
rect 25567 15744 25573 15808
rect 25257 15743 25573 15744
rect 2773 15738 2839 15741
rect 200 15736 2839 15738
rect 200 15680 2778 15736
rect 2834 15680 2839 15736
rect 200 15678 2839 15680
rect 200 15588 800 15678
rect 2773 15675 2839 15678
rect 28625 15738 28691 15741
rect 29200 15738 29800 15828
rect 28625 15736 29800 15738
rect 28625 15680 28630 15736
rect 28686 15680 29800 15736
rect 28625 15678 29800 15680
rect 28625 15675 28691 15678
rect 29200 15588 29800 15678
rect 7892 15264 8208 15265
rect 7892 15200 7898 15264
rect 7962 15200 7978 15264
rect 8042 15200 8058 15264
rect 8122 15200 8138 15264
rect 8202 15200 8208 15264
rect 7892 15199 8208 15200
rect 14838 15264 15154 15265
rect 14838 15200 14844 15264
rect 14908 15200 14924 15264
rect 14988 15200 15004 15264
rect 15068 15200 15084 15264
rect 15148 15200 15154 15264
rect 14838 15199 15154 15200
rect 21784 15264 22100 15265
rect 21784 15200 21790 15264
rect 21854 15200 21870 15264
rect 21934 15200 21950 15264
rect 22014 15200 22030 15264
rect 22094 15200 22100 15264
rect 21784 15199 22100 15200
rect 28730 15264 29046 15265
rect 28730 15200 28736 15264
rect 28800 15200 28816 15264
rect 28880 15200 28896 15264
rect 28960 15200 28976 15264
rect 29040 15200 29046 15264
rect 28730 15199 29046 15200
rect 200 14908 800 15148
rect 25497 15058 25563 15061
rect 29200 15058 29800 15148
rect 25497 15056 29800 15058
rect 25497 15000 25502 15056
rect 25558 15000 29800 15056
rect 25497 14998 29800 15000
rect 25497 14995 25563 14998
rect 29200 14908 29800 14998
rect 4419 14720 4735 14721
rect 4419 14656 4425 14720
rect 4489 14656 4505 14720
rect 4569 14656 4585 14720
rect 4649 14656 4665 14720
rect 4729 14656 4735 14720
rect 4419 14655 4735 14656
rect 11365 14720 11681 14721
rect 11365 14656 11371 14720
rect 11435 14656 11451 14720
rect 11515 14656 11531 14720
rect 11595 14656 11611 14720
rect 11675 14656 11681 14720
rect 11365 14655 11681 14656
rect 18311 14720 18627 14721
rect 18311 14656 18317 14720
rect 18381 14656 18397 14720
rect 18461 14656 18477 14720
rect 18541 14656 18557 14720
rect 18621 14656 18627 14720
rect 18311 14655 18627 14656
rect 25257 14720 25573 14721
rect 25257 14656 25263 14720
rect 25327 14656 25343 14720
rect 25407 14656 25423 14720
rect 25487 14656 25503 14720
rect 25567 14656 25573 14720
rect 25257 14655 25573 14656
rect 200 14378 800 14468
rect 1577 14378 1643 14381
rect 200 14376 1643 14378
rect 200 14320 1582 14376
rect 1638 14320 1643 14376
rect 200 14318 1643 14320
rect 200 14228 800 14318
rect 1577 14315 1643 14318
rect 27521 14378 27587 14381
rect 29200 14378 29800 14468
rect 27521 14376 29800 14378
rect 27521 14320 27526 14376
rect 27582 14320 29800 14376
rect 27521 14318 29800 14320
rect 27521 14315 27587 14318
rect 29200 14228 29800 14318
rect 7892 14176 8208 14177
rect 7892 14112 7898 14176
rect 7962 14112 7978 14176
rect 8042 14112 8058 14176
rect 8122 14112 8138 14176
rect 8202 14112 8208 14176
rect 7892 14111 8208 14112
rect 14838 14176 15154 14177
rect 14838 14112 14844 14176
rect 14908 14112 14924 14176
rect 14988 14112 15004 14176
rect 15068 14112 15084 14176
rect 15148 14112 15154 14176
rect 14838 14111 15154 14112
rect 21784 14176 22100 14177
rect 21784 14112 21790 14176
rect 21854 14112 21870 14176
rect 21934 14112 21950 14176
rect 22014 14112 22030 14176
rect 22094 14112 22100 14176
rect 21784 14111 22100 14112
rect 28730 14176 29046 14177
rect 28730 14112 28736 14176
rect 28800 14112 28816 14176
rect 28880 14112 28896 14176
rect 28960 14112 28976 14176
rect 29040 14112 29046 14176
rect 28730 14111 29046 14112
rect 200 13698 800 13788
rect 1577 13698 1643 13701
rect 200 13696 1643 13698
rect 200 13640 1582 13696
rect 1638 13640 1643 13696
rect 200 13638 1643 13640
rect 200 13548 800 13638
rect 1577 13635 1643 13638
rect 4419 13632 4735 13633
rect 4419 13568 4425 13632
rect 4489 13568 4505 13632
rect 4569 13568 4585 13632
rect 4649 13568 4665 13632
rect 4729 13568 4735 13632
rect 4419 13567 4735 13568
rect 11365 13632 11681 13633
rect 11365 13568 11371 13632
rect 11435 13568 11451 13632
rect 11515 13568 11531 13632
rect 11595 13568 11611 13632
rect 11675 13568 11681 13632
rect 11365 13567 11681 13568
rect 18311 13632 18627 13633
rect 18311 13568 18317 13632
rect 18381 13568 18397 13632
rect 18461 13568 18477 13632
rect 18541 13568 18557 13632
rect 18621 13568 18627 13632
rect 18311 13567 18627 13568
rect 25257 13632 25573 13633
rect 25257 13568 25263 13632
rect 25327 13568 25343 13632
rect 25407 13568 25423 13632
rect 25487 13568 25503 13632
rect 25567 13568 25573 13632
rect 25257 13567 25573 13568
rect 29200 13548 29800 13788
rect 200 12868 800 13108
rect 7892 13088 8208 13089
rect 7892 13024 7898 13088
rect 7962 13024 7978 13088
rect 8042 13024 8058 13088
rect 8122 13024 8138 13088
rect 8202 13024 8208 13088
rect 7892 13023 8208 13024
rect 14838 13088 15154 13089
rect 14838 13024 14844 13088
rect 14908 13024 14924 13088
rect 14988 13024 15004 13088
rect 15068 13024 15084 13088
rect 15148 13024 15154 13088
rect 14838 13023 15154 13024
rect 21784 13088 22100 13089
rect 21784 13024 21790 13088
rect 21854 13024 21870 13088
rect 21934 13024 21950 13088
rect 22014 13024 22030 13088
rect 22094 13024 22100 13088
rect 21784 13023 22100 13024
rect 28730 13088 29046 13089
rect 28730 13024 28736 13088
rect 28800 13024 28816 13088
rect 28880 13024 28896 13088
rect 28960 13024 28976 13088
rect 29040 13024 29046 13088
rect 28730 13023 29046 13024
rect 29200 12868 29800 13108
rect 4419 12544 4735 12545
rect 4419 12480 4425 12544
rect 4489 12480 4505 12544
rect 4569 12480 4585 12544
rect 4649 12480 4665 12544
rect 4729 12480 4735 12544
rect 4419 12479 4735 12480
rect 11365 12544 11681 12545
rect 11365 12480 11371 12544
rect 11435 12480 11451 12544
rect 11515 12480 11531 12544
rect 11595 12480 11611 12544
rect 11675 12480 11681 12544
rect 11365 12479 11681 12480
rect 18311 12544 18627 12545
rect 18311 12480 18317 12544
rect 18381 12480 18397 12544
rect 18461 12480 18477 12544
rect 18541 12480 18557 12544
rect 18621 12480 18627 12544
rect 18311 12479 18627 12480
rect 25257 12544 25573 12545
rect 25257 12480 25263 12544
rect 25327 12480 25343 12544
rect 25407 12480 25423 12544
rect 25487 12480 25503 12544
rect 25567 12480 25573 12544
rect 25257 12479 25573 12480
rect 200 12338 800 12428
rect 3509 12338 3575 12341
rect 200 12336 3575 12338
rect 200 12280 3514 12336
rect 3570 12280 3575 12336
rect 200 12278 3575 12280
rect 200 12188 800 12278
rect 3509 12275 3575 12278
rect 28349 12338 28415 12341
rect 29200 12338 29800 12428
rect 28349 12336 29800 12338
rect 28349 12280 28354 12336
rect 28410 12280 29800 12336
rect 28349 12278 29800 12280
rect 28349 12275 28415 12278
rect 29200 12188 29800 12278
rect 7892 12000 8208 12001
rect 7892 11936 7898 12000
rect 7962 11936 7978 12000
rect 8042 11936 8058 12000
rect 8122 11936 8138 12000
rect 8202 11936 8208 12000
rect 7892 11935 8208 11936
rect 14838 12000 15154 12001
rect 14838 11936 14844 12000
rect 14908 11936 14924 12000
rect 14988 11936 15004 12000
rect 15068 11936 15084 12000
rect 15148 11936 15154 12000
rect 14838 11935 15154 11936
rect 21784 12000 22100 12001
rect 21784 11936 21790 12000
rect 21854 11936 21870 12000
rect 21934 11936 21950 12000
rect 22014 11936 22030 12000
rect 22094 11936 22100 12000
rect 21784 11935 22100 11936
rect 28730 12000 29046 12001
rect 28730 11936 28736 12000
rect 28800 11936 28816 12000
rect 28880 11936 28896 12000
rect 28960 11936 28976 12000
rect 29040 11936 29046 12000
rect 28730 11935 29046 11936
rect 18873 11932 18939 11933
rect 18822 11868 18828 11932
rect 18892 11930 18939 11932
rect 18892 11928 18984 11930
rect 18934 11872 18984 11928
rect 18892 11870 18984 11872
rect 18892 11868 18939 11870
rect 18873 11867 18939 11868
rect 200 11658 800 11748
rect 2773 11658 2839 11661
rect 200 11656 2839 11658
rect 200 11600 2778 11656
rect 2834 11600 2839 11656
rect 200 11598 2839 11600
rect 200 11508 800 11598
rect 2773 11595 2839 11598
rect 4419 11456 4735 11457
rect 4419 11392 4425 11456
rect 4489 11392 4505 11456
rect 4569 11392 4585 11456
rect 4649 11392 4665 11456
rect 4729 11392 4735 11456
rect 4419 11391 4735 11392
rect 11365 11456 11681 11457
rect 11365 11392 11371 11456
rect 11435 11392 11451 11456
rect 11515 11392 11531 11456
rect 11595 11392 11611 11456
rect 11675 11392 11681 11456
rect 11365 11391 11681 11392
rect 18311 11456 18627 11457
rect 18311 11392 18317 11456
rect 18381 11392 18397 11456
rect 18461 11392 18477 11456
rect 18541 11392 18557 11456
rect 18621 11392 18627 11456
rect 18311 11391 18627 11392
rect 25257 11456 25573 11457
rect 25257 11392 25263 11456
rect 25327 11392 25343 11456
rect 25407 11392 25423 11456
rect 25487 11392 25503 11456
rect 25567 11392 25573 11456
rect 25257 11391 25573 11392
rect 29200 10978 29800 11068
rect 29913 10978 29979 10981
rect 29200 10976 29979 10978
rect 29200 10920 29918 10976
rect 29974 10920 29979 10976
rect 29200 10918 29979 10920
rect 7892 10912 8208 10913
rect 7892 10848 7898 10912
rect 7962 10848 7978 10912
rect 8042 10848 8058 10912
rect 8122 10848 8138 10912
rect 8202 10848 8208 10912
rect 7892 10847 8208 10848
rect 14838 10912 15154 10913
rect 14838 10848 14844 10912
rect 14908 10848 14924 10912
rect 14988 10848 15004 10912
rect 15068 10848 15084 10912
rect 15148 10848 15154 10912
rect 14838 10847 15154 10848
rect 21784 10912 22100 10913
rect 21784 10848 21790 10912
rect 21854 10848 21870 10912
rect 21934 10848 21950 10912
rect 22014 10848 22030 10912
rect 22094 10848 22100 10912
rect 21784 10847 22100 10848
rect 28730 10912 29046 10913
rect 28730 10848 28736 10912
rect 28800 10848 28816 10912
rect 28880 10848 28896 10912
rect 28960 10848 28976 10912
rect 29040 10848 29046 10912
rect 28730 10847 29046 10848
rect 29200 10828 29800 10918
rect 29913 10915 29979 10918
rect 200 10148 800 10388
rect 4419 10368 4735 10369
rect 4419 10304 4425 10368
rect 4489 10304 4505 10368
rect 4569 10304 4585 10368
rect 4649 10304 4665 10368
rect 4729 10304 4735 10368
rect 4419 10303 4735 10304
rect 11365 10368 11681 10369
rect 11365 10304 11371 10368
rect 11435 10304 11451 10368
rect 11515 10304 11531 10368
rect 11595 10304 11611 10368
rect 11675 10304 11681 10368
rect 11365 10303 11681 10304
rect 18311 10368 18627 10369
rect 18311 10304 18317 10368
rect 18381 10304 18397 10368
rect 18461 10304 18477 10368
rect 18541 10304 18557 10368
rect 18621 10304 18627 10368
rect 18311 10303 18627 10304
rect 25257 10368 25573 10369
rect 25257 10304 25263 10368
rect 25327 10304 25343 10368
rect 25407 10304 25423 10368
rect 25487 10304 25503 10368
rect 25567 10304 25573 10368
rect 25257 10303 25573 10304
rect 27521 10298 27587 10301
rect 29200 10298 29800 10388
rect 27521 10296 29800 10298
rect 27521 10240 27526 10296
rect 27582 10240 29800 10296
rect 27521 10238 29800 10240
rect 27521 10235 27587 10238
rect 29200 10148 29800 10238
rect 7892 9824 8208 9825
rect 7892 9760 7898 9824
rect 7962 9760 7978 9824
rect 8042 9760 8058 9824
rect 8122 9760 8138 9824
rect 8202 9760 8208 9824
rect 7892 9759 8208 9760
rect 14838 9824 15154 9825
rect 14838 9760 14844 9824
rect 14908 9760 14924 9824
rect 14988 9760 15004 9824
rect 15068 9760 15084 9824
rect 15148 9760 15154 9824
rect 14838 9759 15154 9760
rect 21784 9824 22100 9825
rect 21784 9760 21790 9824
rect 21854 9760 21870 9824
rect 21934 9760 21950 9824
rect 22014 9760 22030 9824
rect 22094 9760 22100 9824
rect 21784 9759 22100 9760
rect 28730 9824 29046 9825
rect 28730 9760 28736 9824
rect 28800 9760 28816 9824
rect 28880 9760 28896 9824
rect 28960 9760 28976 9824
rect 29040 9760 29046 9824
rect 28730 9759 29046 9760
rect 200 9468 800 9708
rect 29200 9468 29800 9708
rect 4419 9280 4735 9281
rect 4419 9216 4425 9280
rect 4489 9216 4505 9280
rect 4569 9216 4585 9280
rect 4649 9216 4665 9280
rect 4729 9216 4735 9280
rect 4419 9215 4735 9216
rect 11365 9280 11681 9281
rect 11365 9216 11371 9280
rect 11435 9216 11451 9280
rect 11515 9216 11531 9280
rect 11595 9216 11611 9280
rect 11675 9216 11681 9280
rect 11365 9215 11681 9216
rect 18311 9280 18627 9281
rect 18311 9216 18317 9280
rect 18381 9216 18397 9280
rect 18461 9216 18477 9280
rect 18541 9216 18557 9280
rect 18621 9216 18627 9280
rect 18311 9215 18627 9216
rect 25257 9280 25573 9281
rect 25257 9216 25263 9280
rect 25327 9216 25343 9280
rect 25407 9216 25423 9280
rect 25487 9216 25503 9280
rect 25567 9216 25573 9280
rect 25257 9215 25573 9216
rect 200 8938 800 9028
rect 2773 8938 2839 8941
rect 200 8936 2839 8938
rect 200 8880 2778 8936
rect 2834 8880 2839 8936
rect 200 8878 2839 8880
rect 200 8788 800 8878
rect 2773 8875 2839 8878
rect 28349 8938 28415 8941
rect 29200 8938 29800 9028
rect 28349 8936 29800 8938
rect 28349 8880 28354 8936
rect 28410 8880 29800 8936
rect 28349 8878 29800 8880
rect 28349 8875 28415 8878
rect 29200 8788 29800 8878
rect 7892 8736 8208 8737
rect 7892 8672 7898 8736
rect 7962 8672 7978 8736
rect 8042 8672 8058 8736
rect 8122 8672 8138 8736
rect 8202 8672 8208 8736
rect 7892 8671 8208 8672
rect 14838 8736 15154 8737
rect 14838 8672 14844 8736
rect 14908 8672 14924 8736
rect 14988 8672 15004 8736
rect 15068 8672 15084 8736
rect 15148 8672 15154 8736
rect 14838 8671 15154 8672
rect 21784 8736 22100 8737
rect 21784 8672 21790 8736
rect 21854 8672 21870 8736
rect 21934 8672 21950 8736
rect 22014 8672 22030 8736
rect 22094 8672 22100 8736
rect 21784 8671 22100 8672
rect 28730 8736 29046 8737
rect 28730 8672 28736 8736
rect 28800 8672 28816 8736
rect 28880 8672 28896 8736
rect 28960 8672 28976 8736
rect 29040 8672 29046 8736
rect 28730 8671 29046 8672
rect 200 8258 800 8348
rect 2957 8258 3023 8261
rect 200 8256 3023 8258
rect 200 8200 2962 8256
rect 3018 8200 3023 8256
rect 200 8198 3023 8200
rect 200 8108 800 8198
rect 2957 8195 3023 8198
rect 26141 8258 26207 8261
rect 29200 8258 29800 8348
rect 26141 8256 29800 8258
rect 26141 8200 26146 8256
rect 26202 8200 29800 8256
rect 26141 8198 29800 8200
rect 26141 8195 26207 8198
rect 4419 8192 4735 8193
rect 4419 8128 4425 8192
rect 4489 8128 4505 8192
rect 4569 8128 4585 8192
rect 4649 8128 4665 8192
rect 4729 8128 4735 8192
rect 4419 8127 4735 8128
rect 11365 8192 11681 8193
rect 11365 8128 11371 8192
rect 11435 8128 11451 8192
rect 11515 8128 11531 8192
rect 11595 8128 11611 8192
rect 11675 8128 11681 8192
rect 11365 8127 11681 8128
rect 18311 8192 18627 8193
rect 18311 8128 18317 8192
rect 18381 8128 18397 8192
rect 18461 8128 18477 8192
rect 18541 8128 18557 8192
rect 18621 8128 18627 8192
rect 18311 8127 18627 8128
rect 25257 8192 25573 8193
rect 25257 8128 25263 8192
rect 25327 8128 25343 8192
rect 25407 8128 25423 8192
rect 25487 8128 25503 8192
rect 25567 8128 25573 8192
rect 25257 8127 25573 8128
rect 29200 8108 29800 8198
rect 200 7578 800 7668
rect 7892 7648 8208 7649
rect 7892 7584 7898 7648
rect 7962 7584 7978 7648
rect 8042 7584 8058 7648
rect 8122 7584 8138 7648
rect 8202 7584 8208 7648
rect 7892 7583 8208 7584
rect 14838 7648 15154 7649
rect 14838 7584 14844 7648
rect 14908 7584 14924 7648
rect 14988 7584 15004 7648
rect 15068 7584 15084 7648
rect 15148 7584 15154 7648
rect 14838 7583 15154 7584
rect 21784 7648 22100 7649
rect 21784 7584 21790 7648
rect 21854 7584 21870 7648
rect 21934 7584 21950 7648
rect 22014 7584 22030 7648
rect 22094 7584 22100 7648
rect 21784 7583 22100 7584
rect 28730 7648 29046 7649
rect 28730 7584 28736 7648
rect 28800 7584 28816 7648
rect 28880 7584 28896 7648
rect 28960 7584 28976 7648
rect 29040 7584 29046 7648
rect 28730 7583 29046 7584
rect 3049 7578 3115 7581
rect 200 7576 3115 7578
rect 200 7520 3054 7576
rect 3110 7520 3115 7576
rect 200 7518 3115 7520
rect 200 7428 800 7518
rect 3049 7515 3115 7518
rect 29200 7578 29800 7668
rect 29913 7578 29979 7581
rect 29200 7576 29979 7578
rect 29200 7520 29918 7576
rect 29974 7520 29979 7576
rect 29200 7518 29979 7520
rect 29200 7428 29800 7518
rect 29913 7515 29979 7518
rect 4419 7104 4735 7105
rect 4419 7040 4425 7104
rect 4489 7040 4505 7104
rect 4569 7040 4585 7104
rect 4649 7040 4665 7104
rect 4729 7040 4735 7104
rect 4419 7039 4735 7040
rect 11365 7104 11681 7105
rect 11365 7040 11371 7104
rect 11435 7040 11451 7104
rect 11515 7040 11531 7104
rect 11595 7040 11611 7104
rect 11675 7040 11681 7104
rect 11365 7039 11681 7040
rect 18311 7104 18627 7105
rect 18311 7040 18317 7104
rect 18381 7040 18397 7104
rect 18461 7040 18477 7104
rect 18541 7040 18557 7104
rect 18621 7040 18627 7104
rect 18311 7039 18627 7040
rect 25257 7104 25573 7105
rect 25257 7040 25263 7104
rect 25327 7040 25343 7104
rect 25407 7040 25423 7104
rect 25487 7040 25503 7104
rect 25567 7040 25573 7104
rect 25257 7039 25573 7040
rect 200 6748 800 6988
rect 28349 6898 28415 6901
rect 29200 6898 29800 6988
rect 28349 6896 29800 6898
rect 28349 6840 28354 6896
rect 28410 6840 29800 6896
rect 28349 6838 29800 6840
rect 28349 6835 28415 6838
rect 29200 6748 29800 6838
rect 7892 6560 8208 6561
rect 7892 6496 7898 6560
rect 7962 6496 7978 6560
rect 8042 6496 8058 6560
rect 8122 6496 8138 6560
rect 8202 6496 8208 6560
rect 7892 6495 8208 6496
rect 14838 6560 15154 6561
rect 14838 6496 14844 6560
rect 14908 6496 14924 6560
rect 14988 6496 15004 6560
rect 15068 6496 15084 6560
rect 15148 6496 15154 6560
rect 14838 6495 15154 6496
rect 21784 6560 22100 6561
rect 21784 6496 21790 6560
rect 21854 6496 21870 6560
rect 21934 6496 21950 6560
rect 22014 6496 22030 6560
rect 22094 6496 22100 6560
rect 21784 6495 22100 6496
rect 28730 6560 29046 6561
rect 28730 6496 28736 6560
rect 28800 6496 28816 6560
rect 28880 6496 28896 6560
rect 28960 6496 28976 6560
rect 29040 6496 29046 6560
rect 28730 6495 29046 6496
rect 200 6218 800 6308
rect 4061 6218 4127 6221
rect 200 6216 4127 6218
rect 200 6160 4066 6216
rect 4122 6160 4127 6216
rect 200 6158 4127 6160
rect 200 6068 800 6158
rect 4061 6155 4127 6158
rect 4419 6016 4735 6017
rect 4419 5952 4425 6016
rect 4489 5952 4505 6016
rect 4569 5952 4585 6016
rect 4649 5952 4665 6016
rect 4729 5952 4735 6016
rect 4419 5951 4735 5952
rect 11365 6016 11681 6017
rect 11365 5952 11371 6016
rect 11435 5952 11451 6016
rect 11515 5952 11531 6016
rect 11595 5952 11611 6016
rect 11675 5952 11681 6016
rect 11365 5951 11681 5952
rect 18311 6016 18627 6017
rect 18311 5952 18317 6016
rect 18381 5952 18397 6016
rect 18461 5952 18477 6016
rect 18541 5952 18557 6016
rect 18621 5952 18627 6016
rect 18311 5951 18627 5952
rect 25257 6016 25573 6017
rect 25257 5952 25263 6016
rect 25327 5952 25343 6016
rect 25407 5952 25423 6016
rect 25487 5952 25503 6016
rect 25567 5952 25573 6016
rect 25257 5951 25573 5952
rect 29200 5538 29800 5628
rect 29200 5478 29930 5538
rect 7892 5472 8208 5473
rect 7892 5408 7898 5472
rect 7962 5408 7978 5472
rect 8042 5408 8058 5472
rect 8122 5408 8138 5472
rect 8202 5408 8208 5472
rect 7892 5407 8208 5408
rect 14838 5472 15154 5473
rect 14838 5408 14844 5472
rect 14908 5408 14924 5472
rect 14988 5408 15004 5472
rect 15068 5408 15084 5472
rect 15148 5408 15154 5472
rect 14838 5407 15154 5408
rect 21784 5472 22100 5473
rect 21784 5408 21790 5472
rect 21854 5408 21870 5472
rect 21934 5408 21950 5472
rect 22014 5408 22030 5472
rect 22094 5408 22100 5472
rect 21784 5407 22100 5408
rect 28730 5472 29046 5473
rect 28730 5408 28736 5472
rect 28800 5408 28816 5472
rect 28880 5408 28896 5472
rect 28960 5408 28976 5472
rect 29040 5408 29046 5472
rect 28730 5407 29046 5408
rect 29200 5402 29800 5478
rect 29870 5402 29930 5478
rect 29200 5388 29930 5402
rect 29318 5342 29930 5388
rect 27521 5266 27587 5269
rect 29318 5266 29378 5342
rect 27521 5264 29378 5266
rect 27521 5208 27526 5264
rect 27582 5208 29378 5264
rect 27521 5206 29378 5208
rect 27521 5203 27587 5206
rect 200 4858 800 4948
rect 4419 4928 4735 4929
rect 4419 4864 4425 4928
rect 4489 4864 4505 4928
rect 4569 4864 4585 4928
rect 4649 4864 4665 4928
rect 4729 4864 4735 4928
rect 4419 4863 4735 4864
rect 11365 4928 11681 4929
rect 11365 4864 11371 4928
rect 11435 4864 11451 4928
rect 11515 4864 11531 4928
rect 11595 4864 11611 4928
rect 11675 4864 11681 4928
rect 11365 4863 11681 4864
rect 18311 4928 18627 4929
rect 18311 4864 18317 4928
rect 18381 4864 18397 4928
rect 18461 4864 18477 4928
rect 18541 4864 18557 4928
rect 18621 4864 18627 4928
rect 18311 4863 18627 4864
rect 25257 4928 25573 4929
rect 25257 4864 25263 4928
rect 25327 4864 25343 4928
rect 25407 4864 25423 4928
rect 25487 4864 25503 4928
rect 25567 4864 25573 4928
rect 25257 4863 25573 4864
rect 3141 4858 3207 4861
rect 200 4856 3207 4858
rect 200 4800 3146 4856
rect 3202 4800 3207 4856
rect 200 4798 3207 4800
rect 200 4708 800 4798
rect 3141 4795 3207 4798
rect 29200 4708 29800 4948
rect 7892 4384 8208 4385
rect 7892 4320 7898 4384
rect 7962 4320 7978 4384
rect 8042 4320 8058 4384
rect 8122 4320 8138 4384
rect 8202 4320 8208 4384
rect 7892 4319 8208 4320
rect 14838 4384 15154 4385
rect 14838 4320 14844 4384
rect 14908 4320 14924 4384
rect 14988 4320 15004 4384
rect 15068 4320 15084 4384
rect 15148 4320 15154 4384
rect 14838 4319 15154 4320
rect 21784 4384 22100 4385
rect 21784 4320 21790 4384
rect 21854 4320 21870 4384
rect 21934 4320 21950 4384
rect 22014 4320 22030 4384
rect 22094 4320 22100 4384
rect 21784 4319 22100 4320
rect 28730 4384 29046 4385
rect 28730 4320 28736 4384
rect 28800 4320 28816 4384
rect 28880 4320 28896 4384
rect 28960 4320 28976 4384
rect 29040 4320 29046 4384
rect 28730 4319 29046 4320
rect 200 4178 800 4268
rect 2773 4178 2839 4181
rect 200 4176 2839 4178
rect 200 4120 2778 4176
rect 2834 4120 2839 4176
rect 200 4118 2839 4120
rect 200 4028 800 4118
rect 2773 4115 2839 4118
rect 29200 4028 29800 4268
rect 4419 3840 4735 3841
rect 4419 3776 4425 3840
rect 4489 3776 4505 3840
rect 4569 3776 4585 3840
rect 4649 3776 4665 3840
rect 4729 3776 4735 3840
rect 4419 3775 4735 3776
rect 11365 3840 11681 3841
rect 11365 3776 11371 3840
rect 11435 3776 11451 3840
rect 11515 3776 11531 3840
rect 11595 3776 11611 3840
rect 11675 3776 11681 3840
rect 11365 3775 11681 3776
rect 18311 3840 18627 3841
rect 18311 3776 18317 3840
rect 18381 3776 18397 3840
rect 18461 3776 18477 3840
rect 18541 3776 18557 3840
rect 18621 3776 18627 3840
rect 18311 3775 18627 3776
rect 25257 3840 25573 3841
rect 25257 3776 25263 3840
rect 25327 3776 25343 3840
rect 25407 3776 25423 3840
rect 25487 3776 25503 3840
rect 25567 3776 25573 3840
rect 25257 3775 25573 3776
rect 200 3498 800 3588
rect 2773 3498 2839 3501
rect 200 3496 2839 3498
rect 200 3440 2778 3496
rect 2834 3440 2839 3496
rect 200 3438 2839 3440
rect 200 3348 800 3438
rect 2773 3435 2839 3438
rect 26141 3498 26207 3501
rect 29200 3498 29800 3588
rect 26141 3496 29800 3498
rect 26141 3440 26146 3496
rect 26202 3440 29800 3496
rect 26141 3438 29800 3440
rect 26141 3435 26207 3438
rect 29200 3348 29800 3438
rect 7892 3296 8208 3297
rect 7892 3232 7898 3296
rect 7962 3232 7978 3296
rect 8042 3232 8058 3296
rect 8122 3232 8138 3296
rect 8202 3232 8208 3296
rect 7892 3231 8208 3232
rect 14838 3296 15154 3297
rect 14838 3232 14844 3296
rect 14908 3232 14924 3296
rect 14988 3232 15004 3296
rect 15068 3232 15084 3296
rect 15148 3232 15154 3296
rect 14838 3231 15154 3232
rect 21784 3296 22100 3297
rect 21784 3232 21790 3296
rect 21854 3232 21870 3296
rect 21934 3232 21950 3296
rect 22014 3232 22030 3296
rect 22094 3232 22100 3296
rect 21784 3231 22100 3232
rect 28730 3296 29046 3297
rect 28730 3232 28736 3296
rect 28800 3232 28816 3296
rect 28880 3232 28896 3296
rect 28960 3232 28976 3296
rect 29040 3232 29046 3296
rect 28730 3231 29046 3232
rect 200 2818 800 2908
rect 1577 2818 1643 2821
rect 200 2816 1643 2818
rect 200 2760 1582 2816
rect 1638 2760 1643 2816
rect 200 2758 1643 2760
rect 200 2668 800 2758
rect 1577 2755 1643 2758
rect 26141 2818 26207 2821
rect 29200 2818 29800 2908
rect 26141 2816 29800 2818
rect 26141 2760 26146 2816
rect 26202 2760 29800 2816
rect 26141 2758 29800 2760
rect 26141 2755 26207 2758
rect 4419 2752 4735 2753
rect 4419 2688 4425 2752
rect 4489 2688 4505 2752
rect 4569 2688 4585 2752
rect 4649 2688 4665 2752
rect 4729 2688 4735 2752
rect 4419 2687 4735 2688
rect 11365 2752 11681 2753
rect 11365 2688 11371 2752
rect 11435 2688 11451 2752
rect 11515 2688 11531 2752
rect 11595 2688 11611 2752
rect 11675 2688 11681 2752
rect 11365 2687 11681 2688
rect 18311 2752 18627 2753
rect 18311 2688 18317 2752
rect 18381 2688 18397 2752
rect 18461 2688 18477 2752
rect 18541 2688 18557 2752
rect 18621 2688 18627 2752
rect 18311 2687 18627 2688
rect 25257 2752 25573 2753
rect 25257 2688 25263 2752
rect 25327 2688 25343 2752
rect 25407 2688 25423 2752
rect 25487 2688 25503 2752
rect 25567 2688 25573 2752
rect 25257 2687 25573 2688
rect 29200 2668 29800 2758
rect 27429 2546 27495 2549
rect 27429 2544 29378 2546
rect 27429 2488 27434 2544
rect 27490 2488 29378 2544
rect 27429 2486 29378 2488
rect 27429 2483 27495 2486
rect 29318 2274 29378 2486
rect 29318 2228 29930 2274
rect 200 2138 800 2228
rect 29200 2214 29930 2228
rect 7892 2208 8208 2209
rect 7892 2144 7898 2208
rect 7962 2144 7978 2208
rect 8042 2144 8058 2208
rect 8122 2144 8138 2208
rect 8202 2144 8208 2208
rect 7892 2143 8208 2144
rect 14838 2208 15154 2209
rect 14838 2144 14844 2208
rect 14908 2144 14924 2208
rect 14988 2144 15004 2208
rect 15068 2144 15084 2208
rect 15148 2144 15154 2208
rect 14838 2143 15154 2144
rect 21784 2208 22100 2209
rect 21784 2144 21790 2208
rect 21854 2144 21870 2208
rect 21934 2144 21950 2208
rect 22014 2144 22030 2208
rect 22094 2144 22100 2208
rect 21784 2143 22100 2144
rect 28730 2208 29046 2209
rect 28730 2144 28736 2208
rect 28800 2144 28816 2208
rect 28880 2144 28896 2208
rect 28960 2144 28976 2208
rect 29040 2144 29046 2208
rect 28730 2143 29046 2144
rect 4061 2138 4127 2141
rect 200 2136 4127 2138
rect 200 2080 4066 2136
rect 4122 2080 4127 2136
rect 200 2078 4127 2080
rect 200 1988 800 2078
rect 4061 2075 4127 2078
rect 29200 2138 29800 2214
rect 29870 2138 29930 2214
rect 29200 2078 29930 2138
rect 29200 1988 29800 2078
rect 200 1458 800 1548
rect 3325 1458 3391 1461
rect 200 1456 3391 1458
rect 200 1400 3330 1456
rect 3386 1400 3391 1456
rect 200 1398 3391 1400
rect 200 1308 800 1398
rect 3325 1395 3391 1398
rect 27521 1458 27587 1461
rect 29200 1458 29800 1548
rect 27521 1456 29800 1458
rect 27521 1400 27526 1456
rect 27582 1400 29800 1456
rect 27521 1398 29800 1400
rect 27521 1395 27587 1398
rect 29200 1308 29800 1398
rect 200 628 800 868
rect 29200 -52 29800 188
<< via3 >>
rect 4425 47356 4489 47360
rect 4425 47300 4429 47356
rect 4429 47300 4485 47356
rect 4485 47300 4489 47356
rect 4425 47296 4489 47300
rect 4505 47356 4569 47360
rect 4505 47300 4509 47356
rect 4509 47300 4565 47356
rect 4565 47300 4569 47356
rect 4505 47296 4569 47300
rect 4585 47356 4649 47360
rect 4585 47300 4589 47356
rect 4589 47300 4645 47356
rect 4645 47300 4649 47356
rect 4585 47296 4649 47300
rect 4665 47356 4729 47360
rect 4665 47300 4669 47356
rect 4669 47300 4725 47356
rect 4725 47300 4729 47356
rect 4665 47296 4729 47300
rect 11371 47356 11435 47360
rect 11371 47300 11375 47356
rect 11375 47300 11431 47356
rect 11431 47300 11435 47356
rect 11371 47296 11435 47300
rect 11451 47356 11515 47360
rect 11451 47300 11455 47356
rect 11455 47300 11511 47356
rect 11511 47300 11515 47356
rect 11451 47296 11515 47300
rect 11531 47356 11595 47360
rect 11531 47300 11535 47356
rect 11535 47300 11591 47356
rect 11591 47300 11595 47356
rect 11531 47296 11595 47300
rect 11611 47356 11675 47360
rect 11611 47300 11615 47356
rect 11615 47300 11671 47356
rect 11671 47300 11675 47356
rect 11611 47296 11675 47300
rect 18317 47356 18381 47360
rect 18317 47300 18321 47356
rect 18321 47300 18377 47356
rect 18377 47300 18381 47356
rect 18317 47296 18381 47300
rect 18397 47356 18461 47360
rect 18397 47300 18401 47356
rect 18401 47300 18457 47356
rect 18457 47300 18461 47356
rect 18397 47296 18461 47300
rect 18477 47356 18541 47360
rect 18477 47300 18481 47356
rect 18481 47300 18537 47356
rect 18537 47300 18541 47356
rect 18477 47296 18541 47300
rect 18557 47356 18621 47360
rect 18557 47300 18561 47356
rect 18561 47300 18617 47356
rect 18617 47300 18621 47356
rect 18557 47296 18621 47300
rect 25263 47356 25327 47360
rect 25263 47300 25267 47356
rect 25267 47300 25323 47356
rect 25323 47300 25327 47356
rect 25263 47296 25327 47300
rect 25343 47356 25407 47360
rect 25343 47300 25347 47356
rect 25347 47300 25403 47356
rect 25403 47300 25407 47356
rect 25343 47296 25407 47300
rect 25423 47356 25487 47360
rect 25423 47300 25427 47356
rect 25427 47300 25483 47356
rect 25483 47300 25487 47356
rect 25423 47296 25487 47300
rect 25503 47356 25567 47360
rect 25503 47300 25507 47356
rect 25507 47300 25563 47356
rect 25563 47300 25567 47356
rect 25503 47296 25567 47300
rect 7898 46812 7962 46816
rect 7898 46756 7902 46812
rect 7902 46756 7958 46812
rect 7958 46756 7962 46812
rect 7898 46752 7962 46756
rect 7978 46812 8042 46816
rect 7978 46756 7982 46812
rect 7982 46756 8038 46812
rect 8038 46756 8042 46812
rect 7978 46752 8042 46756
rect 8058 46812 8122 46816
rect 8058 46756 8062 46812
rect 8062 46756 8118 46812
rect 8118 46756 8122 46812
rect 8058 46752 8122 46756
rect 8138 46812 8202 46816
rect 8138 46756 8142 46812
rect 8142 46756 8198 46812
rect 8198 46756 8202 46812
rect 8138 46752 8202 46756
rect 14844 46812 14908 46816
rect 14844 46756 14848 46812
rect 14848 46756 14904 46812
rect 14904 46756 14908 46812
rect 14844 46752 14908 46756
rect 14924 46812 14988 46816
rect 14924 46756 14928 46812
rect 14928 46756 14984 46812
rect 14984 46756 14988 46812
rect 14924 46752 14988 46756
rect 15004 46812 15068 46816
rect 15004 46756 15008 46812
rect 15008 46756 15064 46812
rect 15064 46756 15068 46812
rect 15004 46752 15068 46756
rect 15084 46812 15148 46816
rect 15084 46756 15088 46812
rect 15088 46756 15144 46812
rect 15144 46756 15148 46812
rect 15084 46752 15148 46756
rect 21790 46812 21854 46816
rect 21790 46756 21794 46812
rect 21794 46756 21850 46812
rect 21850 46756 21854 46812
rect 21790 46752 21854 46756
rect 21870 46812 21934 46816
rect 21870 46756 21874 46812
rect 21874 46756 21930 46812
rect 21930 46756 21934 46812
rect 21870 46752 21934 46756
rect 21950 46812 22014 46816
rect 21950 46756 21954 46812
rect 21954 46756 22010 46812
rect 22010 46756 22014 46812
rect 21950 46752 22014 46756
rect 22030 46812 22094 46816
rect 22030 46756 22034 46812
rect 22034 46756 22090 46812
rect 22090 46756 22094 46812
rect 22030 46752 22094 46756
rect 28736 46812 28800 46816
rect 28736 46756 28740 46812
rect 28740 46756 28796 46812
rect 28796 46756 28800 46812
rect 28736 46752 28800 46756
rect 28816 46812 28880 46816
rect 28816 46756 28820 46812
rect 28820 46756 28876 46812
rect 28876 46756 28880 46812
rect 28816 46752 28880 46756
rect 28896 46812 28960 46816
rect 28896 46756 28900 46812
rect 28900 46756 28956 46812
rect 28956 46756 28960 46812
rect 28896 46752 28960 46756
rect 28976 46812 29040 46816
rect 28976 46756 28980 46812
rect 28980 46756 29036 46812
rect 29036 46756 29040 46812
rect 28976 46752 29040 46756
rect 4425 46268 4489 46272
rect 4425 46212 4429 46268
rect 4429 46212 4485 46268
rect 4485 46212 4489 46268
rect 4425 46208 4489 46212
rect 4505 46268 4569 46272
rect 4505 46212 4509 46268
rect 4509 46212 4565 46268
rect 4565 46212 4569 46268
rect 4505 46208 4569 46212
rect 4585 46268 4649 46272
rect 4585 46212 4589 46268
rect 4589 46212 4645 46268
rect 4645 46212 4649 46268
rect 4585 46208 4649 46212
rect 4665 46268 4729 46272
rect 4665 46212 4669 46268
rect 4669 46212 4725 46268
rect 4725 46212 4729 46268
rect 4665 46208 4729 46212
rect 11371 46268 11435 46272
rect 11371 46212 11375 46268
rect 11375 46212 11431 46268
rect 11431 46212 11435 46268
rect 11371 46208 11435 46212
rect 11451 46268 11515 46272
rect 11451 46212 11455 46268
rect 11455 46212 11511 46268
rect 11511 46212 11515 46268
rect 11451 46208 11515 46212
rect 11531 46268 11595 46272
rect 11531 46212 11535 46268
rect 11535 46212 11591 46268
rect 11591 46212 11595 46268
rect 11531 46208 11595 46212
rect 11611 46268 11675 46272
rect 11611 46212 11615 46268
rect 11615 46212 11671 46268
rect 11671 46212 11675 46268
rect 11611 46208 11675 46212
rect 18317 46268 18381 46272
rect 18317 46212 18321 46268
rect 18321 46212 18377 46268
rect 18377 46212 18381 46268
rect 18317 46208 18381 46212
rect 18397 46268 18461 46272
rect 18397 46212 18401 46268
rect 18401 46212 18457 46268
rect 18457 46212 18461 46268
rect 18397 46208 18461 46212
rect 18477 46268 18541 46272
rect 18477 46212 18481 46268
rect 18481 46212 18537 46268
rect 18537 46212 18541 46268
rect 18477 46208 18541 46212
rect 18557 46268 18621 46272
rect 18557 46212 18561 46268
rect 18561 46212 18617 46268
rect 18617 46212 18621 46268
rect 18557 46208 18621 46212
rect 25263 46268 25327 46272
rect 25263 46212 25267 46268
rect 25267 46212 25323 46268
rect 25323 46212 25327 46268
rect 25263 46208 25327 46212
rect 25343 46268 25407 46272
rect 25343 46212 25347 46268
rect 25347 46212 25403 46268
rect 25403 46212 25407 46268
rect 25343 46208 25407 46212
rect 25423 46268 25487 46272
rect 25423 46212 25427 46268
rect 25427 46212 25483 46268
rect 25483 46212 25487 46268
rect 25423 46208 25487 46212
rect 25503 46268 25567 46272
rect 25503 46212 25507 46268
rect 25507 46212 25563 46268
rect 25563 46212 25567 46268
rect 25503 46208 25567 46212
rect 7898 45724 7962 45728
rect 7898 45668 7902 45724
rect 7902 45668 7958 45724
rect 7958 45668 7962 45724
rect 7898 45664 7962 45668
rect 7978 45724 8042 45728
rect 7978 45668 7982 45724
rect 7982 45668 8038 45724
rect 8038 45668 8042 45724
rect 7978 45664 8042 45668
rect 8058 45724 8122 45728
rect 8058 45668 8062 45724
rect 8062 45668 8118 45724
rect 8118 45668 8122 45724
rect 8058 45664 8122 45668
rect 8138 45724 8202 45728
rect 8138 45668 8142 45724
rect 8142 45668 8198 45724
rect 8198 45668 8202 45724
rect 8138 45664 8202 45668
rect 14844 45724 14908 45728
rect 14844 45668 14848 45724
rect 14848 45668 14904 45724
rect 14904 45668 14908 45724
rect 14844 45664 14908 45668
rect 14924 45724 14988 45728
rect 14924 45668 14928 45724
rect 14928 45668 14984 45724
rect 14984 45668 14988 45724
rect 14924 45664 14988 45668
rect 15004 45724 15068 45728
rect 15004 45668 15008 45724
rect 15008 45668 15064 45724
rect 15064 45668 15068 45724
rect 15004 45664 15068 45668
rect 15084 45724 15148 45728
rect 15084 45668 15088 45724
rect 15088 45668 15144 45724
rect 15144 45668 15148 45724
rect 15084 45664 15148 45668
rect 21790 45724 21854 45728
rect 21790 45668 21794 45724
rect 21794 45668 21850 45724
rect 21850 45668 21854 45724
rect 21790 45664 21854 45668
rect 21870 45724 21934 45728
rect 21870 45668 21874 45724
rect 21874 45668 21930 45724
rect 21930 45668 21934 45724
rect 21870 45664 21934 45668
rect 21950 45724 22014 45728
rect 21950 45668 21954 45724
rect 21954 45668 22010 45724
rect 22010 45668 22014 45724
rect 21950 45664 22014 45668
rect 22030 45724 22094 45728
rect 22030 45668 22034 45724
rect 22034 45668 22090 45724
rect 22090 45668 22094 45724
rect 22030 45664 22094 45668
rect 28736 45724 28800 45728
rect 28736 45668 28740 45724
rect 28740 45668 28796 45724
rect 28796 45668 28800 45724
rect 28736 45664 28800 45668
rect 28816 45724 28880 45728
rect 28816 45668 28820 45724
rect 28820 45668 28876 45724
rect 28876 45668 28880 45724
rect 28816 45664 28880 45668
rect 28896 45724 28960 45728
rect 28896 45668 28900 45724
rect 28900 45668 28956 45724
rect 28956 45668 28960 45724
rect 28896 45664 28960 45668
rect 28976 45724 29040 45728
rect 28976 45668 28980 45724
rect 28980 45668 29036 45724
rect 29036 45668 29040 45724
rect 28976 45664 29040 45668
rect 4425 45180 4489 45184
rect 4425 45124 4429 45180
rect 4429 45124 4485 45180
rect 4485 45124 4489 45180
rect 4425 45120 4489 45124
rect 4505 45180 4569 45184
rect 4505 45124 4509 45180
rect 4509 45124 4565 45180
rect 4565 45124 4569 45180
rect 4505 45120 4569 45124
rect 4585 45180 4649 45184
rect 4585 45124 4589 45180
rect 4589 45124 4645 45180
rect 4645 45124 4649 45180
rect 4585 45120 4649 45124
rect 4665 45180 4729 45184
rect 4665 45124 4669 45180
rect 4669 45124 4725 45180
rect 4725 45124 4729 45180
rect 4665 45120 4729 45124
rect 11371 45180 11435 45184
rect 11371 45124 11375 45180
rect 11375 45124 11431 45180
rect 11431 45124 11435 45180
rect 11371 45120 11435 45124
rect 11451 45180 11515 45184
rect 11451 45124 11455 45180
rect 11455 45124 11511 45180
rect 11511 45124 11515 45180
rect 11451 45120 11515 45124
rect 11531 45180 11595 45184
rect 11531 45124 11535 45180
rect 11535 45124 11591 45180
rect 11591 45124 11595 45180
rect 11531 45120 11595 45124
rect 11611 45180 11675 45184
rect 11611 45124 11615 45180
rect 11615 45124 11671 45180
rect 11671 45124 11675 45180
rect 11611 45120 11675 45124
rect 18317 45180 18381 45184
rect 18317 45124 18321 45180
rect 18321 45124 18377 45180
rect 18377 45124 18381 45180
rect 18317 45120 18381 45124
rect 18397 45180 18461 45184
rect 18397 45124 18401 45180
rect 18401 45124 18457 45180
rect 18457 45124 18461 45180
rect 18397 45120 18461 45124
rect 18477 45180 18541 45184
rect 18477 45124 18481 45180
rect 18481 45124 18537 45180
rect 18537 45124 18541 45180
rect 18477 45120 18541 45124
rect 18557 45180 18621 45184
rect 18557 45124 18561 45180
rect 18561 45124 18617 45180
rect 18617 45124 18621 45180
rect 18557 45120 18621 45124
rect 25263 45180 25327 45184
rect 25263 45124 25267 45180
rect 25267 45124 25323 45180
rect 25323 45124 25327 45180
rect 25263 45120 25327 45124
rect 25343 45180 25407 45184
rect 25343 45124 25347 45180
rect 25347 45124 25403 45180
rect 25403 45124 25407 45180
rect 25343 45120 25407 45124
rect 25423 45180 25487 45184
rect 25423 45124 25427 45180
rect 25427 45124 25483 45180
rect 25483 45124 25487 45180
rect 25423 45120 25487 45124
rect 25503 45180 25567 45184
rect 25503 45124 25507 45180
rect 25507 45124 25563 45180
rect 25563 45124 25567 45180
rect 25503 45120 25567 45124
rect 7898 44636 7962 44640
rect 7898 44580 7902 44636
rect 7902 44580 7958 44636
rect 7958 44580 7962 44636
rect 7898 44576 7962 44580
rect 7978 44636 8042 44640
rect 7978 44580 7982 44636
rect 7982 44580 8038 44636
rect 8038 44580 8042 44636
rect 7978 44576 8042 44580
rect 8058 44636 8122 44640
rect 8058 44580 8062 44636
rect 8062 44580 8118 44636
rect 8118 44580 8122 44636
rect 8058 44576 8122 44580
rect 8138 44636 8202 44640
rect 8138 44580 8142 44636
rect 8142 44580 8198 44636
rect 8198 44580 8202 44636
rect 8138 44576 8202 44580
rect 14844 44636 14908 44640
rect 14844 44580 14848 44636
rect 14848 44580 14904 44636
rect 14904 44580 14908 44636
rect 14844 44576 14908 44580
rect 14924 44636 14988 44640
rect 14924 44580 14928 44636
rect 14928 44580 14984 44636
rect 14984 44580 14988 44636
rect 14924 44576 14988 44580
rect 15004 44636 15068 44640
rect 15004 44580 15008 44636
rect 15008 44580 15064 44636
rect 15064 44580 15068 44636
rect 15004 44576 15068 44580
rect 15084 44636 15148 44640
rect 15084 44580 15088 44636
rect 15088 44580 15144 44636
rect 15144 44580 15148 44636
rect 15084 44576 15148 44580
rect 21790 44636 21854 44640
rect 21790 44580 21794 44636
rect 21794 44580 21850 44636
rect 21850 44580 21854 44636
rect 21790 44576 21854 44580
rect 21870 44636 21934 44640
rect 21870 44580 21874 44636
rect 21874 44580 21930 44636
rect 21930 44580 21934 44636
rect 21870 44576 21934 44580
rect 21950 44636 22014 44640
rect 21950 44580 21954 44636
rect 21954 44580 22010 44636
rect 22010 44580 22014 44636
rect 21950 44576 22014 44580
rect 22030 44636 22094 44640
rect 22030 44580 22034 44636
rect 22034 44580 22090 44636
rect 22090 44580 22094 44636
rect 22030 44576 22094 44580
rect 28736 44636 28800 44640
rect 28736 44580 28740 44636
rect 28740 44580 28796 44636
rect 28796 44580 28800 44636
rect 28736 44576 28800 44580
rect 28816 44636 28880 44640
rect 28816 44580 28820 44636
rect 28820 44580 28876 44636
rect 28876 44580 28880 44636
rect 28816 44576 28880 44580
rect 28896 44636 28960 44640
rect 28896 44580 28900 44636
rect 28900 44580 28956 44636
rect 28956 44580 28960 44636
rect 28896 44576 28960 44580
rect 28976 44636 29040 44640
rect 28976 44580 28980 44636
rect 28980 44580 29036 44636
rect 29036 44580 29040 44636
rect 28976 44576 29040 44580
rect 4425 44092 4489 44096
rect 4425 44036 4429 44092
rect 4429 44036 4485 44092
rect 4485 44036 4489 44092
rect 4425 44032 4489 44036
rect 4505 44092 4569 44096
rect 4505 44036 4509 44092
rect 4509 44036 4565 44092
rect 4565 44036 4569 44092
rect 4505 44032 4569 44036
rect 4585 44092 4649 44096
rect 4585 44036 4589 44092
rect 4589 44036 4645 44092
rect 4645 44036 4649 44092
rect 4585 44032 4649 44036
rect 4665 44092 4729 44096
rect 4665 44036 4669 44092
rect 4669 44036 4725 44092
rect 4725 44036 4729 44092
rect 4665 44032 4729 44036
rect 11371 44092 11435 44096
rect 11371 44036 11375 44092
rect 11375 44036 11431 44092
rect 11431 44036 11435 44092
rect 11371 44032 11435 44036
rect 11451 44092 11515 44096
rect 11451 44036 11455 44092
rect 11455 44036 11511 44092
rect 11511 44036 11515 44092
rect 11451 44032 11515 44036
rect 11531 44092 11595 44096
rect 11531 44036 11535 44092
rect 11535 44036 11591 44092
rect 11591 44036 11595 44092
rect 11531 44032 11595 44036
rect 11611 44092 11675 44096
rect 11611 44036 11615 44092
rect 11615 44036 11671 44092
rect 11671 44036 11675 44092
rect 11611 44032 11675 44036
rect 18317 44092 18381 44096
rect 18317 44036 18321 44092
rect 18321 44036 18377 44092
rect 18377 44036 18381 44092
rect 18317 44032 18381 44036
rect 18397 44092 18461 44096
rect 18397 44036 18401 44092
rect 18401 44036 18457 44092
rect 18457 44036 18461 44092
rect 18397 44032 18461 44036
rect 18477 44092 18541 44096
rect 18477 44036 18481 44092
rect 18481 44036 18537 44092
rect 18537 44036 18541 44092
rect 18477 44032 18541 44036
rect 18557 44092 18621 44096
rect 18557 44036 18561 44092
rect 18561 44036 18617 44092
rect 18617 44036 18621 44092
rect 18557 44032 18621 44036
rect 25263 44092 25327 44096
rect 25263 44036 25267 44092
rect 25267 44036 25323 44092
rect 25323 44036 25327 44092
rect 25263 44032 25327 44036
rect 25343 44092 25407 44096
rect 25343 44036 25347 44092
rect 25347 44036 25403 44092
rect 25403 44036 25407 44092
rect 25343 44032 25407 44036
rect 25423 44092 25487 44096
rect 25423 44036 25427 44092
rect 25427 44036 25483 44092
rect 25483 44036 25487 44092
rect 25423 44032 25487 44036
rect 25503 44092 25567 44096
rect 25503 44036 25507 44092
rect 25507 44036 25563 44092
rect 25563 44036 25567 44092
rect 25503 44032 25567 44036
rect 7898 43548 7962 43552
rect 7898 43492 7902 43548
rect 7902 43492 7958 43548
rect 7958 43492 7962 43548
rect 7898 43488 7962 43492
rect 7978 43548 8042 43552
rect 7978 43492 7982 43548
rect 7982 43492 8038 43548
rect 8038 43492 8042 43548
rect 7978 43488 8042 43492
rect 8058 43548 8122 43552
rect 8058 43492 8062 43548
rect 8062 43492 8118 43548
rect 8118 43492 8122 43548
rect 8058 43488 8122 43492
rect 8138 43548 8202 43552
rect 8138 43492 8142 43548
rect 8142 43492 8198 43548
rect 8198 43492 8202 43548
rect 8138 43488 8202 43492
rect 14844 43548 14908 43552
rect 14844 43492 14848 43548
rect 14848 43492 14904 43548
rect 14904 43492 14908 43548
rect 14844 43488 14908 43492
rect 14924 43548 14988 43552
rect 14924 43492 14928 43548
rect 14928 43492 14984 43548
rect 14984 43492 14988 43548
rect 14924 43488 14988 43492
rect 15004 43548 15068 43552
rect 15004 43492 15008 43548
rect 15008 43492 15064 43548
rect 15064 43492 15068 43548
rect 15004 43488 15068 43492
rect 15084 43548 15148 43552
rect 15084 43492 15088 43548
rect 15088 43492 15144 43548
rect 15144 43492 15148 43548
rect 15084 43488 15148 43492
rect 21790 43548 21854 43552
rect 21790 43492 21794 43548
rect 21794 43492 21850 43548
rect 21850 43492 21854 43548
rect 21790 43488 21854 43492
rect 21870 43548 21934 43552
rect 21870 43492 21874 43548
rect 21874 43492 21930 43548
rect 21930 43492 21934 43548
rect 21870 43488 21934 43492
rect 21950 43548 22014 43552
rect 21950 43492 21954 43548
rect 21954 43492 22010 43548
rect 22010 43492 22014 43548
rect 21950 43488 22014 43492
rect 22030 43548 22094 43552
rect 22030 43492 22034 43548
rect 22034 43492 22090 43548
rect 22090 43492 22094 43548
rect 22030 43488 22094 43492
rect 28736 43548 28800 43552
rect 28736 43492 28740 43548
rect 28740 43492 28796 43548
rect 28796 43492 28800 43548
rect 28736 43488 28800 43492
rect 28816 43548 28880 43552
rect 28816 43492 28820 43548
rect 28820 43492 28876 43548
rect 28876 43492 28880 43548
rect 28816 43488 28880 43492
rect 28896 43548 28960 43552
rect 28896 43492 28900 43548
rect 28900 43492 28956 43548
rect 28956 43492 28960 43548
rect 28896 43488 28960 43492
rect 28976 43548 29040 43552
rect 28976 43492 28980 43548
rect 28980 43492 29036 43548
rect 29036 43492 29040 43548
rect 28976 43488 29040 43492
rect 4425 43004 4489 43008
rect 4425 42948 4429 43004
rect 4429 42948 4485 43004
rect 4485 42948 4489 43004
rect 4425 42944 4489 42948
rect 4505 43004 4569 43008
rect 4505 42948 4509 43004
rect 4509 42948 4565 43004
rect 4565 42948 4569 43004
rect 4505 42944 4569 42948
rect 4585 43004 4649 43008
rect 4585 42948 4589 43004
rect 4589 42948 4645 43004
rect 4645 42948 4649 43004
rect 4585 42944 4649 42948
rect 4665 43004 4729 43008
rect 4665 42948 4669 43004
rect 4669 42948 4725 43004
rect 4725 42948 4729 43004
rect 4665 42944 4729 42948
rect 11371 43004 11435 43008
rect 11371 42948 11375 43004
rect 11375 42948 11431 43004
rect 11431 42948 11435 43004
rect 11371 42944 11435 42948
rect 11451 43004 11515 43008
rect 11451 42948 11455 43004
rect 11455 42948 11511 43004
rect 11511 42948 11515 43004
rect 11451 42944 11515 42948
rect 11531 43004 11595 43008
rect 11531 42948 11535 43004
rect 11535 42948 11591 43004
rect 11591 42948 11595 43004
rect 11531 42944 11595 42948
rect 11611 43004 11675 43008
rect 11611 42948 11615 43004
rect 11615 42948 11671 43004
rect 11671 42948 11675 43004
rect 11611 42944 11675 42948
rect 18317 43004 18381 43008
rect 18317 42948 18321 43004
rect 18321 42948 18377 43004
rect 18377 42948 18381 43004
rect 18317 42944 18381 42948
rect 18397 43004 18461 43008
rect 18397 42948 18401 43004
rect 18401 42948 18457 43004
rect 18457 42948 18461 43004
rect 18397 42944 18461 42948
rect 18477 43004 18541 43008
rect 18477 42948 18481 43004
rect 18481 42948 18537 43004
rect 18537 42948 18541 43004
rect 18477 42944 18541 42948
rect 18557 43004 18621 43008
rect 18557 42948 18561 43004
rect 18561 42948 18617 43004
rect 18617 42948 18621 43004
rect 18557 42944 18621 42948
rect 25263 43004 25327 43008
rect 25263 42948 25267 43004
rect 25267 42948 25323 43004
rect 25323 42948 25327 43004
rect 25263 42944 25327 42948
rect 25343 43004 25407 43008
rect 25343 42948 25347 43004
rect 25347 42948 25403 43004
rect 25403 42948 25407 43004
rect 25343 42944 25407 42948
rect 25423 43004 25487 43008
rect 25423 42948 25427 43004
rect 25427 42948 25483 43004
rect 25483 42948 25487 43004
rect 25423 42944 25487 42948
rect 25503 43004 25567 43008
rect 25503 42948 25507 43004
rect 25507 42948 25563 43004
rect 25563 42948 25567 43004
rect 25503 42944 25567 42948
rect 7898 42460 7962 42464
rect 7898 42404 7902 42460
rect 7902 42404 7958 42460
rect 7958 42404 7962 42460
rect 7898 42400 7962 42404
rect 7978 42460 8042 42464
rect 7978 42404 7982 42460
rect 7982 42404 8038 42460
rect 8038 42404 8042 42460
rect 7978 42400 8042 42404
rect 8058 42460 8122 42464
rect 8058 42404 8062 42460
rect 8062 42404 8118 42460
rect 8118 42404 8122 42460
rect 8058 42400 8122 42404
rect 8138 42460 8202 42464
rect 8138 42404 8142 42460
rect 8142 42404 8198 42460
rect 8198 42404 8202 42460
rect 8138 42400 8202 42404
rect 14844 42460 14908 42464
rect 14844 42404 14848 42460
rect 14848 42404 14904 42460
rect 14904 42404 14908 42460
rect 14844 42400 14908 42404
rect 14924 42460 14988 42464
rect 14924 42404 14928 42460
rect 14928 42404 14984 42460
rect 14984 42404 14988 42460
rect 14924 42400 14988 42404
rect 15004 42460 15068 42464
rect 15004 42404 15008 42460
rect 15008 42404 15064 42460
rect 15064 42404 15068 42460
rect 15004 42400 15068 42404
rect 15084 42460 15148 42464
rect 15084 42404 15088 42460
rect 15088 42404 15144 42460
rect 15144 42404 15148 42460
rect 15084 42400 15148 42404
rect 21790 42460 21854 42464
rect 21790 42404 21794 42460
rect 21794 42404 21850 42460
rect 21850 42404 21854 42460
rect 21790 42400 21854 42404
rect 21870 42460 21934 42464
rect 21870 42404 21874 42460
rect 21874 42404 21930 42460
rect 21930 42404 21934 42460
rect 21870 42400 21934 42404
rect 21950 42460 22014 42464
rect 21950 42404 21954 42460
rect 21954 42404 22010 42460
rect 22010 42404 22014 42460
rect 21950 42400 22014 42404
rect 22030 42460 22094 42464
rect 22030 42404 22034 42460
rect 22034 42404 22090 42460
rect 22090 42404 22094 42460
rect 22030 42400 22094 42404
rect 28736 42460 28800 42464
rect 28736 42404 28740 42460
rect 28740 42404 28796 42460
rect 28796 42404 28800 42460
rect 28736 42400 28800 42404
rect 28816 42460 28880 42464
rect 28816 42404 28820 42460
rect 28820 42404 28876 42460
rect 28876 42404 28880 42460
rect 28816 42400 28880 42404
rect 28896 42460 28960 42464
rect 28896 42404 28900 42460
rect 28900 42404 28956 42460
rect 28956 42404 28960 42460
rect 28896 42400 28960 42404
rect 28976 42460 29040 42464
rect 28976 42404 28980 42460
rect 28980 42404 29036 42460
rect 29036 42404 29040 42460
rect 28976 42400 29040 42404
rect 4425 41916 4489 41920
rect 4425 41860 4429 41916
rect 4429 41860 4485 41916
rect 4485 41860 4489 41916
rect 4425 41856 4489 41860
rect 4505 41916 4569 41920
rect 4505 41860 4509 41916
rect 4509 41860 4565 41916
rect 4565 41860 4569 41916
rect 4505 41856 4569 41860
rect 4585 41916 4649 41920
rect 4585 41860 4589 41916
rect 4589 41860 4645 41916
rect 4645 41860 4649 41916
rect 4585 41856 4649 41860
rect 4665 41916 4729 41920
rect 4665 41860 4669 41916
rect 4669 41860 4725 41916
rect 4725 41860 4729 41916
rect 4665 41856 4729 41860
rect 11371 41916 11435 41920
rect 11371 41860 11375 41916
rect 11375 41860 11431 41916
rect 11431 41860 11435 41916
rect 11371 41856 11435 41860
rect 11451 41916 11515 41920
rect 11451 41860 11455 41916
rect 11455 41860 11511 41916
rect 11511 41860 11515 41916
rect 11451 41856 11515 41860
rect 11531 41916 11595 41920
rect 11531 41860 11535 41916
rect 11535 41860 11591 41916
rect 11591 41860 11595 41916
rect 11531 41856 11595 41860
rect 11611 41916 11675 41920
rect 11611 41860 11615 41916
rect 11615 41860 11671 41916
rect 11671 41860 11675 41916
rect 11611 41856 11675 41860
rect 18317 41916 18381 41920
rect 18317 41860 18321 41916
rect 18321 41860 18377 41916
rect 18377 41860 18381 41916
rect 18317 41856 18381 41860
rect 18397 41916 18461 41920
rect 18397 41860 18401 41916
rect 18401 41860 18457 41916
rect 18457 41860 18461 41916
rect 18397 41856 18461 41860
rect 18477 41916 18541 41920
rect 18477 41860 18481 41916
rect 18481 41860 18537 41916
rect 18537 41860 18541 41916
rect 18477 41856 18541 41860
rect 18557 41916 18621 41920
rect 18557 41860 18561 41916
rect 18561 41860 18617 41916
rect 18617 41860 18621 41916
rect 18557 41856 18621 41860
rect 25263 41916 25327 41920
rect 25263 41860 25267 41916
rect 25267 41860 25323 41916
rect 25323 41860 25327 41916
rect 25263 41856 25327 41860
rect 25343 41916 25407 41920
rect 25343 41860 25347 41916
rect 25347 41860 25403 41916
rect 25403 41860 25407 41916
rect 25343 41856 25407 41860
rect 25423 41916 25487 41920
rect 25423 41860 25427 41916
rect 25427 41860 25483 41916
rect 25483 41860 25487 41916
rect 25423 41856 25487 41860
rect 25503 41916 25567 41920
rect 25503 41860 25507 41916
rect 25507 41860 25563 41916
rect 25563 41860 25567 41916
rect 25503 41856 25567 41860
rect 7898 41372 7962 41376
rect 7898 41316 7902 41372
rect 7902 41316 7958 41372
rect 7958 41316 7962 41372
rect 7898 41312 7962 41316
rect 7978 41372 8042 41376
rect 7978 41316 7982 41372
rect 7982 41316 8038 41372
rect 8038 41316 8042 41372
rect 7978 41312 8042 41316
rect 8058 41372 8122 41376
rect 8058 41316 8062 41372
rect 8062 41316 8118 41372
rect 8118 41316 8122 41372
rect 8058 41312 8122 41316
rect 8138 41372 8202 41376
rect 8138 41316 8142 41372
rect 8142 41316 8198 41372
rect 8198 41316 8202 41372
rect 8138 41312 8202 41316
rect 14844 41372 14908 41376
rect 14844 41316 14848 41372
rect 14848 41316 14904 41372
rect 14904 41316 14908 41372
rect 14844 41312 14908 41316
rect 14924 41372 14988 41376
rect 14924 41316 14928 41372
rect 14928 41316 14984 41372
rect 14984 41316 14988 41372
rect 14924 41312 14988 41316
rect 15004 41372 15068 41376
rect 15004 41316 15008 41372
rect 15008 41316 15064 41372
rect 15064 41316 15068 41372
rect 15004 41312 15068 41316
rect 15084 41372 15148 41376
rect 15084 41316 15088 41372
rect 15088 41316 15144 41372
rect 15144 41316 15148 41372
rect 15084 41312 15148 41316
rect 21790 41372 21854 41376
rect 21790 41316 21794 41372
rect 21794 41316 21850 41372
rect 21850 41316 21854 41372
rect 21790 41312 21854 41316
rect 21870 41372 21934 41376
rect 21870 41316 21874 41372
rect 21874 41316 21930 41372
rect 21930 41316 21934 41372
rect 21870 41312 21934 41316
rect 21950 41372 22014 41376
rect 21950 41316 21954 41372
rect 21954 41316 22010 41372
rect 22010 41316 22014 41372
rect 21950 41312 22014 41316
rect 22030 41372 22094 41376
rect 22030 41316 22034 41372
rect 22034 41316 22090 41372
rect 22090 41316 22094 41372
rect 22030 41312 22094 41316
rect 28736 41372 28800 41376
rect 28736 41316 28740 41372
rect 28740 41316 28796 41372
rect 28796 41316 28800 41372
rect 28736 41312 28800 41316
rect 28816 41372 28880 41376
rect 28816 41316 28820 41372
rect 28820 41316 28876 41372
rect 28876 41316 28880 41372
rect 28816 41312 28880 41316
rect 28896 41372 28960 41376
rect 28896 41316 28900 41372
rect 28900 41316 28956 41372
rect 28956 41316 28960 41372
rect 28896 41312 28960 41316
rect 28976 41372 29040 41376
rect 28976 41316 28980 41372
rect 28980 41316 29036 41372
rect 29036 41316 29040 41372
rect 28976 41312 29040 41316
rect 4425 40828 4489 40832
rect 4425 40772 4429 40828
rect 4429 40772 4485 40828
rect 4485 40772 4489 40828
rect 4425 40768 4489 40772
rect 4505 40828 4569 40832
rect 4505 40772 4509 40828
rect 4509 40772 4565 40828
rect 4565 40772 4569 40828
rect 4505 40768 4569 40772
rect 4585 40828 4649 40832
rect 4585 40772 4589 40828
rect 4589 40772 4645 40828
rect 4645 40772 4649 40828
rect 4585 40768 4649 40772
rect 4665 40828 4729 40832
rect 4665 40772 4669 40828
rect 4669 40772 4725 40828
rect 4725 40772 4729 40828
rect 4665 40768 4729 40772
rect 11371 40828 11435 40832
rect 11371 40772 11375 40828
rect 11375 40772 11431 40828
rect 11431 40772 11435 40828
rect 11371 40768 11435 40772
rect 11451 40828 11515 40832
rect 11451 40772 11455 40828
rect 11455 40772 11511 40828
rect 11511 40772 11515 40828
rect 11451 40768 11515 40772
rect 11531 40828 11595 40832
rect 11531 40772 11535 40828
rect 11535 40772 11591 40828
rect 11591 40772 11595 40828
rect 11531 40768 11595 40772
rect 11611 40828 11675 40832
rect 11611 40772 11615 40828
rect 11615 40772 11671 40828
rect 11671 40772 11675 40828
rect 11611 40768 11675 40772
rect 18317 40828 18381 40832
rect 18317 40772 18321 40828
rect 18321 40772 18377 40828
rect 18377 40772 18381 40828
rect 18317 40768 18381 40772
rect 18397 40828 18461 40832
rect 18397 40772 18401 40828
rect 18401 40772 18457 40828
rect 18457 40772 18461 40828
rect 18397 40768 18461 40772
rect 18477 40828 18541 40832
rect 18477 40772 18481 40828
rect 18481 40772 18537 40828
rect 18537 40772 18541 40828
rect 18477 40768 18541 40772
rect 18557 40828 18621 40832
rect 18557 40772 18561 40828
rect 18561 40772 18617 40828
rect 18617 40772 18621 40828
rect 18557 40768 18621 40772
rect 25263 40828 25327 40832
rect 25263 40772 25267 40828
rect 25267 40772 25323 40828
rect 25323 40772 25327 40828
rect 25263 40768 25327 40772
rect 25343 40828 25407 40832
rect 25343 40772 25347 40828
rect 25347 40772 25403 40828
rect 25403 40772 25407 40828
rect 25343 40768 25407 40772
rect 25423 40828 25487 40832
rect 25423 40772 25427 40828
rect 25427 40772 25483 40828
rect 25483 40772 25487 40828
rect 25423 40768 25487 40772
rect 25503 40828 25567 40832
rect 25503 40772 25507 40828
rect 25507 40772 25563 40828
rect 25563 40772 25567 40828
rect 25503 40768 25567 40772
rect 7898 40284 7962 40288
rect 7898 40228 7902 40284
rect 7902 40228 7958 40284
rect 7958 40228 7962 40284
rect 7898 40224 7962 40228
rect 7978 40284 8042 40288
rect 7978 40228 7982 40284
rect 7982 40228 8038 40284
rect 8038 40228 8042 40284
rect 7978 40224 8042 40228
rect 8058 40284 8122 40288
rect 8058 40228 8062 40284
rect 8062 40228 8118 40284
rect 8118 40228 8122 40284
rect 8058 40224 8122 40228
rect 8138 40284 8202 40288
rect 8138 40228 8142 40284
rect 8142 40228 8198 40284
rect 8198 40228 8202 40284
rect 8138 40224 8202 40228
rect 14844 40284 14908 40288
rect 14844 40228 14848 40284
rect 14848 40228 14904 40284
rect 14904 40228 14908 40284
rect 14844 40224 14908 40228
rect 14924 40284 14988 40288
rect 14924 40228 14928 40284
rect 14928 40228 14984 40284
rect 14984 40228 14988 40284
rect 14924 40224 14988 40228
rect 15004 40284 15068 40288
rect 15004 40228 15008 40284
rect 15008 40228 15064 40284
rect 15064 40228 15068 40284
rect 15004 40224 15068 40228
rect 15084 40284 15148 40288
rect 15084 40228 15088 40284
rect 15088 40228 15144 40284
rect 15144 40228 15148 40284
rect 15084 40224 15148 40228
rect 21790 40284 21854 40288
rect 21790 40228 21794 40284
rect 21794 40228 21850 40284
rect 21850 40228 21854 40284
rect 21790 40224 21854 40228
rect 21870 40284 21934 40288
rect 21870 40228 21874 40284
rect 21874 40228 21930 40284
rect 21930 40228 21934 40284
rect 21870 40224 21934 40228
rect 21950 40284 22014 40288
rect 21950 40228 21954 40284
rect 21954 40228 22010 40284
rect 22010 40228 22014 40284
rect 21950 40224 22014 40228
rect 22030 40284 22094 40288
rect 22030 40228 22034 40284
rect 22034 40228 22090 40284
rect 22090 40228 22094 40284
rect 22030 40224 22094 40228
rect 28736 40284 28800 40288
rect 28736 40228 28740 40284
rect 28740 40228 28796 40284
rect 28796 40228 28800 40284
rect 28736 40224 28800 40228
rect 28816 40284 28880 40288
rect 28816 40228 28820 40284
rect 28820 40228 28876 40284
rect 28876 40228 28880 40284
rect 28816 40224 28880 40228
rect 28896 40284 28960 40288
rect 28896 40228 28900 40284
rect 28900 40228 28956 40284
rect 28956 40228 28960 40284
rect 28896 40224 28960 40228
rect 28976 40284 29040 40288
rect 28976 40228 28980 40284
rect 28980 40228 29036 40284
rect 29036 40228 29040 40284
rect 28976 40224 29040 40228
rect 4425 39740 4489 39744
rect 4425 39684 4429 39740
rect 4429 39684 4485 39740
rect 4485 39684 4489 39740
rect 4425 39680 4489 39684
rect 4505 39740 4569 39744
rect 4505 39684 4509 39740
rect 4509 39684 4565 39740
rect 4565 39684 4569 39740
rect 4505 39680 4569 39684
rect 4585 39740 4649 39744
rect 4585 39684 4589 39740
rect 4589 39684 4645 39740
rect 4645 39684 4649 39740
rect 4585 39680 4649 39684
rect 4665 39740 4729 39744
rect 4665 39684 4669 39740
rect 4669 39684 4725 39740
rect 4725 39684 4729 39740
rect 4665 39680 4729 39684
rect 11371 39740 11435 39744
rect 11371 39684 11375 39740
rect 11375 39684 11431 39740
rect 11431 39684 11435 39740
rect 11371 39680 11435 39684
rect 11451 39740 11515 39744
rect 11451 39684 11455 39740
rect 11455 39684 11511 39740
rect 11511 39684 11515 39740
rect 11451 39680 11515 39684
rect 11531 39740 11595 39744
rect 11531 39684 11535 39740
rect 11535 39684 11591 39740
rect 11591 39684 11595 39740
rect 11531 39680 11595 39684
rect 11611 39740 11675 39744
rect 11611 39684 11615 39740
rect 11615 39684 11671 39740
rect 11671 39684 11675 39740
rect 11611 39680 11675 39684
rect 18317 39740 18381 39744
rect 18317 39684 18321 39740
rect 18321 39684 18377 39740
rect 18377 39684 18381 39740
rect 18317 39680 18381 39684
rect 18397 39740 18461 39744
rect 18397 39684 18401 39740
rect 18401 39684 18457 39740
rect 18457 39684 18461 39740
rect 18397 39680 18461 39684
rect 18477 39740 18541 39744
rect 18477 39684 18481 39740
rect 18481 39684 18537 39740
rect 18537 39684 18541 39740
rect 18477 39680 18541 39684
rect 18557 39740 18621 39744
rect 18557 39684 18561 39740
rect 18561 39684 18617 39740
rect 18617 39684 18621 39740
rect 18557 39680 18621 39684
rect 25263 39740 25327 39744
rect 25263 39684 25267 39740
rect 25267 39684 25323 39740
rect 25323 39684 25327 39740
rect 25263 39680 25327 39684
rect 25343 39740 25407 39744
rect 25343 39684 25347 39740
rect 25347 39684 25403 39740
rect 25403 39684 25407 39740
rect 25343 39680 25407 39684
rect 25423 39740 25487 39744
rect 25423 39684 25427 39740
rect 25427 39684 25483 39740
rect 25483 39684 25487 39740
rect 25423 39680 25487 39684
rect 25503 39740 25567 39744
rect 25503 39684 25507 39740
rect 25507 39684 25563 39740
rect 25563 39684 25567 39740
rect 25503 39680 25567 39684
rect 7898 39196 7962 39200
rect 7898 39140 7902 39196
rect 7902 39140 7958 39196
rect 7958 39140 7962 39196
rect 7898 39136 7962 39140
rect 7978 39196 8042 39200
rect 7978 39140 7982 39196
rect 7982 39140 8038 39196
rect 8038 39140 8042 39196
rect 7978 39136 8042 39140
rect 8058 39196 8122 39200
rect 8058 39140 8062 39196
rect 8062 39140 8118 39196
rect 8118 39140 8122 39196
rect 8058 39136 8122 39140
rect 8138 39196 8202 39200
rect 8138 39140 8142 39196
rect 8142 39140 8198 39196
rect 8198 39140 8202 39196
rect 8138 39136 8202 39140
rect 14844 39196 14908 39200
rect 14844 39140 14848 39196
rect 14848 39140 14904 39196
rect 14904 39140 14908 39196
rect 14844 39136 14908 39140
rect 14924 39196 14988 39200
rect 14924 39140 14928 39196
rect 14928 39140 14984 39196
rect 14984 39140 14988 39196
rect 14924 39136 14988 39140
rect 15004 39196 15068 39200
rect 15004 39140 15008 39196
rect 15008 39140 15064 39196
rect 15064 39140 15068 39196
rect 15004 39136 15068 39140
rect 15084 39196 15148 39200
rect 15084 39140 15088 39196
rect 15088 39140 15144 39196
rect 15144 39140 15148 39196
rect 15084 39136 15148 39140
rect 21790 39196 21854 39200
rect 21790 39140 21794 39196
rect 21794 39140 21850 39196
rect 21850 39140 21854 39196
rect 21790 39136 21854 39140
rect 21870 39196 21934 39200
rect 21870 39140 21874 39196
rect 21874 39140 21930 39196
rect 21930 39140 21934 39196
rect 21870 39136 21934 39140
rect 21950 39196 22014 39200
rect 21950 39140 21954 39196
rect 21954 39140 22010 39196
rect 22010 39140 22014 39196
rect 21950 39136 22014 39140
rect 22030 39196 22094 39200
rect 22030 39140 22034 39196
rect 22034 39140 22090 39196
rect 22090 39140 22094 39196
rect 22030 39136 22094 39140
rect 28736 39196 28800 39200
rect 28736 39140 28740 39196
rect 28740 39140 28796 39196
rect 28796 39140 28800 39196
rect 28736 39136 28800 39140
rect 28816 39196 28880 39200
rect 28816 39140 28820 39196
rect 28820 39140 28876 39196
rect 28876 39140 28880 39196
rect 28816 39136 28880 39140
rect 28896 39196 28960 39200
rect 28896 39140 28900 39196
rect 28900 39140 28956 39196
rect 28956 39140 28960 39196
rect 28896 39136 28960 39140
rect 28976 39196 29040 39200
rect 28976 39140 28980 39196
rect 28980 39140 29036 39196
rect 29036 39140 29040 39196
rect 28976 39136 29040 39140
rect 4425 38652 4489 38656
rect 4425 38596 4429 38652
rect 4429 38596 4485 38652
rect 4485 38596 4489 38652
rect 4425 38592 4489 38596
rect 4505 38652 4569 38656
rect 4505 38596 4509 38652
rect 4509 38596 4565 38652
rect 4565 38596 4569 38652
rect 4505 38592 4569 38596
rect 4585 38652 4649 38656
rect 4585 38596 4589 38652
rect 4589 38596 4645 38652
rect 4645 38596 4649 38652
rect 4585 38592 4649 38596
rect 4665 38652 4729 38656
rect 4665 38596 4669 38652
rect 4669 38596 4725 38652
rect 4725 38596 4729 38652
rect 4665 38592 4729 38596
rect 11371 38652 11435 38656
rect 11371 38596 11375 38652
rect 11375 38596 11431 38652
rect 11431 38596 11435 38652
rect 11371 38592 11435 38596
rect 11451 38652 11515 38656
rect 11451 38596 11455 38652
rect 11455 38596 11511 38652
rect 11511 38596 11515 38652
rect 11451 38592 11515 38596
rect 11531 38652 11595 38656
rect 11531 38596 11535 38652
rect 11535 38596 11591 38652
rect 11591 38596 11595 38652
rect 11531 38592 11595 38596
rect 11611 38652 11675 38656
rect 11611 38596 11615 38652
rect 11615 38596 11671 38652
rect 11671 38596 11675 38652
rect 11611 38592 11675 38596
rect 18317 38652 18381 38656
rect 18317 38596 18321 38652
rect 18321 38596 18377 38652
rect 18377 38596 18381 38652
rect 18317 38592 18381 38596
rect 18397 38652 18461 38656
rect 18397 38596 18401 38652
rect 18401 38596 18457 38652
rect 18457 38596 18461 38652
rect 18397 38592 18461 38596
rect 18477 38652 18541 38656
rect 18477 38596 18481 38652
rect 18481 38596 18537 38652
rect 18537 38596 18541 38652
rect 18477 38592 18541 38596
rect 18557 38652 18621 38656
rect 18557 38596 18561 38652
rect 18561 38596 18617 38652
rect 18617 38596 18621 38652
rect 18557 38592 18621 38596
rect 25263 38652 25327 38656
rect 25263 38596 25267 38652
rect 25267 38596 25323 38652
rect 25323 38596 25327 38652
rect 25263 38592 25327 38596
rect 25343 38652 25407 38656
rect 25343 38596 25347 38652
rect 25347 38596 25403 38652
rect 25403 38596 25407 38652
rect 25343 38592 25407 38596
rect 25423 38652 25487 38656
rect 25423 38596 25427 38652
rect 25427 38596 25483 38652
rect 25483 38596 25487 38652
rect 25423 38592 25487 38596
rect 25503 38652 25567 38656
rect 25503 38596 25507 38652
rect 25507 38596 25563 38652
rect 25563 38596 25567 38652
rect 25503 38592 25567 38596
rect 7898 38108 7962 38112
rect 7898 38052 7902 38108
rect 7902 38052 7958 38108
rect 7958 38052 7962 38108
rect 7898 38048 7962 38052
rect 7978 38108 8042 38112
rect 7978 38052 7982 38108
rect 7982 38052 8038 38108
rect 8038 38052 8042 38108
rect 7978 38048 8042 38052
rect 8058 38108 8122 38112
rect 8058 38052 8062 38108
rect 8062 38052 8118 38108
rect 8118 38052 8122 38108
rect 8058 38048 8122 38052
rect 8138 38108 8202 38112
rect 8138 38052 8142 38108
rect 8142 38052 8198 38108
rect 8198 38052 8202 38108
rect 8138 38048 8202 38052
rect 14844 38108 14908 38112
rect 14844 38052 14848 38108
rect 14848 38052 14904 38108
rect 14904 38052 14908 38108
rect 14844 38048 14908 38052
rect 14924 38108 14988 38112
rect 14924 38052 14928 38108
rect 14928 38052 14984 38108
rect 14984 38052 14988 38108
rect 14924 38048 14988 38052
rect 15004 38108 15068 38112
rect 15004 38052 15008 38108
rect 15008 38052 15064 38108
rect 15064 38052 15068 38108
rect 15004 38048 15068 38052
rect 15084 38108 15148 38112
rect 15084 38052 15088 38108
rect 15088 38052 15144 38108
rect 15144 38052 15148 38108
rect 15084 38048 15148 38052
rect 21790 38108 21854 38112
rect 21790 38052 21794 38108
rect 21794 38052 21850 38108
rect 21850 38052 21854 38108
rect 21790 38048 21854 38052
rect 21870 38108 21934 38112
rect 21870 38052 21874 38108
rect 21874 38052 21930 38108
rect 21930 38052 21934 38108
rect 21870 38048 21934 38052
rect 21950 38108 22014 38112
rect 21950 38052 21954 38108
rect 21954 38052 22010 38108
rect 22010 38052 22014 38108
rect 21950 38048 22014 38052
rect 22030 38108 22094 38112
rect 22030 38052 22034 38108
rect 22034 38052 22090 38108
rect 22090 38052 22094 38108
rect 22030 38048 22094 38052
rect 28736 38108 28800 38112
rect 28736 38052 28740 38108
rect 28740 38052 28796 38108
rect 28796 38052 28800 38108
rect 28736 38048 28800 38052
rect 28816 38108 28880 38112
rect 28816 38052 28820 38108
rect 28820 38052 28876 38108
rect 28876 38052 28880 38108
rect 28816 38048 28880 38052
rect 28896 38108 28960 38112
rect 28896 38052 28900 38108
rect 28900 38052 28956 38108
rect 28956 38052 28960 38108
rect 28896 38048 28960 38052
rect 28976 38108 29040 38112
rect 28976 38052 28980 38108
rect 28980 38052 29036 38108
rect 29036 38052 29040 38108
rect 28976 38048 29040 38052
rect 4425 37564 4489 37568
rect 4425 37508 4429 37564
rect 4429 37508 4485 37564
rect 4485 37508 4489 37564
rect 4425 37504 4489 37508
rect 4505 37564 4569 37568
rect 4505 37508 4509 37564
rect 4509 37508 4565 37564
rect 4565 37508 4569 37564
rect 4505 37504 4569 37508
rect 4585 37564 4649 37568
rect 4585 37508 4589 37564
rect 4589 37508 4645 37564
rect 4645 37508 4649 37564
rect 4585 37504 4649 37508
rect 4665 37564 4729 37568
rect 4665 37508 4669 37564
rect 4669 37508 4725 37564
rect 4725 37508 4729 37564
rect 4665 37504 4729 37508
rect 11371 37564 11435 37568
rect 11371 37508 11375 37564
rect 11375 37508 11431 37564
rect 11431 37508 11435 37564
rect 11371 37504 11435 37508
rect 11451 37564 11515 37568
rect 11451 37508 11455 37564
rect 11455 37508 11511 37564
rect 11511 37508 11515 37564
rect 11451 37504 11515 37508
rect 11531 37564 11595 37568
rect 11531 37508 11535 37564
rect 11535 37508 11591 37564
rect 11591 37508 11595 37564
rect 11531 37504 11595 37508
rect 11611 37564 11675 37568
rect 11611 37508 11615 37564
rect 11615 37508 11671 37564
rect 11671 37508 11675 37564
rect 11611 37504 11675 37508
rect 18317 37564 18381 37568
rect 18317 37508 18321 37564
rect 18321 37508 18377 37564
rect 18377 37508 18381 37564
rect 18317 37504 18381 37508
rect 18397 37564 18461 37568
rect 18397 37508 18401 37564
rect 18401 37508 18457 37564
rect 18457 37508 18461 37564
rect 18397 37504 18461 37508
rect 18477 37564 18541 37568
rect 18477 37508 18481 37564
rect 18481 37508 18537 37564
rect 18537 37508 18541 37564
rect 18477 37504 18541 37508
rect 18557 37564 18621 37568
rect 18557 37508 18561 37564
rect 18561 37508 18617 37564
rect 18617 37508 18621 37564
rect 18557 37504 18621 37508
rect 25263 37564 25327 37568
rect 25263 37508 25267 37564
rect 25267 37508 25323 37564
rect 25323 37508 25327 37564
rect 25263 37504 25327 37508
rect 25343 37564 25407 37568
rect 25343 37508 25347 37564
rect 25347 37508 25403 37564
rect 25403 37508 25407 37564
rect 25343 37504 25407 37508
rect 25423 37564 25487 37568
rect 25423 37508 25427 37564
rect 25427 37508 25483 37564
rect 25483 37508 25487 37564
rect 25423 37504 25487 37508
rect 25503 37564 25567 37568
rect 25503 37508 25507 37564
rect 25507 37508 25563 37564
rect 25563 37508 25567 37564
rect 25503 37504 25567 37508
rect 7898 37020 7962 37024
rect 7898 36964 7902 37020
rect 7902 36964 7958 37020
rect 7958 36964 7962 37020
rect 7898 36960 7962 36964
rect 7978 37020 8042 37024
rect 7978 36964 7982 37020
rect 7982 36964 8038 37020
rect 8038 36964 8042 37020
rect 7978 36960 8042 36964
rect 8058 37020 8122 37024
rect 8058 36964 8062 37020
rect 8062 36964 8118 37020
rect 8118 36964 8122 37020
rect 8058 36960 8122 36964
rect 8138 37020 8202 37024
rect 8138 36964 8142 37020
rect 8142 36964 8198 37020
rect 8198 36964 8202 37020
rect 8138 36960 8202 36964
rect 14844 37020 14908 37024
rect 14844 36964 14848 37020
rect 14848 36964 14904 37020
rect 14904 36964 14908 37020
rect 14844 36960 14908 36964
rect 14924 37020 14988 37024
rect 14924 36964 14928 37020
rect 14928 36964 14984 37020
rect 14984 36964 14988 37020
rect 14924 36960 14988 36964
rect 15004 37020 15068 37024
rect 15004 36964 15008 37020
rect 15008 36964 15064 37020
rect 15064 36964 15068 37020
rect 15004 36960 15068 36964
rect 15084 37020 15148 37024
rect 15084 36964 15088 37020
rect 15088 36964 15144 37020
rect 15144 36964 15148 37020
rect 15084 36960 15148 36964
rect 21790 37020 21854 37024
rect 21790 36964 21794 37020
rect 21794 36964 21850 37020
rect 21850 36964 21854 37020
rect 21790 36960 21854 36964
rect 21870 37020 21934 37024
rect 21870 36964 21874 37020
rect 21874 36964 21930 37020
rect 21930 36964 21934 37020
rect 21870 36960 21934 36964
rect 21950 37020 22014 37024
rect 21950 36964 21954 37020
rect 21954 36964 22010 37020
rect 22010 36964 22014 37020
rect 21950 36960 22014 36964
rect 22030 37020 22094 37024
rect 22030 36964 22034 37020
rect 22034 36964 22090 37020
rect 22090 36964 22094 37020
rect 22030 36960 22094 36964
rect 28736 37020 28800 37024
rect 28736 36964 28740 37020
rect 28740 36964 28796 37020
rect 28796 36964 28800 37020
rect 28736 36960 28800 36964
rect 28816 37020 28880 37024
rect 28816 36964 28820 37020
rect 28820 36964 28876 37020
rect 28876 36964 28880 37020
rect 28816 36960 28880 36964
rect 28896 37020 28960 37024
rect 28896 36964 28900 37020
rect 28900 36964 28956 37020
rect 28956 36964 28960 37020
rect 28896 36960 28960 36964
rect 28976 37020 29040 37024
rect 28976 36964 28980 37020
rect 28980 36964 29036 37020
rect 29036 36964 29040 37020
rect 28976 36960 29040 36964
rect 4425 36476 4489 36480
rect 4425 36420 4429 36476
rect 4429 36420 4485 36476
rect 4485 36420 4489 36476
rect 4425 36416 4489 36420
rect 4505 36476 4569 36480
rect 4505 36420 4509 36476
rect 4509 36420 4565 36476
rect 4565 36420 4569 36476
rect 4505 36416 4569 36420
rect 4585 36476 4649 36480
rect 4585 36420 4589 36476
rect 4589 36420 4645 36476
rect 4645 36420 4649 36476
rect 4585 36416 4649 36420
rect 4665 36476 4729 36480
rect 4665 36420 4669 36476
rect 4669 36420 4725 36476
rect 4725 36420 4729 36476
rect 4665 36416 4729 36420
rect 11371 36476 11435 36480
rect 11371 36420 11375 36476
rect 11375 36420 11431 36476
rect 11431 36420 11435 36476
rect 11371 36416 11435 36420
rect 11451 36476 11515 36480
rect 11451 36420 11455 36476
rect 11455 36420 11511 36476
rect 11511 36420 11515 36476
rect 11451 36416 11515 36420
rect 11531 36476 11595 36480
rect 11531 36420 11535 36476
rect 11535 36420 11591 36476
rect 11591 36420 11595 36476
rect 11531 36416 11595 36420
rect 11611 36476 11675 36480
rect 11611 36420 11615 36476
rect 11615 36420 11671 36476
rect 11671 36420 11675 36476
rect 11611 36416 11675 36420
rect 18317 36476 18381 36480
rect 18317 36420 18321 36476
rect 18321 36420 18377 36476
rect 18377 36420 18381 36476
rect 18317 36416 18381 36420
rect 18397 36476 18461 36480
rect 18397 36420 18401 36476
rect 18401 36420 18457 36476
rect 18457 36420 18461 36476
rect 18397 36416 18461 36420
rect 18477 36476 18541 36480
rect 18477 36420 18481 36476
rect 18481 36420 18537 36476
rect 18537 36420 18541 36476
rect 18477 36416 18541 36420
rect 18557 36476 18621 36480
rect 18557 36420 18561 36476
rect 18561 36420 18617 36476
rect 18617 36420 18621 36476
rect 18557 36416 18621 36420
rect 25263 36476 25327 36480
rect 25263 36420 25267 36476
rect 25267 36420 25323 36476
rect 25323 36420 25327 36476
rect 25263 36416 25327 36420
rect 25343 36476 25407 36480
rect 25343 36420 25347 36476
rect 25347 36420 25403 36476
rect 25403 36420 25407 36476
rect 25343 36416 25407 36420
rect 25423 36476 25487 36480
rect 25423 36420 25427 36476
rect 25427 36420 25483 36476
rect 25483 36420 25487 36476
rect 25423 36416 25487 36420
rect 25503 36476 25567 36480
rect 25503 36420 25507 36476
rect 25507 36420 25563 36476
rect 25563 36420 25567 36476
rect 25503 36416 25567 36420
rect 7898 35932 7962 35936
rect 7898 35876 7902 35932
rect 7902 35876 7958 35932
rect 7958 35876 7962 35932
rect 7898 35872 7962 35876
rect 7978 35932 8042 35936
rect 7978 35876 7982 35932
rect 7982 35876 8038 35932
rect 8038 35876 8042 35932
rect 7978 35872 8042 35876
rect 8058 35932 8122 35936
rect 8058 35876 8062 35932
rect 8062 35876 8118 35932
rect 8118 35876 8122 35932
rect 8058 35872 8122 35876
rect 8138 35932 8202 35936
rect 8138 35876 8142 35932
rect 8142 35876 8198 35932
rect 8198 35876 8202 35932
rect 8138 35872 8202 35876
rect 14844 35932 14908 35936
rect 14844 35876 14848 35932
rect 14848 35876 14904 35932
rect 14904 35876 14908 35932
rect 14844 35872 14908 35876
rect 14924 35932 14988 35936
rect 14924 35876 14928 35932
rect 14928 35876 14984 35932
rect 14984 35876 14988 35932
rect 14924 35872 14988 35876
rect 15004 35932 15068 35936
rect 15004 35876 15008 35932
rect 15008 35876 15064 35932
rect 15064 35876 15068 35932
rect 15004 35872 15068 35876
rect 15084 35932 15148 35936
rect 15084 35876 15088 35932
rect 15088 35876 15144 35932
rect 15144 35876 15148 35932
rect 15084 35872 15148 35876
rect 21790 35932 21854 35936
rect 21790 35876 21794 35932
rect 21794 35876 21850 35932
rect 21850 35876 21854 35932
rect 21790 35872 21854 35876
rect 21870 35932 21934 35936
rect 21870 35876 21874 35932
rect 21874 35876 21930 35932
rect 21930 35876 21934 35932
rect 21870 35872 21934 35876
rect 21950 35932 22014 35936
rect 21950 35876 21954 35932
rect 21954 35876 22010 35932
rect 22010 35876 22014 35932
rect 21950 35872 22014 35876
rect 22030 35932 22094 35936
rect 22030 35876 22034 35932
rect 22034 35876 22090 35932
rect 22090 35876 22094 35932
rect 22030 35872 22094 35876
rect 28736 35932 28800 35936
rect 28736 35876 28740 35932
rect 28740 35876 28796 35932
rect 28796 35876 28800 35932
rect 28736 35872 28800 35876
rect 28816 35932 28880 35936
rect 28816 35876 28820 35932
rect 28820 35876 28876 35932
rect 28876 35876 28880 35932
rect 28816 35872 28880 35876
rect 28896 35932 28960 35936
rect 28896 35876 28900 35932
rect 28900 35876 28956 35932
rect 28956 35876 28960 35932
rect 28896 35872 28960 35876
rect 28976 35932 29040 35936
rect 28976 35876 28980 35932
rect 28980 35876 29036 35932
rect 29036 35876 29040 35932
rect 28976 35872 29040 35876
rect 4425 35388 4489 35392
rect 4425 35332 4429 35388
rect 4429 35332 4485 35388
rect 4485 35332 4489 35388
rect 4425 35328 4489 35332
rect 4505 35388 4569 35392
rect 4505 35332 4509 35388
rect 4509 35332 4565 35388
rect 4565 35332 4569 35388
rect 4505 35328 4569 35332
rect 4585 35388 4649 35392
rect 4585 35332 4589 35388
rect 4589 35332 4645 35388
rect 4645 35332 4649 35388
rect 4585 35328 4649 35332
rect 4665 35388 4729 35392
rect 4665 35332 4669 35388
rect 4669 35332 4725 35388
rect 4725 35332 4729 35388
rect 4665 35328 4729 35332
rect 11371 35388 11435 35392
rect 11371 35332 11375 35388
rect 11375 35332 11431 35388
rect 11431 35332 11435 35388
rect 11371 35328 11435 35332
rect 11451 35388 11515 35392
rect 11451 35332 11455 35388
rect 11455 35332 11511 35388
rect 11511 35332 11515 35388
rect 11451 35328 11515 35332
rect 11531 35388 11595 35392
rect 11531 35332 11535 35388
rect 11535 35332 11591 35388
rect 11591 35332 11595 35388
rect 11531 35328 11595 35332
rect 11611 35388 11675 35392
rect 11611 35332 11615 35388
rect 11615 35332 11671 35388
rect 11671 35332 11675 35388
rect 11611 35328 11675 35332
rect 18317 35388 18381 35392
rect 18317 35332 18321 35388
rect 18321 35332 18377 35388
rect 18377 35332 18381 35388
rect 18317 35328 18381 35332
rect 18397 35388 18461 35392
rect 18397 35332 18401 35388
rect 18401 35332 18457 35388
rect 18457 35332 18461 35388
rect 18397 35328 18461 35332
rect 18477 35388 18541 35392
rect 18477 35332 18481 35388
rect 18481 35332 18537 35388
rect 18537 35332 18541 35388
rect 18477 35328 18541 35332
rect 18557 35388 18621 35392
rect 18557 35332 18561 35388
rect 18561 35332 18617 35388
rect 18617 35332 18621 35388
rect 18557 35328 18621 35332
rect 25263 35388 25327 35392
rect 25263 35332 25267 35388
rect 25267 35332 25323 35388
rect 25323 35332 25327 35388
rect 25263 35328 25327 35332
rect 25343 35388 25407 35392
rect 25343 35332 25347 35388
rect 25347 35332 25403 35388
rect 25403 35332 25407 35388
rect 25343 35328 25407 35332
rect 25423 35388 25487 35392
rect 25423 35332 25427 35388
rect 25427 35332 25483 35388
rect 25483 35332 25487 35388
rect 25423 35328 25487 35332
rect 25503 35388 25567 35392
rect 25503 35332 25507 35388
rect 25507 35332 25563 35388
rect 25563 35332 25567 35388
rect 25503 35328 25567 35332
rect 7898 34844 7962 34848
rect 7898 34788 7902 34844
rect 7902 34788 7958 34844
rect 7958 34788 7962 34844
rect 7898 34784 7962 34788
rect 7978 34844 8042 34848
rect 7978 34788 7982 34844
rect 7982 34788 8038 34844
rect 8038 34788 8042 34844
rect 7978 34784 8042 34788
rect 8058 34844 8122 34848
rect 8058 34788 8062 34844
rect 8062 34788 8118 34844
rect 8118 34788 8122 34844
rect 8058 34784 8122 34788
rect 8138 34844 8202 34848
rect 8138 34788 8142 34844
rect 8142 34788 8198 34844
rect 8198 34788 8202 34844
rect 8138 34784 8202 34788
rect 14844 34844 14908 34848
rect 14844 34788 14848 34844
rect 14848 34788 14904 34844
rect 14904 34788 14908 34844
rect 14844 34784 14908 34788
rect 14924 34844 14988 34848
rect 14924 34788 14928 34844
rect 14928 34788 14984 34844
rect 14984 34788 14988 34844
rect 14924 34784 14988 34788
rect 15004 34844 15068 34848
rect 15004 34788 15008 34844
rect 15008 34788 15064 34844
rect 15064 34788 15068 34844
rect 15004 34784 15068 34788
rect 15084 34844 15148 34848
rect 15084 34788 15088 34844
rect 15088 34788 15144 34844
rect 15144 34788 15148 34844
rect 15084 34784 15148 34788
rect 21790 34844 21854 34848
rect 21790 34788 21794 34844
rect 21794 34788 21850 34844
rect 21850 34788 21854 34844
rect 21790 34784 21854 34788
rect 21870 34844 21934 34848
rect 21870 34788 21874 34844
rect 21874 34788 21930 34844
rect 21930 34788 21934 34844
rect 21870 34784 21934 34788
rect 21950 34844 22014 34848
rect 21950 34788 21954 34844
rect 21954 34788 22010 34844
rect 22010 34788 22014 34844
rect 21950 34784 22014 34788
rect 22030 34844 22094 34848
rect 22030 34788 22034 34844
rect 22034 34788 22090 34844
rect 22090 34788 22094 34844
rect 22030 34784 22094 34788
rect 28736 34844 28800 34848
rect 28736 34788 28740 34844
rect 28740 34788 28796 34844
rect 28796 34788 28800 34844
rect 28736 34784 28800 34788
rect 28816 34844 28880 34848
rect 28816 34788 28820 34844
rect 28820 34788 28876 34844
rect 28876 34788 28880 34844
rect 28816 34784 28880 34788
rect 28896 34844 28960 34848
rect 28896 34788 28900 34844
rect 28900 34788 28956 34844
rect 28956 34788 28960 34844
rect 28896 34784 28960 34788
rect 28976 34844 29040 34848
rect 28976 34788 28980 34844
rect 28980 34788 29036 34844
rect 29036 34788 29040 34844
rect 28976 34784 29040 34788
rect 4425 34300 4489 34304
rect 4425 34244 4429 34300
rect 4429 34244 4485 34300
rect 4485 34244 4489 34300
rect 4425 34240 4489 34244
rect 4505 34300 4569 34304
rect 4505 34244 4509 34300
rect 4509 34244 4565 34300
rect 4565 34244 4569 34300
rect 4505 34240 4569 34244
rect 4585 34300 4649 34304
rect 4585 34244 4589 34300
rect 4589 34244 4645 34300
rect 4645 34244 4649 34300
rect 4585 34240 4649 34244
rect 4665 34300 4729 34304
rect 4665 34244 4669 34300
rect 4669 34244 4725 34300
rect 4725 34244 4729 34300
rect 4665 34240 4729 34244
rect 11371 34300 11435 34304
rect 11371 34244 11375 34300
rect 11375 34244 11431 34300
rect 11431 34244 11435 34300
rect 11371 34240 11435 34244
rect 11451 34300 11515 34304
rect 11451 34244 11455 34300
rect 11455 34244 11511 34300
rect 11511 34244 11515 34300
rect 11451 34240 11515 34244
rect 11531 34300 11595 34304
rect 11531 34244 11535 34300
rect 11535 34244 11591 34300
rect 11591 34244 11595 34300
rect 11531 34240 11595 34244
rect 11611 34300 11675 34304
rect 11611 34244 11615 34300
rect 11615 34244 11671 34300
rect 11671 34244 11675 34300
rect 11611 34240 11675 34244
rect 18317 34300 18381 34304
rect 18317 34244 18321 34300
rect 18321 34244 18377 34300
rect 18377 34244 18381 34300
rect 18317 34240 18381 34244
rect 18397 34300 18461 34304
rect 18397 34244 18401 34300
rect 18401 34244 18457 34300
rect 18457 34244 18461 34300
rect 18397 34240 18461 34244
rect 18477 34300 18541 34304
rect 18477 34244 18481 34300
rect 18481 34244 18537 34300
rect 18537 34244 18541 34300
rect 18477 34240 18541 34244
rect 18557 34300 18621 34304
rect 18557 34244 18561 34300
rect 18561 34244 18617 34300
rect 18617 34244 18621 34300
rect 18557 34240 18621 34244
rect 25263 34300 25327 34304
rect 25263 34244 25267 34300
rect 25267 34244 25323 34300
rect 25323 34244 25327 34300
rect 25263 34240 25327 34244
rect 25343 34300 25407 34304
rect 25343 34244 25347 34300
rect 25347 34244 25403 34300
rect 25403 34244 25407 34300
rect 25343 34240 25407 34244
rect 25423 34300 25487 34304
rect 25423 34244 25427 34300
rect 25427 34244 25483 34300
rect 25483 34244 25487 34300
rect 25423 34240 25487 34244
rect 25503 34300 25567 34304
rect 25503 34244 25507 34300
rect 25507 34244 25563 34300
rect 25563 34244 25567 34300
rect 25503 34240 25567 34244
rect 7898 33756 7962 33760
rect 7898 33700 7902 33756
rect 7902 33700 7958 33756
rect 7958 33700 7962 33756
rect 7898 33696 7962 33700
rect 7978 33756 8042 33760
rect 7978 33700 7982 33756
rect 7982 33700 8038 33756
rect 8038 33700 8042 33756
rect 7978 33696 8042 33700
rect 8058 33756 8122 33760
rect 8058 33700 8062 33756
rect 8062 33700 8118 33756
rect 8118 33700 8122 33756
rect 8058 33696 8122 33700
rect 8138 33756 8202 33760
rect 8138 33700 8142 33756
rect 8142 33700 8198 33756
rect 8198 33700 8202 33756
rect 8138 33696 8202 33700
rect 14844 33756 14908 33760
rect 14844 33700 14848 33756
rect 14848 33700 14904 33756
rect 14904 33700 14908 33756
rect 14844 33696 14908 33700
rect 14924 33756 14988 33760
rect 14924 33700 14928 33756
rect 14928 33700 14984 33756
rect 14984 33700 14988 33756
rect 14924 33696 14988 33700
rect 15004 33756 15068 33760
rect 15004 33700 15008 33756
rect 15008 33700 15064 33756
rect 15064 33700 15068 33756
rect 15004 33696 15068 33700
rect 15084 33756 15148 33760
rect 15084 33700 15088 33756
rect 15088 33700 15144 33756
rect 15144 33700 15148 33756
rect 15084 33696 15148 33700
rect 21790 33756 21854 33760
rect 21790 33700 21794 33756
rect 21794 33700 21850 33756
rect 21850 33700 21854 33756
rect 21790 33696 21854 33700
rect 21870 33756 21934 33760
rect 21870 33700 21874 33756
rect 21874 33700 21930 33756
rect 21930 33700 21934 33756
rect 21870 33696 21934 33700
rect 21950 33756 22014 33760
rect 21950 33700 21954 33756
rect 21954 33700 22010 33756
rect 22010 33700 22014 33756
rect 21950 33696 22014 33700
rect 22030 33756 22094 33760
rect 22030 33700 22034 33756
rect 22034 33700 22090 33756
rect 22090 33700 22094 33756
rect 22030 33696 22094 33700
rect 28736 33756 28800 33760
rect 28736 33700 28740 33756
rect 28740 33700 28796 33756
rect 28796 33700 28800 33756
rect 28736 33696 28800 33700
rect 28816 33756 28880 33760
rect 28816 33700 28820 33756
rect 28820 33700 28876 33756
rect 28876 33700 28880 33756
rect 28816 33696 28880 33700
rect 28896 33756 28960 33760
rect 28896 33700 28900 33756
rect 28900 33700 28956 33756
rect 28956 33700 28960 33756
rect 28896 33696 28960 33700
rect 28976 33756 29040 33760
rect 28976 33700 28980 33756
rect 28980 33700 29036 33756
rect 29036 33700 29040 33756
rect 28976 33696 29040 33700
rect 4425 33212 4489 33216
rect 4425 33156 4429 33212
rect 4429 33156 4485 33212
rect 4485 33156 4489 33212
rect 4425 33152 4489 33156
rect 4505 33212 4569 33216
rect 4505 33156 4509 33212
rect 4509 33156 4565 33212
rect 4565 33156 4569 33212
rect 4505 33152 4569 33156
rect 4585 33212 4649 33216
rect 4585 33156 4589 33212
rect 4589 33156 4645 33212
rect 4645 33156 4649 33212
rect 4585 33152 4649 33156
rect 4665 33212 4729 33216
rect 4665 33156 4669 33212
rect 4669 33156 4725 33212
rect 4725 33156 4729 33212
rect 4665 33152 4729 33156
rect 11371 33212 11435 33216
rect 11371 33156 11375 33212
rect 11375 33156 11431 33212
rect 11431 33156 11435 33212
rect 11371 33152 11435 33156
rect 11451 33212 11515 33216
rect 11451 33156 11455 33212
rect 11455 33156 11511 33212
rect 11511 33156 11515 33212
rect 11451 33152 11515 33156
rect 11531 33212 11595 33216
rect 11531 33156 11535 33212
rect 11535 33156 11591 33212
rect 11591 33156 11595 33212
rect 11531 33152 11595 33156
rect 11611 33212 11675 33216
rect 11611 33156 11615 33212
rect 11615 33156 11671 33212
rect 11671 33156 11675 33212
rect 11611 33152 11675 33156
rect 18317 33212 18381 33216
rect 18317 33156 18321 33212
rect 18321 33156 18377 33212
rect 18377 33156 18381 33212
rect 18317 33152 18381 33156
rect 18397 33212 18461 33216
rect 18397 33156 18401 33212
rect 18401 33156 18457 33212
rect 18457 33156 18461 33212
rect 18397 33152 18461 33156
rect 18477 33212 18541 33216
rect 18477 33156 18481 33212
rect 18481 33156 18537 33212
rect 18537 33156 18541 33212
rect 18477 33152 18541 33156
rect 18557 33212 18621 33216
rect 18557 33156 18561 33212
rect 18561 33156 18617 33212
rect 18617 33156 18621 33212
rect 18557 33152 18621 33156
rect 25263 33212 25327 33216
rect 25263 33156 25267 33212
rect 25267 33156 25323 33212
rect 25323 33156 25327 33212
rect 25263 33152 25327 33156
rect 25343 33212 25407 33216
rect 25343 33156 25347 33212
rect 25347 33156 25403 33212
rect 25403 33156 25407 33212
rect 25343 33152 25407 33156
rect 25423 33212 25487 33216
rect 25423 33156 25427 33212
rect 25427 33156 25483 33212
rect 25483 33156 25487 33212
rect 25423 33152 25487 33156
rect 25503 33212 25567 33216
rect 25503 33156 25507 33212
rect 25507 33156 25563 33212
rect 25563 33156 25567 33212
rect 25503 33152 25567 33156
rect 7898 32668 7962 32672
rect 7898 32612 7902 32668
rect 7902 32612 7958 32668
rect 7958 32612 7962 32668
rect 7898 32608 7962 32612
rect 7978 32668 8042 32672
rect 7978 32612 7982 32668
rect 7982 32612 8038 32668
rect 8038 32612 8042 32668
rect 7978 32608 8042 32612
rect 8058 32668 8122 32672
rect 8058 32612 8062 32668
rect 8062 32612 8118 32668
rect 8118 32612 8122 32668
rect 8058 32608 8122 32612
rect 8138 32668 8202 32672
rect 8138 32612 8142 32668
rect 8142 32612 8198 32668
rect 8198 32612 8202 32668
rect 8138 32608 8202 32612
rect 14844 32668 14908 32672
rect 14844 32612 14848 32668
rect 14848 32612 14904 32668
rect 14904 32612 14908 32668
rect 14844 32608 14908 32612
rect 14924 32668 14988 32672
rect 14924 32612 14928 32668
rect 14928 32612 14984 32668
rect 14984 32612 14988 32668
rect 14924 32608 14988 32612
rect 15004 32668 15068 32672
rect 15004 32612 15008 32668
rect 15008 32612 15064 32668
rect 15064 32612 15068 32668
rect 15004 32608 15068 32612
rect 15084 32668 15148 32672
rect 15084 32612 15088 32668
rect 15088 32612 15144 32668
rect 15144 32612 15148 32668
rect 15084 32608 15148 32612
rect 21790 32668 21854 32672
rect 21790 32612 21794 32668
rect 21794 32612 21850 32668
rect 21850 32612 21854 32668
rect 21790 32608 21854 32612
rect 21870 32668 21934 32672
rect 21870 32612 21874 32668
rect 21874 32612 21930 32668
rect 21930 32612 21934 32668
rect 21870 32608 21934 32612
rect 21950 32668 22014 32672
rect 21950 32612 21954 32668
rect 21954 32612 22010 32668
rect 22010 32612 22014 32668
rect 21950 32608 22014 32612
rect 22030 32668 22094 32672
rect 22030 32612 22034 32668
rect 22034 32612 22090 32668
rect 22090 32612 22094 32668
rect 22030 32608 22094 32612
rect 28736 32668 28800 32672
rect 28736 32612 28740 32668
rect 28740 32612 28796 32668
rect 28796 32612 28800 32668
rect 28736 32608 28800 32612
rect 28816 32668 28880 32672
rect 28816 32612 28820 32668
rect 28820 32612 28876 32668
rect 28876 32612 28880 32668
rect 28816 32608 28880 32612
rect 28896 32668 28960 32672
rect 28896 32612 28900 32668
rect 28900 32612 28956 32668
rect 28956 32612 28960 32668
rect 28896 32608 28960 32612
rect 28976 32668 29040 32672
rect 28976 32612 28980 32668
rect 28980 32612 29036 32668
rect 29036 32612 29040 32668
rect 28976 32608 29040 32612
rect 4425 32124 4489 32128
rect 4425 32068 4429 32124
rect 4429 32068 4485 32124
rect 4485 32068 4489 32124
rect 4425 32064 4489 32068
rect 4505 32124 4569 32128
rect 4505 32068 4509 32124
rect 4509 32068 4565 32124
rect 4565 32068 4569 32124
rect 4505 32064 4569 32068
rect 4585 32124 4649 32128
rect 4585 32068 4589 32124
rect 4589 32068 4645 32124
rect 4645 32068 4649 32124
rect 4585 32064 4649 32068
rect 4665 32124 4729 32128
rect 4665 32068 4669 32124
rect 4669 32068 4725 32124
rect 4725 32068 4729 32124
rect 4665 32064 4729 32068
rect 11371 32124 11435 32128
rect 11371 32068 11375 32124
rect 11375 32068 11431 32124
rect 11431 32068 11435 32124
rect 11371 32064 11435 32068
rect 11451 32124 11515 32128
rect 11451 32068 11455 32124
rect 11455 32068 11511 32124
rect 11511 32068 11515 32124
rect 11451 32064 11515 32068
rect 11531 32124 11595 32128
rect 11531 32068 11535 32124
rect 11535 32068 11591 32124
rect 11591 32068 11595 32124
rect 11531 32064 11595 32068
rect 11611 32124 11675 32128
rect 11611 32068 11615 32124
rect 11615 32068 11671 32124
rect 11671 32068 11675 32124
rect 11611 32064 11675 32068
rect 18317 32124 18381 32128
rect 18317 32068 18321 32124
rect 18321 32068 18377 32124
rect 18377 32068 18381 32124
rect 18317 32064 18381 32068
rect 18397 32124 18461 32128
rect 18397 32068 18401 32124
rect 18401 32068 18457 32124
rect 18457 32068 18461 32124
rect 18397 32064 18461 32068
rect 18477 32124 18541 32128
rect 18477 32068 18481 32124
rect 18481 32068 18537 32124
rect 18537 32068 18541 32124
rect 18477 32064 18541 32068
rect 18557 32124 18621 32128
rect 18557 32068 18561 32124
rect 18561 32068 18617 32124
rect 18617 32068 18621 32124
rect 18557 32064 18621 32068
rect 25263 32124 25327 32128
rect 25263 32068 25267 32124
rect 25267 32068 25323 32124
rect 25323 32068 25327 32124
rect 25263 32064 25327 32068
rect 25343 32124 25407 32128
rect 25343 32068 25347 32124
rect 25347 32068 25403 32124
rect 25403 32068 25407 32124
rect 25343 32064 25407 32068
rect 25423 32124 25487 32128
rect 25423 32068 25427 32124
rect 25427 32068 25483 32124
rect 25483 32068 25487 32124
rect 25423 32064 25487 32068
rect 25503 32124 25567 32128
rect 25503 32068 25507 32124
rect 25507 32068 25563 32124
rect 25563 32068 25567 32124
rect 25503 32064 25567 32068
rect 7898 31580 7962 31584
rect 7898 31524 7902 31580
rect 7902 31524 7958 31580
rect 7958 31524 7962 31580
rect 7898 31520 7962 31524
rect 7978 31580 8042 31584
rect 7978 31524 7982 31580
rect 7982 31524 8038 31580
rect 8038 31524 8042 31580
rect 7978 31520 8042 31524
rect 8058 31580 8122 31584
rect 8058 31524 8062 31580
rect 8062 31524 8118 31580
rect 8118 31524 8122 31580
rect 8058 31520 8122 31524
rect 8138 31580 8202 31584
rect 8138 31524 8142 31580
rect 8142 31524 8198 31580
rect 8198 31524 8202 31580
rect 8138 31520 8202 31524
rect 14844 31580 14908 31584
rect 14844 31524 14848 31580
rect 14848 31524 14904 31580
rect 14904 31524 14908 31580
rect 14844 31520 14908 31524
rect 14924 31580 14988 31584
rect 14924 31524 14928 31580
rect 14928 31524 14984 31580
rect 14984 31524 14988 31580
rect 14924 31520 14988 31524
rect 15004 31580 15068 31584
rect 15004 31524 15008 31580
rect 15008 31524 15064 31580
rect 15064 31524 15068 31580
rect 15004 31520 15068 31524
rect 15084 31580 15148 31584
rect 15084 31524 15088 31580
rect 15088 31524 15144 31580
rect 15144 31524 15148 31580
rect 15084 31520 15148 31524
rect 21790 31580 21854 31584
rect 21790 31524 21794 31580
rect 21794 31524 21850 31580
rect 21850 31524 21854 31580
rect 21790 31520 21854 31524
rect 21870 31580 21934 31584
rect 21870 31524 21874 31580
rect 21874 31524 21930 31580
rect 21930 31524 21934 31580
rect 21870 31520 21934 31524
rect 21950 31580 22014 31584
rect 21950 31524 21954 31580
rect 21954 31524 22010 31580
rect 22010 31524 22014 31580
rect 21950 31520 22014 31524
rect 22030 31580 22094 31584
rect 22030 31524 22034 31580
rect 22034 31524 22090 31580
rect 22090 31524 22094 31580
rect 22030 31520 22094 31524
rect 28736 31580 28800 31584
rect 28736 31524 28740 31580
rect 28740 31524 28796 31580
rect 28796 31524 28800 31580
rect 28736 31520 28800 31524
rect 28816 31580 28880 31584
rect 28816 31524 28820 31580
rect 28820 31524 28876 31580
rect 28876 31524 28880 31580
rect 28816 31520 28880 31524
rect 28896 31580 28960 31584
rect 28896 31524 28900 31580
rect 28900 31524 28956 31580
rect 28956 31524 28960 31580
rect 28896 31520 28960 31524
rect 28976 31580 29040 31584
rect 28976 31524 28980 31580
rect 28980 31524 29036 31580
rect 29036 31524 29040 31580
rect 28976 31520 29040 31524
rect 4425 31036 4489 31040
rect 4425 30980 4429 31036
rect 4429 30980 4485 31036
rect 4485 30980 4489 31036
rect 4425 30976 4489 30980
rect 4505 31036 4569 31040
rect 4505 30980 4509 31036
rect 4509 30980 4565 31036
rect 4565 30980 4569 31036
rect 4505 30976 4569 30980
rect 4585 31036 4649 31040
rect 4585 30980 4589 31036
rect 4589 30980 4645 31036
rect 4645 30980 4649 31036
rect 4585 30976 4649 30980
rect 4665 31036 4729 31040
rect 4665 30980 4669 31036
rect 4669 30980 4725 31036
rect 4725 30980 4729 31036
rect 4665 30976 4729 30980
rect 11371 31036 11435 31040
rect 11371 30980 11375 31036
rect 11375 30980 11431 31036
rect 11431 30980 11435 31036
rect 11371 30976 11435 30980
rect 11451 31036 11515 31040
rect 11451 30980 11455 31036
rect 11455 30980 11511 31036
rect 11511 30980 11515 31036
rect 11451 30976 11515 30980
rect 11531 31036 11595 31040
rect 11531 30980 11535 31036
rect 11535 30980 11591 31036
rect 11591 30980 11595 31036
rect 11531 30976 11595 30980
rect 11611 31036 11675 31040
rect 11611 30980 11615 31036
rect 11615 30980 11671 31036
rect 11671 30980 11675 31036
rect 11611 30976 11675 30980
rect 18317 31036 18381 31040
rect 18317 30980 18321 31036
rect 18321 30980 18377 31036
rect 18377 30980 18381 31036
rect 18317 30976 18381 30980
rect 18397 31036 18461 31040
rect 18397 30980 18401 31036
rect 18401 30980 18457 31036
rect 18457 30980 18461 31036
rect 18397 30976 18461 30980
rect 18477 31036 18541 31040
rect 18477 30980 18481 31036
rect 18481 30980 18537 31036
rect 18537 30980 18541 31036
rect 18477 30976 18541 30980
rect 18557 31036 18621 31040
rect 18557 30980 18561 31036
rect 18561 30980 18617 31036
rect 18617 30980 18621 31036
rect 18557 30976 18621 30980
rect 25263 31036 25327 31040
rect 25263 30980 25267 31036
rect 25267 30980 25323 31036
rect 25323 30980 25327 31036
rect 25263 30976 25327 30980
rect 25343 31036 25407 31040
rect 25343 30980 25347 31036
rect 25347 30980 25403 31036
rect 25403 30980 25407 31036
rect 25343 30976 25407 30980
rect 25423 31036 25487 31040
rect 25423 30980 25427 31036
rect 25427 30980 25483 31036
rect 25483 30980 25487 31036
rect 25423 30976 25487 30980
rect 25503 31036 25567 31040
rect 25503 30980 25507 31036
rect 25507 30980 25563 31036
rect 25563 30980 25567 31036
rect 25503 30976 25567 30980
rect 7898 30492 7962 30496
rect 7898 30436 7902 30492
rect 7902 30436 7958 30492
rect 7958 30436 7962 30492
rect 7898 30432 7962 30436
rect 7978 30492 8042 30496
rect 7978 30436 7982 30492
rect 7982 30436 8038 30492
rect 8038 30436 8042 30492
rect 7978 30432 8042 30436
rect 8058 30492 8122 30496
rect 8058 30436 8062 30492
rect 8062 30436 8118 30492
rect 8118 30436 8122 30492
rect 8058 30432 8122 30436
rect 8138 30492 8202 30496
rect 8138 30436 8142 30492
rect 8142 30436 8198 30492
rect 8198 30436 8202 30492
rect 8138 30432 8202 30436
rect 14844 30492 14908 30496
rect 14844 30436 14848 30492
rect 14848 30436 14904 30492
rect 14904 30436 14908 30492
rect 14844 30432 14908 30436
rect 14924 30492 14988 30496
rect 14924 30436 14928 30492
rect 14928 30436 14984 30492
rect 14984 30436 14988 30492
rect 14924 30432 14988 30436
rect 15004 30492 15068 30496
rect 15004 30436 15008 30492
rect 15008 30436 15064 30492
rect 15064 30436 15068 30492
rect 15004 30432 15068 30436
rect 15084 30492 15148 30496
rect 15084 30436 15088 30492
rect 15088 30436 15144 30492
rect 15144 30436 15148 30492
rect 15084 30432 15148 30436
rect 21790 30492 21854 30496
rect 21790 30436 21794 30492
rect 21794 30436 21850 30492
rect 21850 30436 21854 30492
rect 21790 30432 21854 30436
rect 21870 30492 21934 30496
rect 21870 30436 21874 30492
rect 21874 30436 21930 30492
rect 21930 30436 21934 30492
rect 21870 30432 21934 30436
rect 21950 30492 22014 30496
rect 21950 30436 21954 30492
rect 21954 30436 22010 30492
rect 22010 30436 22014 30492
rect 21950 30432 22014 30436
rect 22030 30492 22094 30496
rect 22030 30436 22034 30492
rect 22034 30436 22090 30492
rect 22090 30436 22094 30492
rect 22030 30432 22094 30436
rect 28736 30492 28800 30496
rect 28736 30436 28740 30492
rect 28740 30436 28796 30492
rect 28796 30436 28800 30492
rect 28736 30432 28800 30436
rect 28816 30492 28880 30496
rect 28816 30436 28820 30492
rect 28820 30436 28876 30492
rect 28876 30436 28880 30492
rect 28816 30432 28880 30436
rect 28896 30492 28960 30496
rect 28896 30436 28900 30492
rect 28900 30436 28956 30492
rect 28956 30436 28960 30492
rect 28896 30432 28960 30436
rect 28976 30492 29040 30496
rect 28976 30436 28980 30492
rect 28980 30436 29036 30492
rect 29036 30436 29040 30492
rect 28976 30432 29040 30436
rect 4425 29948 4489 29952
rect 4425 29892 4429 29948
rect 4429 29892 4485 29948
rect 4485 29892 4489 29948
rect 4425 29888 4489 29892
rect 4505 29948 4569 29952
rect 4505 29892 4509 29948
rect 4509 29892 4565 29948
rect 4565 29892 4569 29948
rect 4505 29888 4569 29892
rect 4585 29948 4649 29952
rect 4585 29892 4589 29948
rect 4589 29892 4645 29948
rect 4645 29892 4649 29948
rect 4585 29888 4649 29892
rect 4665 29948 4729 29952
rect 4665 29892 4669 29948
rect 4669 29892 4725 29948
rect 4725 29892 4729 29948
rect 4665 29888 4729 29892
rect 11371 29948 11435 29952
rect 11371 29892 11375 29948
rect 11375 29892 11431 29948
rect 11431 29892 11435 29948
rect 11371 29888 11435 29892
rect 11451 29948 11515 29952
rect 11451 29892 11455 29948
rect 11455 29892 11511 29948
rect 11511 29892 11515 29948
rect 11451 29888 11515 29892
rect 11531 29948 11595 29952
rect 11531 29892 11535 29948
rect 11535 29892 11591 29948
rect 11591 29892 11595 29948
rect 11531 29888 11595 29892
rect 11611 29948 11675 29952
rect 11611 29892 11615 29948
rect 11615 29892 11671 29948
rect 11671 29892 11675 29948
rect 11611 29888 11675 29892
rect 18317 29948 18381 29952
rect 18317 29892 18321 29948
rect 18321 29892 18377 29948
rect 18377 29892 18381 29948
rect 18317 29888 18381 29892
rect 18397 29948 18461 29952
rect 18397 29892 18401 29948
rect 18401 29892 18457 29948
rect 18457 29892 18461 29948
rect 18397 29888 18461 29892
rect 18477 29948 18541 29952
rect 18477 29892 18481 29948
rect 18481 29892 18537 29948
rect 18537 29892 18541 29948
rect 18477 29888 18541 29892
rect 18557 29948 18621 29952
rect 18557 29892 18561 29948
rect 18561 29892 18617 29948
rect 18617 29892 18621 29948
rect 18557 29888 18621 29892
rect 25263 29948 25327 29952
rect 25263 29892 25267 29948
rect 25267 29892 25323 29948
rect 25323 29892 25327 29948
rect 25263 29888 25327 29892
rect 25343 29948 25407 29952
rect 25343 29892 25347 29948
rect 25347 29892 25403 29948
rect 25403 29892 25407 29948
rect 25343 29888 25407 29892
rect 25423 29948 25487 29952
rect 25423 29892 25427 29948
rect 25427 29892 25483 29948
rect 25483 29892 25487 29948
rect 25423 29888 25487 29892
rect 25503 29948 25567 29952
rect 25503 29892 25507 29948
rect 25507 29892 25563 29948
rect 25563 29892 25567 29948
rect 25503 29888 25567 29892
rect 7898 29404 7962 29408
rect 7898 29348 7902 29404
rect 7902 29348 7958 29404
rect 7958 29348 7962 29404
rect 7898 29344 7962 29348
rect 7978 29404 8042 29408
rect 7978 29348 7982 29404
rect 7982 29348 8038 29404
rect 8038 29348 8042 29404
rect 7978 29344 8042 29348
rect 8058 29404 8122 29408
rect 8058 29348 8062 29404
rect 8062 29348 8118 29404
rect 8118 29348 8122 29404
rect 8058 29344 8122 29348
rect 8138 29404 8202 29408
rect 8138 29348 8142 29404
rect 8142 29348 8198 29404
rect 8198 29348 8202 29404
rect 8138 29344 8202 29348
rect 14844 29404 14908 29408
rect 14844 29348 14848 29404
rect 14848 29348 14904 29404
rect 14904 29348 14908 29404
rect 14844 29344 14908 29348
rect 14924 29404 14988 29408
rect 14924 29348 14928 29404
rect 14928 29348 14984 29404
rect 14984 29348 14988 29404
rect 14924 29344 14988 29348
rect 15004 29404 15068 29408
rect 15004 29348 15008 29404
rect 15008 29348 15064 29404
rect 15064 29348 15068 29404
rect 15004 29344 15068 29348
rect 15084 29404 15148 29408
rect 15084 29348 15088 29404
rect 15088 29348 15144 29404
rect 15144 29348 15148 29404
rect 15084 29344 15148 29348
rect 21790 29404 21854 29408
rect 21790 29348 21794 29404
rect 21794 29348 21850 29404
rect 21850 29348 21854 29404
rect 21790 29344 21854 29348
rect 21870 29404 21934 29408
rect 21870 29348 21874 29404
rect 21874 29348 21930 29404
rect 21930 29348 21934 29404
rect 21870 29344 21934 29348
rect 21950 29404 22014 29408
rect 21950 29348 21954 29404
rect 21954 29348 22010 29404
rect 22010 29348 22014 29404
rect 21950 29344 22014 29348
rect 22030 29404 22094 29408
rect 22030 29348 22034 29404
rect 22034 29348 22090 29404
rect 22090 29348 22094 29404
rect 22030 29344 22094 29348
rect 28736 29404 28800 29408
rect 28736 29348 28740 29404
rect 28740 29348 28796 29404
rect 28796 29348 28800 29404
rect 28736 29344 28800 29348
rect 28816 29404 28880 29408
rect 28816 29348 28820 29404
rect 28820 29348 28876 29404
rect 28876 29348 28880 29404
rect 28816 29344 28880 29348
rect 28896 29404 28960 29408
rect 28896 29348 28900 29404
rect 28900 29348 28956 29404
rect 28956 29348 28960 29404
rect 28896 29344 28960 29348
rect 28976 29404 29040 29408
rect 28976 29348 28980 29404
rect 28980 29348 29036 29404
rect 29036 29348 29040 29404
rect 28976 29344 29040 29348
rect 4425 28860 4489 28864
rect 4425 28804 4429 28860
rect 4429 28804 4485 28860
rect 4485 28804 4489 28860
rect 4425 28800 4489 28804
rect 4505 28860 4569 28864
rect 4505 28804 4509 28860
rect 4509 28804 4565 28860
rect 4565 28804 4569 28860
rect 4505 28800 4569 28804
rect 4585 28860 4649 28864
rect 4585 28804 4589 28860
rect 4589 28804 4645 28860
rect 4645 28804 4649 28860
rect 4585 28800 4649 28804
rect 4665 28860 4729 28864
rect 4665 28804 4669 28860
rect 4669 28804 4725 28860
rect 4725 28804 4729 28860
rect 4665 28800 4729 28804
rect 11371 28860 11435 28864
rect 11371 28804 11375 28860
rect 11375 28804 11431 28860
rect 11431 28804 11435 28860
rect 11371 28800 11435 28804
rect 11451 28860 11515 28864
rect 11451 28804 11455 28860
rect 11455 28804 11511 28860
rect 11511 28804 11515 28860
rect 11451 28800 11515 28804
rect 11531 28860 11595 28864
rect 11531 28804 11535 28860
rect 11535 28804 11591 28860
rect 11591 28804 11595 28860
rect 11531 28800 11595 28804
rect 11611 28860 11675 28864
rect 11611 28804 11615 28860
rect 11615 28804 11671 28860
rect 11671 28804 11675 28860
rect 11611 28800 11675 28804
rect 18317 28860 18381 28864
rect 18317 28804 18321 28860
rect 18321 28804 18377 28860
rect 18377 28804 18381 28860
rect 18317 28800 18381 28804
rect 18397 28860 18461 28864
rect 18397 28804 18401 28860
rect 18401 28804 18457 28860
rect 18457 28804 18461 28860
rect 18397 28800 18461 28804
rect 18477 28860 18541 28864
rect 18477 28804 18481 28860
rect 18481 28804 18537 28860
rect 18537 28804 18541 28860
rect 18477 28800 18541 28804
rect 18557 28860 18621 28864
rect 18557 28804 18561 28860
rect 18561 28804 18617 28860
rect 18617 28804 18621 28860
rect 18557 28800 18621 28804
rect 25263 28860 25327 28864
rect 25263 28804 25267 28860
rect 25267 28804 25323 28860
rect 25323 28804 25327 28860
rect 25263 28800 25327 28804
rect 25343 28860 25407 28864
rect 25343 28804 25347 28860
rect 25347 28804 25403 28860
rect 25403 28804 25407 28860
rect 25343 28800 25407 28804
rect 25423 28860 25487 28864
rect 25423 28804 25427 28860
rect 25427 28804 25483 28860
rect 25483 28804 25487 28860
rect 25423 28800 25487 28804
rect 25503 28860 25567 28864
rect 25503 28804 25507 28860
rect 25507 28804 25563 28860
rect 25563 28804 25567 28860
rect 25503 28800 25567 28804
rect 7898 28316 7962 28320
rect 7898 28260 7902 28316
rect 7902 28260 7958 28316
rect 7958 28260 7962 28316
rect 7898 28256 7962 28260
rect 7978 28316 8042 28320
rect 7978 28260 7982 28316
rect 7982 28260 8038 28316
rect 8038 28260 8042 28316
rect 7978 28256 8042 28260
rect 8058 28316 8122 28320
rect 8058 28260 8062 28316
rect 8062 28260 8118 28316
rect 8118 28260 8122 28316
rect 8058 28256 8122 28260
rect 8138 28316 8202 28320
rect 8138 28260 8142 28316
rect 8142 28260 8198 28316
rect 8198 28260 8202 28316
rect 8138 28256 8202 28260
rect 14844 28316 14908 28320
rect 14844 28260 14848 28316
rect 14848 28260 14904 28316
rect 14904 28260 14908 28316
rect 14844 28256 14908 28260
rect 14924 28316 14988 28320
rect 14924 28260 14928 28316
rect 14928 28260 14984 28316
rect 14984 28260 14988 28316
rect 14924 28256 14988 28260
rect 15004 28316 15068 28320
rect 15004 28260 15008 28316
rect 15008 28260 15064 28316
rect 15064 28260 15068 28316
rect 15004 28256 15068 28260
rect 15084 28316 15148 28320
rect 15084 28260 15088 28316
rect 15088 28260 15144 28316
rect 15144 28260 15148 28316
rect 15084 28256 15148 28260
rect 21790 28316 21854 28320
rect 21790 28260 21794 28316
rect 21794 28260 21850 28316
rect 21850 28260 21854 28316
rect 21790 28256 21854 28260
rect 21870 28316 21934 28320
rect 21870 28260 21874 28316
rect 21874 28260 21930 28316
rect 21930 28260 21934 28316
rect 21870 28256 21934 28260
rect 21950 28316 22014 28320
rect 21950 28260 21954 28316
rect 21954 28260 22010 28316
rect 22010 28260 22014 28316
rect 21950 28256 22014 28260
rect 22030 28316 22094 28320
rect 22030 28260 22034 28316
rect 22034 28260 22090 28316
rect 22090 28260 22094 28316
rect 22030 28256 22094 28260
rect 28736 28316 28800 28320
rect 28736 28260 28740 28316
rect 28740 28260 28796 28316
rect 28796 28260 28800 28316
rect 28736 28256 28800 28260
rect 28816 28316 28880 28320
rect 28816 28260 28820 28316
rect 28820 28260 28876 28316
rect 28876 28260 28880 28316
rect 28816 28256 28880 28260
rect 28896 28316 28960 28320
rect 28896 28260 28900 28316
rect 28900 28260 28956 28316
rect 28956 28260 28960 28316
rect 28896 28256 28960 28260
rect 28976 28316 29040 28320
rect 28976 28260 28980 28316
rect 28980 28260 29036 28316
rect 29036 28260 29040 28316
rect 28976 28256 29040 28260
rect 18828 27976 18892 27980
rect 18828 27920 18878 27976
rect 18878 27920 18892 27976
rect 18828 27916 18892 27920
rect 4425 27772 4489 27776
rect 4425 27716 4429 27772
rect 4429 27716 4485 27772
rect 4485 27716 4489 27772
rect 4425 27712 4489 27716
rect 4505 27772 4569 27776
rect 4505 27716 4509 27772
rect 4509 27716 4565 27772
rect 4565 27716 4569 27772
rect 4505 27712 4569 27716
rect 4585 27772 4649 27776
rect 4585 27716 4589 27772
rect 4589 27716 4645 27772
rect 4645 27716 4649 27772
rect 4585 27712 4649 27716
rect 4665 27772 4729 27776
rect 4665 27716 4669 27772
rect 4669 27716 4725 27772
rect 4725 27716 4729 27772
rect 4665 27712 4729 27716
rect 11371 27772 11435 27776
rect 11371 27716 11375 27772
rect 11375 27716 11431 27772
rect 11431 27716 11435 27772
rect 11371 27712 11435 27716
rect 11451 27772 11515 27776
rect 11451 27716 11455 27772
rect 11455 27716 11511 27772
rect 11511 27716 11515 27772
rect 11451 27712 11515 27716
rect 11531 27772 11595 27776
rect 11531 27716 11535 27772
rect 11535 27716 11591 27772
rect 11591 27716 11595 27772
rect 11531 27712 11595 27716
rect 11611 27772 11675 27776
rect 11611 27716 11615 27772
rect 11615 27716 11671 27772
rect 11671 27716 11675 27772
rect 11611 27712 11675 27716
rect 18317 27772 18381 27776
rect 18317 27716 18321 27772
rect 18321 27716 18377 27772
rect 18377 27716 18381 27772
rect 18317 27712 18381 27716
rect 18397 27772 18461 27776
rect 18397 27716 18401 27772
rect 18401 27716 18457 27772
rect 18457 27716 18461 27772
rect 18397 27712 18461 27716
rect 18477 27772 18541 27776
rect 18477 27716 18481 27772
rect 18481 27716 18537 27772
rect 18537 27716 18541 27772
rect 18477 27712 18541 27716
rect 18557 27772 18621 27776
rect 18557 27716 18561 27772
rect 18561 27716 18617 27772
rect 18617 27716 18621 27772
rect 18557 27712 18621 27716
rect 25263 27772 25327 27776
rect 25263 27716 25267 27772
rect 25267 27716 25323 27772
rect 25323 27716 25327 27772
rect 25263 27712 25327 27716
rect 25343 27772 25407 27776
rect 25343 27716 25347 27772
rect 25347 27716 25403 27772
rect 25403 27716 25407 27772
rect 25343 27712 25407 27716
rect 25423 27772 25487 27776
rect 25423 27716 25427 27772
rect 25427 27716 25483 27772
rect 25483 27716 25487 27772
rect 25423 27712 25487 27716
rect 25503 27772 25567 27776
rect 25503 27716 25507 27772
rect 25507 27716 25563 27772
rect 25563 27716 25567 27772
rect 25503 27712 25567 27716
rect 7898 27228 7962 27232
rect 7898 27172 7902 27228
rect 7902 27172 7958 27228
rect 7958 27172 7962 27228
rect 7898 27168 7962 27172
rect 7978 27228 8042 27232
rect 7978 27172 7982 27228
rect 7982 27172 8038 27228
rect 8038 27172 8042 27228
rect 7978 27168 8042 27172
rect 8058 27228 8122 27232
rect 8058 27172 8062 27228
rect 8062 27172 8118 27228
rect 8118 27172 8122 27228
rect 8058 27168 8122 27172
rect 8138 27228 8202 27232
rect 8138 27172 8142 27228
rect 8142 27172 8198 27228
rect 8198 27172 8202 27228
rect 8138 27168 8202 27172
rect 14844 27228 14908 27232
rect 14844 27172 14848 27228
rect 14848 27172 14904 27228
rect 14904 27172 14908 27228
rect 14844 27168 14908 27172
rect 14924 27228 14988 27232
rect 14924 27172 14928 27228
rect 14928 27172 14984 27228
rect 14984 27172 14988 27228
rect 14924 27168 14988 27172
rect 15004 27228 15068 27232
rect 15004 27172 15008 27228
rect 15008 27172 15064 27228
rect 15064 27172 15068 27228
rect 15004 27168 15068 27172
rect 15084 27228 15148 27232
rect 15084 27172 15088 27228
rect 15088 27172 15144 27228
rect 15144 27172 15148 27228
rect 15084 27168 15148 27172
rect 21790 27228 21854 27232
rect 21790 27172 21794 27228
rect 21794 27172 21850 27228
rect 21850 27172 21854 27228
rect 21790 27168 21854 27172
rect 21870 27228 21934 27232
rect 21870 27172 21874 27228
rect 21874 27172 21930 27228
rect 21930 27172 21934 27228
rect 21870 27168 21934 27172
rect 21950 27228 22014 27232
rect 21950 27172 21954 27228
rect 21954 27172 22010 27228
rect 22010 27172 22014 27228
rect 21950 27168 22014 27172
rect 22030 27228 22094 27232
rect 22030 27172 22034 27228
rect 22034 27172 22090 27228
rect 22090 27172 22094 27228
rect 22030 27168 22094 27172
rect 28736 27228 28800 27232
rect 28736 27172 28740 27228
rect 28740 27172 28796 27228
rect 28796 27172 28800 27228
rect 28736 27168 28800 27172
rect 28816 27228 28880 27232
rect 28816 27172 28820 27228
rect 28820 27172 28876 27228
rect 28876 27172 28880 27228
rect 28816 27168 28880 27172
rect 28896 27228 28960 27232
rect 28896 27172 28900 27228
rect 28900 27172 28956 27228
rect 28956 27172 28960 27228
rect 28896 27168 28960 27172
rect 28976 27228 29040 27232
rect 28976 27172 28980 27228
rect 28980 27172 29036 27228
rect 29036 27172 29040 27228
rect 28976 27168 29040 27172
rect 4425 26684 4489 26688
rect 4425 26628 4429 26684
rect 4429 26628 4485 26684
rect 4485 26628 4489 26684
rect 4425 26624 4489 26628
rect 4505 26684 4569 26688
rect 4505 26628 4509 26684
rect 4509 26628 4565 26684
rect 4565 26628 4569 26684
rect 4505 26624 4569 26628
rect 4585 26684 4649 26688
rect 4585 26628 4589 26684
rect 4589 26628 4645 26684
rect 4645 26628 4649 26684
rect 4585 26624 4649 26628
rect 4665 26684 4729 26688
rect 4665 26628 4669 26684
rect 4669 26628 4725 26684
rect 4725 26628 4729 26684
rect 4665 26624 4729 26628
rect 11371 26684 11435 26688
rect 11371 26628 11375 26684
rect 11375 26628 11431 26684
rect 11431 26628 11435 26684
rect 11371 26624 11435 26628
rect 11451 26684 11515 26688
rect 11451 26628 11455 26684
rect 11455 26628 11511 26684
rect 11511 26628 11515 26684
rect 11451 26624 11515 26628
rect 11531 26684 11595 26688
rect 11531 26628 11535 26684
rect 11535 26628 11591 26684
rect 11591 26628 11595 26684
rect 11531 26624 11595 26628
rect 11611 26684 11675 26688
rect 11611 26628 11615 26684
rect 11615 26628 11671 26684
rect 11671 26628 11675 26684
rect 11611 26624 11675 26628
rect 18317 26684 18381 26688
rect 18317 26628 18321 26684
rect 18321 26628 18377 26684
rect 18377 26628 18381 26684
rect 18317 26624 18381 26628
rect 18397 26684 18461 26688
rect 18397 26628 18401 26684
rect 18401 26628 18457 26684
rect 18457 26628 18461 26684
rect 18397 26624 18461 26628
rect 18477 26684 18541 26688
rect 18477 26628 18481 26684
rect 18481 26628 18537 26684
rect 18537 26628 18541 26684
rect 18477 26624 18541 26628
rect 18557 26684 18621 26688
rect 18557 26628 18561 26684
rect 18561 26628 18617 26684
rect 18617 26628 18621 26684
rect 18557 26624 18621 26628
rect 25263 26684 25327 26688
rect 25263 26628 25267 26684
rect 25267 26628 25323 26684
rect 25323 26628 25327 26684
rect 25263 26624 25327 26628
rect 25343 26684 25407 26688
rect 25343 26628 25347 26684
rect 25347 26628 25403 26684
rect 25403 26628 25407 26684
rect 25343 26624 25407 26628
rect 25423 26684 25487 26688
rect 25423 26628 25427 26684
rect 25427 26628 25483 26684
rect 25483 26628 25487 26684
rect 25423 26624 25487 26628
rect 25503 26684 25567 26688
rect 25503 26628 25507 26684
rect 25507 26628 25563 26684
rect 25563 26628 25567 26684
rect 25503 26624 25567 26628
rect 7898 26140 7962 26144
rect 7898 26084 7902 26140
rect 7902 26084 7958 26140
rect 7958 26084 7962 26140
rect 7898 26080 7962 26084
rect 7978 26140 8042 26144
rect 7978 26084 7982 26140
rect 7982 26084 8038 26140
rect 8038 26084 8042 26140
rect 7978 26080 8042 26084
rect 8058 26140 8122 26144
rect 8058 26084 8062 26140
rect 8062 26084 8118 26140
rect 8118 26084 8122 26140
rect 8058 26080 8122 26084
rect 8138 26140 8202 26144
rect 8138 26084 8142 26140
rect 8142 26084 8198 26140
rect 8198 26084 8202 26140
rect 8138 26080 8202 26084
rect 14844 26140 14908 26144
rect 14844 26084 14848 26140
rect 14848 26084 14904 26140
rect 14904 26084 14908 26140
rect 14844 26080 14908 26084
rect 14924 26140 14988 26144
rect 14924 26084 14928 26140
rect 14928 26084 14984 26140
rect 14984 26084 14988 26140
rect 14924 26080 14988 26084
rect 15004 26140 15068 26144
rect 15004 26084 15008 26140
rect 15008 26084 15064 26140
rect 15064 26084 15068 26140
rect 15004 26080 15068 26084
rect 15084 26140 15148 26144
rect 15084 26084 15088 26140
rect 15088 26084 15144 26140
rect 15144 26084 15148 26140
rect 15084 26080 15148 26084
rect 21790 26140 21854 26144
rect 21790 26084 21794 26140
rect 21794 26084 21850 26140
rect 21850 26084 21854 26140
rect 21790 26080 21854 26084
rect 21870 26140 21934 26144
rect 21870 26084 21874 26140
rect 21874 26084 21930 26140
rect 21930 26084 21934 26140
rect 21870 26080 21934 26084
rect 21950 26140 22014 26144
rect 21950 26084 21954 26140
rect 21954 26084 22010 26140
rect 22010 26084 22014 26140
rect 21950 26080 22014 26084
rect 22030 26140 22094 26144
rect 22030 26084 22034 26140
rect 22034 26084 22090 26140
rect 22090 26084 22094 26140
rect 22030 26080 22094 26084
rect 28736 26140 28800 26144
rect 28736 26084 28740 26140
rect 28740 26084 28796 26140
rect 28796 26084 28800 26140
rect 28736 26080 28800 26084
rect 28816 26140 28880 26144
rect 28816 26084 28820 26140
rect 28820 26084 28876 26140
rect 28876 26084 28880 26140
rect 28816 26080 28880 26084
rect 28896 26140 28960 26144
rect 28896 26084 28900 26140
rect 28900 26084 28956 26140
rect 28956 26084 28960 26140
rect 28896 26080 28960 26084
rect 28976 26140 29040 26144
rect 28976 26084 28980 26140
rect 28980 26084 29036 26140
rect 29036 26084 29040 26140
rect 28976 26080 29040 26084
rect 4425 25596 4489 25600
rect 4425 25540 4429 25596
rect 4429 25540 4485 25596
rect 4485 25540 4489 25596
rect 4425 25536 4489 25540
rect 4505 25596 4569 25600
rect 4505 25540 4509 25596
rect 4509 25540 4565 25596
rect 4565 25540 4569 25596
rect 4505 25536 4569 25540
rect 4585 25596 4649 25600
rect 4585 25540 4589 25596
rect 4589 25540 4645 25596
rect 4645 25540 4649 25596
rect 4585 25536 4649 25540
rect 4665 25596 4729 25600
rect 4665 25540 4669 25596
rect 4669 25540 4725 25596
rect 4725 25540 4729 25596
rect 4665 25536 4729 25540
rect 11371 25596 11435 25600
rect 11371 25540 11375 25596
rect 11375 25540 11431 25596
rect 11431 25540 11435 25596
rect 11371 25536 11435 25540
rect 11451 25596 11515 25600
rect 11451 25540 11455 25596
rect 11455 25540 11511 25596
rect 11511 25540 11515 25596
rect 11451 25536 11515 25540
rect 11531 25596 11595 25600
rect 11531 25540 11535 25596
rect 11535 25540 11591 25596
rect 11591 25540 11595 25596
rect 11531 25536 11595 25540
rect 11611 25596 11675 25600
rect 11611 25540 11615 25596
rect 11615 25540 11671 25596
rect 11671 25540 11675 25596
rect 11611 25536 11675 25540
rect 18317 25596 18381 25600
rect 18317 25540 18321 25596
rect 18321 25540 18377 25596
rect 18377 25540 18381 25596
rect 18317 25536 18381 25540
rect 18397 25596 18461 25600
rect 18397 25540 18401 25596
rect 18401 25540 18457 25596
rect 18457 25540 18461 25596
rect 18397 25536 18461 25540
rect 18477 25596 18541 25600
rect 18477 25540 18481 25596
rect 18481 25540 18537 25596
rect 18537 25540 18541 25596
rect 18477 25536 18541 25540
rect 18557 25596 18621 25600
rect 18557 25540 18561 25596
rect 18561 25540 18617 25596
rect 18617 25540 18621 25596
rect 18557 25536 18621 25540
rect 25263 25596 25327 25600
rect 25263 25540 25267 25596
rect 25267 25540 25323 25596
rect 25323 25540 25327 25596
rect 25263 25536 25327 25540
rect 25343 25596 25407 25600
rect 25343 25540 25347 25596
rect 25347 25540 25403 25596
rect 25403 25540 25407 25596
rect 25343 25536 25407 25540
rect 25423 25596 25487 25600
rect 25423 25540 25427 25596
rect 25427 25540 25483 25596
rect 25483 25540 25487 25596
rect 25423 25536 25487 25540
rect 25503 25596 25567 25600
rect 25503 25540 25507 25596
rect 25507 25540 25563 25596
rect 25563 25540 25567 25596
rect 25503 25536 25567 25540
rect 7898 25052 7962 25056
rect 7898 24996 7902 25052
rect 7902 24996 7958 25052
rect 7958 24996 7962 25052
rect 7898 24992 7962 24996
rect 7978 25052 8042 25056
rect 7978 24996 7982 25052
rect 7982 24996 8038 25052
rect 8038 24996 8042 25052
rect 7978 24992 8042 24996
rect 8058 25052 8122 25056
rect 8058 24996 8062 25052
rect 8062 24996 8118 25052
rect 8118 24996 8122 25052
rect 8058 24992 8122 24996
rect 8138 25052 8202 25056
rect 8138 24996 8142 25052
rect 8142 24996 8198 25052
rect 8198 24996 8202 25052
rect 8138 24992 8202 24996
rect 14844 25052 14908 25056
rect 14844 24996 14848 25052
rect 14848 24996 14904 25052
rect 14904 24996 14908 25052
rect 14844 24992 14908 24996
rect 14924 25052 14988 25056
rect 14924 24996 14928 25052
rect 14928 24996 14984 25052
rect 14984 24996 14988 25052
rect 14924 24992 14988 24996
rect 15004 25052 15068 25056
rect 15004 24996 15008 25052
rect 15008 24996 15064 25052
rect 15064 24996 15068 25052
rect 15004 24992 15068 24996
rect 15084 25052 15148 25056
rect 15084 24996 15088 25052
rect 15088 24996 15144 25052
rect 15144 24996 15148 25052
rect 15084 24992 15148 24996
rect 21790 25052 21854 25056
rect 21790 24996 21794 25052
rect 21794 24996 21850 25052
rect 21850 24996 21854 25052
rect 21790 24992 21854 24996
rect 21870 25052 21934 25056
rect 21870 24996 21874 25052
rect 21874 24996 21930 25052
rect 21930 24996 21934 25052
rect 21870 24992 21934 24996
rect 21950 25052 22014 25056
rect 21950 24996 21954 25052
rect 21954 24996 22010 25052
rect 22010 24996 22014 25052
rect 21950 24992 22014 24996
rect 22030 25052 22094 25056
rect 22030 24996 22034 25052
rect 22034 24996 22090 25052
rect 22090 24996 22094 25052
rect 22030 24992 22094 24996
rect 28736 25052 28800 25056
rect 28736 24996 28740 25052
rect 28740 24996 28796 25052
rect 28796 24996 28800 25052
rect 28736 24992 28800 24996
rect 28816 25052 28880 25056
rect 28816 24996 28820 25052
rect 28820 24996 28876 25052
rect 28876 24996 28880 25052
rect 28816 24992 28880 24996
rect 28896 25052 28960 25056
rect 28896 24996 28900 25052
rect 28900 24996 28956 25052
rect 28956 24996 28960 25052
rect 28896 24992 28960 24996
rect 28976 25052 29040 25056
rect 28976 24996 28980 25052
rect 28980 24996 29036 25052
rect 29036 24996 29040 25052
rect 28976 24992 29040 24996
rect 4425 24508 4489 24512
rect 4425 24452 4429 24508
rect 4429 24452 4485 24508
rect 4485 24452 4489 24508
rect 4425 24448 4489 24452
rect 4505 24508 4569 24512
rect 4505 24452 4509 24508
rect 4509 24452 4565 24508
rect 4565 24452 4569 24508
rect 4505 24448 4569 24452
rect 4585 24508 4649 24512
rect 4585 24452 4589 24508
rect 4589 24452 4645 24508
rect 4645 24452 4649 24508
rect 4585 24448 4649 24452
rect 4665 24508 4729 24512
rect 4665 24452 4669 24508
rect 4669 24452 4725 24508
rect 4725 24452 4729 24508
rect 4665 24448 4729 24452
rect 11371 24508 11435 24512
rect 11371 24452 11375 24508
rect 11375 24452 11431 24508
rect 11431 24452 11435 24508
rect 11371 24448 11435 24452
rect 11451 24508 11515 24512
rect 11451 24452 11455 24508
rect 11455 24452 11511 24508
rect 11511 24452 11515 24508
rect 11451 24448 11515 24452
rect 11531 24508 11595 24512
rect 11531 24452 11535 24508
rect 11535 24452 11591 24508
rect 11591 24452 11595 24508
rect 11531 24448 11595 24452
rect 11611 24508 11675 24512
rect 11611 24452 11615 24508
rect 11615 24452 11671 24508
rect 11671 24452 11675 24508
rect 11611 24448 11675 24452
rect 18317 24508 18381 24512
rect 18317 24452 18321 24508
rect 18321 24452 18377 24508
rect 18377 24452 18381 24508
rect 18317 24448 18381 24452
rect 18397 24508 18461 24512
rect 18397 24452 18401 24508
rect 18401 24452 18457 24508
rect 18457 24452 18461 24508
rect 18397 24448 18461 24452
rect 18477 24508 18541 24512
rect 18477 24452 18481 24508
rect 18481 24452 18537 24508
rect 18537 24452 18541 24508
rect 18477 24448 18541 24452
rect 18557 24508 18621 24512
rect 18557 24452 18561 24508
rect 18561 24452 18617 24508
rect 18617 24452 18621 24508
rect 18557 24448 18621 24452
rect 25263 24508 25327 24512
rect 25263 24452 25267 24508
rect 25267 24452 25323 24508
rect 25323 24452 25327 24508
rect 25263 24448 25327 24452
rect 25343 24508 25407 24512
rect 25343 24452 25347 24508
rect 25347 24452 25403 24508
rect 25403 24452 25407 24508
rect 25343 24448 25407 24452
rect 25423 24508 25487 24512
rect 25423 24452 25427 24508
rect 25427 24452 25483 24508
rect 25483 24452 25487 24508
rect 25423 24448 25487 24452
rect 25503 24508 25567 24512
rect 25503 24452 25507 24508
rect 25507 24452 25563 24508
rect 25563 24452 25567 24508
rect 25503 24448 25567 24452
rect 7898 23964 7962 23968
rect 7898 23908 7902 23964
rect 7902 23908 7958 23964
rect 7958 23908 7962 23964
rect 7898 23904 7962 23908
rect 7978 23964 8042 23968
rect 7978 23908 7982 23964
rect 7982 23908 8038 23964
rect 8038 23908 8042 23964
rect 7978 23904 8042 23908
rect 8058 23964 8122 23968
rect 8058 23908 8062 23964
rect 8062 23908 8118 23964
rect 8118 23908 8122 23964
rect 8058 23904 8122 23908
rect 8138 23964 8202 23968
rect 8138 23908 8142 23964
rect 8142 23908 8198 23964
rect 8198 23908 8202 23964
rect 8138 23904 8202 23908
rect 14844 23964 14908 23968
rect 14844 23908 14848 23964
rect 14848 23908 14904 23964
rect 14904 23908 14908 23964
rect 14844 23904 14908 23908
rect 14924 23964 14988 23968
rect 14924 23908 14928 23964
rect 14928 23908 14984 23964
rect 14984 23908 14988 23964
rect 14924 23904 14988 23908
rect 15004 23964 15068 23968
rect 15004 23908 15008 23964
rect 15008 23908 15064 23964
rect 15064 23908 15068 23964
rect 15004 23904 15068 23908
rect 15084 23964 15148 23968
rect 15084 23908 15088 23964
rect 15088 23908 15144 23964
rect 15144 23908 15148 23964
rect 15084 23904 15148 23908
rect 21790 23964 21854 23968
rect 21790 23908 21794 23964
rect 21794 23908 21850 23964
rect 21850 23908 21854 23964
rect 21790 23904 21854 23908
rect 21870 23964 21934 23968
rect 21870 23908 21874 23964
rect 21874 23908 21930 23964
rect 21930 23908 21934 23964
rect 21870 23904 21934 23908
rect 21950 23964 22014 23968
rect 21950 23908 21954 23964
rect 21954 23908 22010 23964
rect 22010 23908 22014 23964
rect 21950 23904 22014 23908
rect 22030 23964 22094 23968
rect 22030 23908 22034 23964
rect 22034 23908 22090 23964
rect 22090 23908 22094 23964
rect 22030 23904 22094 23908
rect 28736 23964 28800 23968
rect 28736 23908 28740 23964
rect 28740 23908 28796 23964
rect 28796 23908 28800 23964
rect 28736 23904 28800 23908
rect 28816 23964 28880 23968
rect 28816 23908 28820 23964
rect 28820 23908 28876 23964
rect 28876 23908 28880 23964
rect 28816 23904 28880 23908
rect 28896 23964 28960 23968
rect 28896 23908 28900 23964
rect 28900 23908 28956 23964
rect 28956 23908 28960 23964
rect 28896 23904 28960 23908
rect 28976 23964 29040 23968
rect 28976 23908 28980 23964
rect 28980 23908 29036 23964
rect 29036 23908 29040 23964
rect 28976 23904 29040 23908
rect 4425 23420 4489 23424
rect 4425 23364 4429 23420
rect 4429 23364 4485 23420
rect 4485 23364 4489 23420
rect 4425 23360 4489 23364
rect 4505 23420 4569 23424
rect 4505 23364 4509 23420
rect 4509 23364 4565 23420
rect 4565 23364 4569 23420
rect 4505 23360 4569 23364
rect 4585 23420 4649 23424
rect 4585 23364 4589 23420
rect 4589 23364 4645 23420
rect 4645 23364 4649 23420
rect 4585 23360 4649 23364
rect 4665 23420 4729 23424
rect 4665 23364 4669 23420
rect 4669 23364 4725 23420
rect 4725 23364 4729 23420
rect 4665 23360 4729 23364
rect 11371 23420 11435 23424
rect 11371 23364 11375 23420
rect 11375 23364 11431 23420
rect 11431 23364 11435 23420
rect 11371 23360 11435 23364
rect 11451 23420 11515 23424
rect 11451 23364 11455 23420
rect 11455 23364 11511 23420
rect 11511 23364 11515 23420
rect 11451 23360 11515 23364
rect 11531 23420 11595 23424
rect 11531 23364 11535 23420
rect 11535 23364 11591 23420
rect 11591 23364 11595 23420
rect 11531 23360 11595 23364
rect 11611 23420 11675 23424
rect 11611 23364 11615 23420
rect 11615 23364 11671 23420
rect 11671 23364 11675 23420
rect 11611 23360 11675 23364
rect 18317 23420 18381 23424
rect 18317 23364 18321 23420
rect 18321 23364 18377 23420
rect 18377 23364 18381 23420
rect 18317 23360 18381 23364
rect 18397 23420 18461 23424
rect 18397 23364 18401 23420
rect 18401 23364 18457 23420
rect 18457 23364 18461 23420
rect 18397 23360 18461 23364
rect 18477 23420 18541 23424
rect 18477 23364 18481 23420
rect 18481 23364 18537 23420
rect 18537 23364 18541 23420
rect 18477 23360 18541 23364
rect 18557 23420 18621 23424
rect 18557 23364 18561 23420
rect 18561 23364 18617 23420
rect 18617 23364 18621 23420
rect 18557 23360 18621 23364
rect 25263 23420 25327 23424
rect 25263 23364 25267 23420
rect 25267 23364 25323 23420
rect 25323 23364 25327 23420
rect 25263 23360 25327 23364
rect 25343 23420 25407 23424
rect 25343 23364 25347 23420
rect 25347 23364 25403 23420
rect 25403 23364 25407 23420
rect 25343 23360 25407 23364
rect 25423 23420 25487 23424
rect 25423 23364 25427 23420
rect 25427 23364 25483 23420
rect 25483 23364 25487 23420
rect 25423 23360 25487 23364
rect 25503 23420 25567 23424
rect 25503 23364 25507 23420
rect 25507 23364 25563 23420
rect 25563 23364 25567 23420
rect 25503 23360 25567 23364
rect 7898 22876 7962 22880
rect 7898 22820 7902 22876
rect 7902 22820 7958 22876
rect 7958 22820 7962 22876
rect 7898 22816 7962 22820
rect 7978 22876 8042 22880
rect 7978 22820 7982 22876
rect 7982 22820 8038 22876
rect 8038 22820 8042 22876
rect 7978 22816 8042 22820
rect 8058 22876 8122 22880
rect 8058 22820 8062 22876
rect 8062 22820 8118 22876
rect 8118 22820 8122 22876
rect 8058 22816 8122 22820
rect 8138 22876 8202 22880
rect 8138 22820 8142 22876
rect 8142 22820 8198 22876
rect 8198 22820 8202 22876
rect 8138 22816 8202 22820
rect 14844 22876 14908 22880
rect 14844 22820 14848 22876
rect 14848 22820 14904 22876
rect 14904 22820 14908 22876
rect 14844 22816 14908 22820
rect 14924 22876 14988 22880
rect 14924 22820 14928 22876
rect 14928 22820 14984 22876
rect 14984 22820 14988 22876
rect 14924 22816 14988 22820
rect 15004 22876 15068 22880
rect 15004 22820 15008 22876
rect 15008 22820 15064 22876
rect 15064 22820 15068 22876
rect 15004 22816 15068 22820
rect 15084 22876 15148 22880
rect 15084 22820 15088 22876
rect 15088 22820 15144 22876
rect 15144 22820 15148 22876
rect 15084 22816 15148 22820
rect 21790 22876 21854 22880
rect 21790 22820 21794 22876
rect 21794 22820 21850 22876
rect 21850 22820 21854 22876
rect 21790 22816 21854 22820
rect 21870 22876 21934 22880
rect 21870 22820 21874 22876
rect 21874 22820 21930 22876
rect 21930 22820 21934 22876
rect 21870 22816 21934 22820
rect 21950 22876 22014 22880
rect 21950 22820 21954 22876
rect 21954 22820 22010 22876
rect 22010 22820 22014 22876
rect 21950 22816 22014 22820
rect 22030 22876 22094 22880
rect 22030 22820 22034 22876
rect 22034 22820 22090 22876
rect 22090 22820 22094 22876
rect 22030 22816 22094 22820
rect 28736 22876 28800 22880
rect 28736 22820 28740 22876
rect 28740 22820 28796 22876
rect 28796 22820 28800 22876
rect 28736 22816 28800 22820
rect 28816 22876 28880 22880
rect 28816 22820 28820 22876
rect 28820 22820 28876 22876
rect 28876 22820 28880 22876
rect 28816 22816 28880 22820
rect 28896 22876 28960 22880
rect 28896 22820 28900 22876
rect 28900 22820 28956 22876
rect 28956 22820 28960 22876
rect 28896 22816 28960 22820
rect 28976 22876 29040 22880
rect 28976 22820 28980 22876
rect 28980 22820 29036 22876
rect 29036 22820 29040 22876
rect 28976 22816 29040 22820
rect 4425 22332 4489 22336
rect 4425 22276 4429 22332
rect 4429 22276 4485 22332
rect 4485 22276 4489 22332
rect 4425 22272 4489 22276
rect 4505 22332 4569 22336
rect 4505 22276 4509 22332
rect 4509 22276 4565 22332
rect 4565 22276 4569 22332
rect 4505 22272 4569 22276
rect 4585 22332 4649 22336
rect 4585 22276 4589 22332
rect 4589 22276 4645 22332
rect 4645 22276 4649 22332
rect 4585 22272 4649 22276
rect 4665 22332 4729 22336
rect 4665 22276 4669 22332
rect 4669 22276 4725 22332
rect 4725 22276 4729 22332
rect 4665 22272 4729 22276
rect 11371 22332 11435 22336
rect 11371 22276 11375 22332
rect 11375 22276 11431 22332
rect 11431 22276 11435 22332
rect 11371 22272 11435 22276
rect 11451 22332 11515 22336
rect 11451 22276 11455 22332
rect 11455 22276 11511 22332
rect 11511 22276 11515 22332
rect 11451 22272 11515 22276
rect 11531 22332 11595 22336
rect 11531 22276 11535 22332
rect 11535 22276 11591 22332
rect 11591 22276 11595 22332
rect 11531 22272 11595 22276
rect 11611 22332 11675 22336
rect 11611 22276 11615 22332
rect 11615 22276 11671 22332
rect 11671 22276 11675 22332
rect 11611 22272 11675 22276
rect 18317 22332 18381 22336
rect 18317 22276 18321 22332
rect 18321 22276 18377 22332
rect 18377 22276 18381 22332
rect 18317 22272 18381 22276
rect 18397 22332 18461 22336
rect 18397 22276 18401 22332
rect 18401 22276 18457 22332
rect 18457 22276 18461 22332
rect 18397 22272 18461 22276
rect 18477 22332 18541 22336
rect 18477 22276 18481 22332
rect 18481 22276 18537 22332
rect 18537 22276 18541 22332
rect 18477 22272 18541 22276
rect 18557 22332 18621 22336
rect 18557 22276 18561 22332
rect 18561 22276 18617 22332
rect 18617 22276 18621 22332
rect 18557 22272 18621 22276
rect 25263 22332 25327 22336
rect 25263 22276 25267 22332
rect 25267 22276 25323 22332
rect 25323 22276 25327 22332
rect 25263 22272 25327 22276
rect 25343 22332 25407 22336
rect 25343 22276 25347 22332
rect 25347 22276 25403 22332
rect 25403 22276 25407 22332
rect 25343 22272 25407 22276
rect 25423 22332 25487 22336
rect 25423 22276 25427 22332
rect 25427 22276 25483 22332
rect 25483 22276 25487 22332
rect 25423 22272 25487 22276
rect 25503 22332 25567 22336
rect 25503 22276 25507 22332
rect 25507 22276 25563 22332
rect 25563 22276 25567 22332
rect 25503 22272 25567 22276
rect 7898 21788 7962 21792
rect 7898 21732 7902 21788
rect 7902 21732 7958 21788
rect 7958 21732 7962 21788
rect 7898 21728 7962 21732
rect 7978 21788 8042 21792
rect 7978 21732 7982 21788
rect 7982 21732 8038 21788
rect 8038 21732 8042 21788
rect 7978 21728 8042 21732
rect 8058 21788 8122 21792
rect 8058 21732 8062 21788
rect 8062 21732 8118 21788
rect 8118 21732 8122 21788
rect 8058 21728 8122 21732
rect 8138 21788 8202 21792
rect 8138 21732 8142 21788
rect 8142 21732 8198 21788
rect 8198 21732 8202 21788
rect 8138 21728 8202 21732
rect 14844 21788 14908 21792
rect 14844 21732 14848 21788
rect 14848 21732 14904 21788
rect 14904 21732 14908 21788
rect 14844 21728 14908 21732
rect 14924 21788 14988 21792
rect 14924 21732 14928 21788
rect 14928 21732 14984 21788
rect 14984 21732 14988 21788
rect 14924 21728 14988 21732
rect 15004 21788 15068 21792
rect 15004 21732 15008 21788
rect 15008 21732 15064 21788
rect 15064 21732 15068 21788
rect 15004 21728 15068 21732
rect 15084 21788 15148 21792
rect 15084 21732 15088 21788
rect 15088 21732 15144 21788
rect 15144 21732 15148 21788
rect 15084 21728 15148 21732
rect 21790 21788 21854 21792
rect 21790 21732 21794 21788
rect 21794 21732 21850 21788
rect 21850 21732 21854 21788
rect 21790 21728 21854 21732
rect 21870 21788 21934 21792
rect 21870 21732 21874 21788
rect 21874 21732 21930 21788
rect 21930 21732 21934 21788
rect 21870 21728 21934 21732
rect 21950 21788 22014 21792
rect 21950 21732 21954 21788
rect 21954 21732 22010 21788
rect 22010 21732 22014 21788
rect 21950 21728 22014 21732
rect 22030 21788 22094 21792
rect 22030 21732 22034 21788
rect 22034 21732 22090 21788
rect 22090 21732 22094 21788
rect 22030 21728 22094 21732
rect 28736 21788 28800 21792
rect 28736 21732 28740 21788
rect 28740 21732 28796 21788
rect 28796 21732 28800 21788
rect 28736 21728 28800 21732
rect 28816 21788 28880 21792
rect 28816 21732 28820 21788
rect 28820 21732 28876 21788
rect 28876 21732 28880 21788
rect 28816 21728 28880 21732
rect 28896 21788 28960 21792
rect 28896 21732 28900 21788
rect 28900 21732 28956 21788
rect 28956 21732 28960 21788
rect 28896 21728 28960 21732
rect 28976 21788 29040 21792
rect 28976 21732 28980 21788
rect 28980 21732 29036 21788
rect 29036 21732 29040 21788
rect 28976 21728 29040 21732
rect 4425 21244 4489 21248
rect 4425 21188 4429 21244
rect 4429 21188 4485 21244
rect 4485 21188 4489 21244
rect 4425 21184 4489 21188
rect 4505 21244 4569 21248
rect 4505 21188 4509 21244
rect 4509 21188 4565 21244
rect 4565 21188 4569 21244
rect 4505 21184 4569 21188
rect 4585 21244 4649 21248
rect 4585 21188 4589 21244
rect 4589 21188 4645 21244
rect 4645 21188 4649 21244
rect 4585 21184 4649 21188
rect 4665 21244 4729 21248
rect 4665 21188 4669 21244
rect 4669 21188 4725 21244
rect 4725 21188 4729 21244
rect 4665 21184 4729 21188
rect 11371 21244 11435 21248
rect 11371 21188 11375 21244
rect 11375 21188 11431 21244
rect 11431 21188 11435 21244
rect 11371 21184 11435 21188
rect 11451 21244 11515 21248
rect 11451 21188 11455 21244
rect 11455 21188 11511 21244
rect 11511 21188 11515 21244
rect 11451 21184 11515 21188
rect 11531 21244 11595 21248
rect 11531 21188 11535 21244
rect 11535 21188 11591 21244
rect 11591 21188 11595 21244
rect 11531 21184 11595 21188
rect 11611 21244 11675 21248
rect 11611 21188 11615 21244
rect 11615 21188 11671 21244
rect 11671 21188 11675 21244
rect 11611 21184 11675 21188
rect 18317 21244 18381 21248
rect 18317 21188 18321 21244
rect 18321 21188 18377 21244
rect 18377 21188 18381 21244
rect 18317 21184 18381 21188
rect 18397 21244 18461 21248
rect 18397 21188 18401 21244
rect 18401 21188 18457 21244
rect 18457 21188 18461 21244
rect 18397 21184 18461 21188
rect 18477 21244 18541 21248
rect 18477 21188 18481 21244
rect 18481 21188 18537 21244
rect 18537 21188 18541 21244
rect 18477 21184 18541 21188
rect 18557 21244 18621 21248
rect 18557 21188 18561 21244
rect 18561 21188 18617 21244
rect 18617 21188 18621 21244
rect 18557 21184 18621 21188
rect 25263 21244 25327 21248
rect 25263 21188 25267 21244
rect 25267 21188 25323 21244
rect 25323 21188 25327 21244
rect 25263 21184 25327 21188
rect 25343 21244 25407 21248
rect 25343 21188 25347 21244
rect 25347 21188 25403 21244
rect 25403 21188 25407 21244
rect 25343 21184 25407 21188
rect 25423 21244 25487 21248
rect 25423 21188 25427 21244
rect 25427 21188 25483 21244
rect 25483 21188 25487 21244
rect 25423 21184 25487 21188
rect 25503 21244 25567 21248
rect 25503 21188 25507 21244
rect 25507 21188 25563 21244
rect 25563 21188 25567 21244
rect 25503 21184 25567 21188
rect 7898 20700 7962 20704
rect 7898 20644 7902 20700
rect 7902 20644 7958 20700
rect 7958 20644 7962 20700
rect 7898 20640 7962 20644
rect 7978 20700 8042 20704
rect 7978 20644 7982 20700
rect 7982 20644 8038 20700
rect 8038 20644 8042 20700
rect 7978 20640 8042 20644
rect 8058 20700 8122 20704
rect 8058 20644 8062 20700
rect 8062 20644 8118 20700
rect 8118 20644 8122 20700
rect 8058 20640 8122 20644
rect 8138 20700 8202 20704
rect 8138 20644 8142 20700
rect 8142 20644 8198 20700
rect 8198 20644 8202 20700
rect 8138 20640 8202 20644
rect 14844 20700 14908 20704
rect 14844 20644 14848 20700
rect 14848 20644 14904 20700
rect 14904 20644 14908 20700
rect 14844 20640 14908 20644
rect 14924 20700 14988 20704
rect 14924 20644 14928 20700
rect 14928 20644 14984 20700
rect 14984 20644 14988 20700
rect 14924 20640 14988 20644
rect 15004 20700 15068 20704
rect 15004 20644 15008 20700
rect 15008 20644 15064 20700
rect 15064 20644 15068 20700
rect 15004 20640 15068 20644
rect 15084 20700 15148 20704
rect 15084 20644 15088 20700
rect 15088 20644 15144 20700
rect 15144 20644 15148 20700
rect 15084 20640 15148 20644
rect 21790 20700 21854 20704
rect 21790 20644 21794 20700
rect 21794 20644 21850 20700
rect 21850 20644 21854 20700
rect 21790 20640 21854 20644
rect 21870 20700 21934 20704
rect 21870 20644 21874 20700
rect 21874 20644 21930 20700
rect 21930 20644 21934 20700
rect 21870 20640 21934 20644
rect 21950 20700 22014 20704
rect 21950 20644 21954 20700
rect 21954 20644 22010 20700
rect 22010 20644 22014 20700
rect 21950 20640 22014 20644
rect 22030 20700 22094 20704
rect 22030 20644 22034 20700
rect 22034 20644 22090 20700
rect 22090 20644 22094 20700
rect 22030 20640 22094 20644
rect 28736 20700 28800 20704
rect 28736 20644 28740 20700
rect 28740 20644 28796 20700
rect 28796 20644 28800 20700
rect 28736 20640 28800 20644
rect 28816 20700 28880 20704
rect 28816 20644 28820 20700
rect 28820 20644 28876 20700
rect 28876 20644 28880 20700
rect 28816 20640 28880 20644
rect 28896 20700 28960 20704
rect 28896 20644 28900 20700
rect 28900 20644 28956 20700
rect 28956 20644 28960 20700
rect 28896 20640 28960 20644
rect 28976 20700 29040 20704
rect 28976 20644 28980 20700
rect 28980 20644 29036 20700
rect 29036 20644 29040 20700
rect 28976 20640 29040 20644
rect 4425 20156 4489 20160
rect 4425 20100 4429 20156
rect 4429 20100 4485 20156
rect 4485 20100 4489 20156
rect 4425 20096 4489 20100
rect 4505 20156 4569 20160
rect 4505 20100 4509 20156
rect 4509 20100 4565 20156
rect 4565 20100 4569 20156
rect 4505 20096 4569 20100
rect 4585 20156 4649 20160
rect 4585 20100 4589 20156
rect 4589 20100 4645 20156
rect 4645 20100 4649 20156
rect 4585 20096 4649 20100
rect 4665 20156 4729 20160
rect 4665 20100 4669 20156
rect 4669 20100 4725 20156
rect 4725 20100 4729 20156
rect 4665 20096 4729 20100
rect 11371 20156 11435 20160
rect 11371 20100 11375 20156
rect 11375 20100 11431 20156
rect 11431 20100 11435 20156
rect 11371 20096 11435 20100
rect 11451 20156 11515 20160
rect 11451 20100 11455 20156
rect 11455 20100 11511 20156
rect 11511 20100 11515 20156
rect 11451 20096 11515 20100
rect 11531 20156 11595 20160
rect 11531 20100 11535 20156
rect 11535 20100 11591 20156
rect 11591 20100 11595 20156
rect 11531 20096 11595 20100
rect 11611 20156 11675 20160
rect 11611 20100 11615 20156
rect 11615 20100 11671 20156
rect 11671 20100 11675 20156
rect 11611 20096 11675 20100
rect 18317 20156 18381 20160
rect 18317 20100 18321 20156
rect 18321 20100 18377 20156
rect 18377 20100 18381 20156
rect 18317 20096 18381 20100
rect 18397 20156 18461 20160
rect 18397 20100 18401 20156
rect 18401 20100 18457 20156
rect 18457 20100 18461 20156
rect 18397 20096 18461 20100
rect 18477 20156 18541 20160
rect 18477 20100 18481 20156
rect 18481 20100 18537 20156
rect 18537 20100 18541 20156
rect 18477 20096 18541 20100
rect 18557 20156 18621 20160
rect 18557 20100 18561 20156
rect 18561 20100 18617 20156
rect 18617 20100 18621 20156
rect 18557 20096 18621 20100
rect 25263 20156 25327 20160
rect 25263 20100 25267 20156
rect 25267 20100 25323 20156
rect 25323 20100 25327 20156
rect 25263 20096 25327 20100
rect 25343 20156 25407 20160
rect 25343 20100 25347 20156
rect 25347 20100 25403 20156
rect 25403 20100 25407 20156
rect 25343 20096 25407 20100
rect 25423 20156 25487 20160
rect 25423 20100 25427 20156
rect 25427 20100 25483 20156
rect 25483 20100 25487 20156
rect 25423 20096 25487 20100
rect 25503 20156 25567 20160
rect 25503 20100 25507 20156
rect 25507 20100 25563 20156
rect 25563 20100 25567 20156
rect 25503 20096 25567 20100
rect 7898 19612 7962 19616
rect 7898 19556 7902 19612
rect 7902 19556 7958 19612
rect 7958 19556 7962 19612
rect 7898 19552 7962 19556
rect 7978 19612 8042 19616
rect 7978 19556 7982 19612
rect 7982 19556 8038 19612
rect 8038 19556 8042 19612
rect 7978 19552 8042 19556
rect 8058 19612 8122 19616
rect 8058 19556 8062 19612
rect 8062 19556 8118 19612
rect 8118 19556 8122 19612
rect 8058 19552 8122 19556
rect 8138 19612 8202 19616
rect 8138 19556 8142 19612
rect 8142 19556 8198 19612
rect 8198 19556 8202 19612
rect 8138 19552 8202 19556
rect 14844 19612 14908 19616
rect 14844 19556 14848 19612
rect 14848 19556 14904 19612
rect 14904 19556 14908 19612
rect 14844 19552 14908 19556
rect 14924 19612 14988 19616
rect 14924 19556 14928 19612
rect 14928 19556 14984 19612
rect 14984 19556 14988 19612
rect 14924 19552 14988 19556
rect 15004 19612 15068 19616
rect 15004 19556 15008 19612
rect 15008 19556 15064 19612
rect 15064 19556 15068 19612
rect 15004 19552 15068 19556
rect 15084 19612 15148 19616
rect 15084 19556 15088 19612
rect 15088 19556 15144 19612
rect 15144 19556 15148 19612
rect 15084 19552 15148 19556
rect 21790 19612 21854 19616
rect 21790 19556 21794 19612
rect 21794 19556 21850 19612
rect 21850 19556 21854 19612
rect 21790 19552 21854 19556
rect 21870 19612 21934 19616
rect 21870 19556 21874 19612
rect 21874 19556 21930 19612
rect 21930 19556 21934 19612
rect 21870 19552 21934 19556
rect 21950 19612 22014 19616
rect 21950 19556 21954 19612
rect 21954 19556 22010 19612
rect 22010 19556 22014 19612
rect 21950 19552 22014 19556
rect 22030 19612 22094 19616
rect 22030 19556 22034 19612
rect 22034 19556 22090 19612
rect 22090 19556 22094 19612
rect 22030 19552 22094 19556
rect 28736 19612 28800 19616
rect 28736 19556 28740 19612
rect 28740 19556 28796 19612
rect 28796 19556 28800 19612
rect 28736 19552 28800 19556
rect 28816 19612 28880 19616
rect 28816 19556 28820 19612
rect 28820 19556 28876 19612
rect 28876 19556 28880 19612
rect 28816 19552 28880 19556
rect 28896 19612 28960 19616
rect 28896 19556 28900 19612
rect 28900 19556 28956 19612
rect 28956 19556 28960 19612
rect 28896 19552 28960 19556
rect 28976 19612 29040 19616
rect 28976 19556 28980 19612
rect 28980 19556 29036 19612
rect 29036 19556 29040 19612
rect 28976 19552 29040 19556
rect 4425 19068 4489 19072
rect 4425 19012 4429 19068
rect 4429 19012 4485 19068
rect 4485 19012 4489 19068
rect 4425 19008 4489 19012
rect 4505 19068 4569 19072
rect 4505 19012 4509 19068
rect 4509 19012 4565 19068
rect 4565 19012 4569 19068
rect 4505 19008 4569 19012
rect 4585 19068 4649 19072
rect 4585 19012 4589 19068
rect 4589 19012 4645 19068
rect 4645 19012 4649 19068
rect 4585 19008 4649 19012
rect 4665 19068 4729 19072
rect 4665 19012 4669 19068
rect 4669 19012 4725 19068
rect 4725 19012 4729 19068
rect 4665 19008 4729 19012
rect 11371 19068 11435 19072
rect 11371 19012 11375 19068
rect 11375 19012 11431 19068
rect 11431 19012 11435 19068
rect 11371 19008 11435 19012
rect 11451 19068 11515 19072
rect 11451 19012 11455 19068
rect 11455 19012 11511 19068
rect 11511 19012 11515 19068
rect 11451 19008 11515 19012
rect 11531 19068 11595 19072
rect 11531 19012 11535 19068
rect 11535 19012 11591 19068
rect 11591 19012 11595 19068
rect 11531 19008 11595 19012
rect 11611 19068 11675 19072
rect 11611 19012 11615 19068
rect 11615 19012 11671 19068
rect 11671 19012 11675 19068
rect 11611 19008 11675 19012
rect 18317 19068 18381 19072
rect 18317 19012 18321 19068
rect 18321 19012 18377 19068
rect 18377 19012 18381 19068
rect 18317 19008 18381 19012
rect 18397 19068 18461 19072
rect 18397 19012 18401 19068
rect 18401 19012 18457 19068
rect 18457 19012 18461 19068
rect 18397 19008 18461 19012
rect 18477 19068 18541 19072
rect 18477 19012 18481 19068
rect 18481 19012 18537 19068
rect 18537 19012 18541 19068
rect 18477 19008 18541 19012
rect 18557 19068 18621 19072
rect 18557 19012 18561 19068
rect 18561 19012 18617 19068
rect 18617 19012 18621 19068
rect 18557 19008 18621 19012
rect 25263 19068 25327 19072
rect 25263 19012 25267 19068
rect 25267 19012 25323 19068
rect 25323 19012 25327 19068
rect 25263 19008 25327 19012
rect 25343 19068 25407 19072
rect 25343 19012 25347 19068
rect 25347 19012 25403 19068
rect 25403 19012 25407 19068
rect 25343 19008 25407 19012
rect 25423 19068 25487 19072
rect 25423 19012 25427 19068
rect 25427 19012 25483 19068
rect 25483 19012 25487 19068
rect 25423 19008 25487 19012
rect 25503 19068 25567 19072
rect 25503 19012 25507 19068
rect 25507 19012 25563 19068
rect 25563 19012 25567 19068
rect 25503 19008 25567 19012
rect 7898 18524 7962 18528
rect 7898 18468 7902 18524
rect 7902 18468 7958 18524
rect 7958 18468 7962 18524
rect 7898 18464 7962 18468
rect 7978 18524 8042 18528
rect 7978 18468 7982 18524
rect 7982 18468 8038 18524
rect 8038 18468 8042 18524
rect 7978 18464 8042 18468
rect 8058 18524 8122 18528
rect 8058 18468 8062 18524
rect 8062 18468 8118 18524
rect 8118 18468 8122 18524
rect 8058 18464 8122 18468
rect 8138 18524 8202 18528
rect 8138 18468 8142 18524
rect 8142 18468 8198 18524
rect 8198 18468 8202 18524
rect 8138 18464 8202 18468
rect 14844 18524 14908 18528
rect 14844 18468 14848 18524
rect 14848 18468 14904 18524
rect 14904 18468 14908 18524
rect 14844 18464 14908 18468
rect 14924 18524 14988 18528
rect 14924 18468 14928 18524
rect 14928 18468 14984 18524
rect 14984 18468 14988 18524
rect 14924 18464 14988 18468
rect 15004 18524 15068 18528
rect 15004 18468 15008 18524
rect 15008 18468 15064 18524
rect 15064 18468 15068 18524
rect 15004 18464 15068 18468
rect 15084 18524 15148 18528
rect 15084 18468 15088 18524
rect 15088 18468 15144 18524
rect 15144 18468 15148 18524
rect 15084 18464 15148 18468
rect 21790 18524 21854 18528
rect 21790 18468 21794 18524
rect 21794 18468 21850 18524
rect 21850 18468 21854 18524
rect 21790 18464 21854 18468
rect 21870 18524 21934 18528
rect 21870 18468 21874 18524
rect 21874 18468 21930 18524
rect 21930 18468 21934 18524
rect 21870 18464 21934 18468
rect 21950 18524 22014 18528
rect 21950 18468 21954 18524
rect 21954 18468 22010 18524
rect 22010 18468 22014 18524
rect 21950 18464 22014 18468
rect 22030 18524 22094 18528
rect 22030 18468 22034 18524
rect 22034 18468 22090 18524
rect 22090 18468 22094 18524
rect 22030 18464 22094 18468
rect 28736 18524 28800 18528
rect 28736 18468 28740 18524
rect 28740 18468 28796 18524
rect 28796 18468 28800 18524
rect 28736 18464 28800 18468
rect 28816 18524 28880 18528
rect 28816 18468 28820 18524
rect 28820 18468 28876 18524
rect 28876 18468 28880 18524
rect 28816 18464 28880 18468
rect 28896 18524 28960 18528
rect 28896 18468 28900 18524
rect 28900 18468 28956 18524
rect 28956 18468 28960 18524
rect 28896 18464 28960 18468
rect 28976 18524 29040 18528
rect 28976 18468 28980 18524
rect 28980 18468 29036 18524
rect 29036 18468 29040 18524
rect 28976 18464 29040 18468
rect 4425 17980 4489 17984
rect 4425 17924 4429 17980
rect 4429 17924 4485 17980
rect 4485 17924 4489 17980
rect 4425 17920 4489 17924
rect 4505 17980 4569 17984
rect 4505 17924 4509 17980
rect 4509 17924 4565 17980
rect 4565 17924 4569 17980
rect 4505 17920 4569 17924
rect 4585 17980 4649 17984
rect 4585 17924 4589 17980
rect 4589 17924 4645 17980
rect 4645 17924 4649 17980
rect 4585 17920 4649 17924
rect 4665 17980 4729 17984
rect 4665 17924 4669 17980
rect 4669 17924 4725 17980
rect 4725 17924 4729 17980
rect 4665 17920 4729 17924
rect 11371 17980 11435 17984
rect 11371 17924 11375 17980
rect 11375 17924 11431 17980
rect 11431 17924 11435 17980
rect 11371 17920 11435 17924
rect 11451 17980 11515 17984
rect 11451 17924 11455 17980
rect 11455 17924 11511 17980
rect 11511 17924 11515 17980
rect 11451 17920 11515 17924
rect 11531 17980 11595 17984
rect 11531 17924 11535 17980
rect 11535 17924 11591 17980
rect 11591 17924 11595 17980
rect 11531 17920 11595 17924
rect 11611 17980 11675 17984
rect 11611 17924 11615 17980
rect 11615 17924 11671 17980
rect 11671 17924 11675 17980
rect 11611 17920 11675 17924
rect 18317 17980 18381 17984
rect 18317 17924 18321 17980
rect 18321 17924 18377 17980
rect 18377 17924 18381 17980
rect 18317 17920 18381 17924
rect 18397 17980 18461 17984
rect 18397 17924 18401 17980
rect 18401 17924 18457 17980
rect 18457 17924 18461 17980
rect 18397 17920 18461 17924
rect 18477 17980 18541 17984
rect 18477 17924 18481 17980
rect 18481 17924 18537 17980
rect 18537 17924 18541 17980
rect 18477 17920 18541 17924
rect 18557 17980 18621 17984
rect 18557 17924 18561 17980
rect 18561 17924 18617 17980
rect 18617 17924 18621 17980
rect 18557 17920 18621 17924
rect 25263 17980 25327 17984
rect 25263 17924 25267 17980
rect 25267 17924 25323 17980
rect 25323 17924 25327 17980
rect 25263 17920 25327 17924
rect 25343 17980 25407 17984
rect 25343 17924 25347 17980
rect 25347 17924 25403 17980
rect 25403 17924 25407 17980
rect 25343 17920 25407 17924
rect 25423 17980 25487 17984
rect 25423 17924 25427 17980
rect 25427 17924 25483 17980
rect 25483 17924 25487 17980
rect 25423 17920 25487 17924
rect 25503 17980 25567 17984
rect 25503 17924 25507 17980
rect 25507 17924 25563 17980
rect 25563 17924 25567 17980
rect 25503 17920 25567 17924
rect 7898 17436 7962 17440
rect 7898 17380 7902 17436
rect 7902 17380 7958 17436
rect 7958 17380 7962 17436
rect 7898 17376 7962 17380
rect 7978 17436 8042 17440
rect 7978 17380 7982 17436
rect 7982 17380 8038 17436
rect 8038 17380 8042 17436
rect 7978 17376 8042 17380
rect 8058 17436 8122 17440
rect 8058 17380 8062 17436
rect 8062 17380 8118 17436
rect 8118 17380 8122 17436
rect 8058 17376 8122 17380
rect 8138 17436 8202 17440
rect 8138 17380 8142 17436
rect 8142 17380 8198 17436
rect 8198 17380 8202 17436
rect 8138 17376 8202 17380
rect 14844 17436 14908 17440
rect 14844 17380 14848 17436
rect 14848 17380 14904 17436
rect 14904 17380 14908 17436
rect 14844 17376 14908 17380
rect 14924 17436 14988 17440
rect 14924 17380 14928 17436
rect 14928 17380 14984 17436
rect 14984 17380 14988 17436
rect 14924 17376 14988 17380
rect 15004 17436 15068 17440
rect 15004 17380 15008 17436
rect 15008 17380 15064 17436
rect 15064 17380 15068 17436
rect 15004 17376 15068 17380
rect 15084 17436 15148 17440
rect 15084 17380 15088 17436
rect 15088 17380 15144 17436
rect 15144 17380 15148 17436
rect 15084 17376 15148 17380
rect 21790 17436 21854 17440
rect 21790 17380 21794 17436
rect 21794 17380 21850 17436
rect 21850 17380 21854 17436
rect 21790 17376 21854 17380
rect 21870 17436 21934 17440
rect 21870 17380 21874 17436
rect 21874 17380 21930 17436
rect 21930 17380 21934 17436
rect 21870 17376 21934 17380
rect 21950 17436 22014 17440
rect 21950 17380 21954 17436
rect 21954 17380 22010 17436
rect 22010 17380 22014 17436
rect 21950 17376 22014 17380
rect 22030 17436 22094 17440
rect 22030 17380 22034 17436
rect 22034 17380 22090 17436
rect 22090 17380 22094 17436
rect 22030 17376 22094 17380
rect 28736 17436 28800 17440
rect 28736 17380 28740 17436
rect 28740 17380 28796 17436
rect 28796 17380 28800 17436
rect 28736 17376 28800 17380
rect 28816 17436 28880 17440
rect 28816 17380 28820 17436
rect 28820 17380 28876 17436
rect 28876 17380 28880 17436
rect 28816 17376 28880 17380
rect 28896 17436 28960 17440
rect 28896 17380 28900 17436
rect 28900 17380 28956 17436
rect 28956 17380 28960 17436
rect 28896 17376 28960 17380
rect 28976 17436 29040 17440
rect 28976 17380 28980 17436
rect 28980 17380 29036 17436
rect 29036 17380 29040 17436
rect 28976 17376 29040 17380
rect 4425 16892 4489 16896
rect 4425 16836 4429 16892
rect 4429 16836 4485 16892
rect 4485 16836 4489 16892
rect 4425 16832 4489 16836
rect 4505 16892 4569 16896
rect 4505 16836 4509 16892
rect 4509 16836 4565 16892
rect 4565 16836 4569 16892
rect 4505 16832 4569 16836
rect 4585 16892 4649 16896
rect 4585 16836 4589 16892
rect 4589 16836 4645 16892
rect 4645 16836 4649 16892
rect 4585 16832 4649 16836
rect 4665 16892 4729 16896
rect 4665 16836 4669 16892
rect 4669 16836 4725 16892
rect 4725 16836 4729 16892
rect 4665 16832 4729 16836
rect 11371 16892 11435 16896
rect 11371 16836 11375 16892
rect 11375 16836 11431 16892
rect 11431 16836 11435 16892
rect 11371 16832 11435 16836
rect 11451 16892 11515 16896
rect 11451 16836 11455 16892
rect 11455 16836 11511 16892
rect 11511 16836 11515 16892
rect 11451 16832 11515 16836
rect 11531 16892 11595 16896
rect 11531 16836 11535 16892
rect 11535 16836 11591 16892
rect 11591 16836 11595 16892
rect 11531 16832 11595 16836
rect 11611 16892 11675 16896
rect 11611 16836 11615 16892
rect 11615 16836 11671 16892
rect 11671 16836 11675 16892
rect 11611 16832 11675 16836
rect 18317 16892 18381 16896
rect 18317 16836 18321 16892
rect 18321 16836 18377 16892
rect 18377 16836 18381 16892
rect 18317 16832 18381 16836
rect 18397 16892 18461 16896
rect 18397 16836 18401 16892
rect 18401 16836 18457 16892
rect 18457 16836 18461 16892
rect 18397 16832 18461 16836
rect 18477 16892 18541 16896
rect 18477 16836 18481 16892
rect 18481 16836 18537 16892
rect 18537 16836 18541 16892
rect 18477 16832 18541 16836
rect 18557 16892 18621 16896
rect 18557 16836 18561 16892
rect 18561 16836 18617 16892
rect 18617 16836 18621 16892
rect 18557 16832 18621 16836
rect 25263 16892 25327 16896
rect 25263 16836 25267 16892
rect 25267 16836 25323 16892
rect 25323 16836 25327 16892
rect 25263 16832 25327 16836
rect 25343 16892 25407 16896
rect 25343 16836 25347 16892
rect 25347 16836 25403 16892
rect 25403 16836 25407 16892
rect 25343 16832 25407 16836
rect 25423 16892 25487 16896
rect 25423 16836 25427 16892
rect 25427 16836 25483 16892
rect 25483 16836 25487 16892
rect 25423 16832 25487 16836
rect 25503 16892 25567 16896
rect 25503 16836 25507 16892
rect 25507 16836 25563 16892
rect 25563 16836 25567 16892
rect 25503 16832 25567 16836
rect 7898 16348 7962 16352
rect 7898 16292 7902 16348
rect 7902 16292 7958 16348
rect 7958 16292 7962 16348
rect 7898 16288 7962 16292
rect 7978 16348 8042 16352
rect 7978 16292 7982 16348
rect 7982 16292 8038 16348
rect 8038 16292 8042 16348
rect 7978 16288 8042 16292
rect 8058 16348 8122 16352
rect 8058 16292 8062 16348
rect 8062 16292 8118 16348
rect 8118 16292 8122 16348
rect 8058 16288 8122 16292
rect 8138 16348 8202 16352
rect 8138 16292 8142 16348
rect 8142 16292 8198 16348
rect 8198 16292 8202 16348
rect 8138 16288 8202 16292
rect 14844 16348 14908 16352
rect 14844 16292 14848 16348
rect 14848 16292 14904 16348
rect 14904 16292 14908 16348
rect 14844 16288 14908 16292
rect 14924 16348 14988 16352
rect 14924 16292 14928 16348
rect 14928 16292 14984 16348
rect 14984 16292 14988 16348
rect 14924 16288 14988 16292
rect 15004 16348 15068 16352
rect 15004 16292 15008 16348
rect 15008 16292 15064 16348
rect 15064 16292 15068 16348
rect 15004 16288 15068 16292
rect 15084 16348 15148 16352
rect 15084 16292 15088 16348
rect 15088 16292 15144 16348
rect 15144 16292 15148 16348
rect 15084 16288 15148 16292
rect 21790 16348 21854 16352
rect 21790 16292 21794 16348
rect 21794 16292 21850 16348
rect 21850 16292 21854 16348
rect 21790 16288 21854 16292
rect 21870 16348 21934 16352
rect 21870 16292 21874 16348
rect 21874 16292 21930 16348
rect 21930 16292 21934 16348
rect 21870 16288 21934 16292
rect 21950 16348 22014 16352
rect 21950 16292 21954 16348
rect 21954 16292 22010 16348
rect 22010 16292 22014 16348
rect 21950 16288 22014 16292
rect 22030 16348 22094 16352
rect 22030 16292 22034 16348
rect 22034 16292 22090 16348
rect 22090 16292 22094 16348
rect 22030 16288 22094 16292
rect 28736 16348 28800 16352
rect 28736 16292 28740 16348
rect 28740 16292 28796 16348
rect 28796 16292 28800 16348
rect 28736 16288 28800 16292
rect 28816 16348 28880 16352
rect 28816 16292 28820 16348
rect 28820 16292 28876 16348
rect 28876 16292 28880 16348
rect 28816 16288 28880 16292
rect 28896 16348 28960 16352
rect 28896 16292 28900 16348
rect 28900 16292 28956 16348
rect 28956 16292 28960 16348
rect 28896 16288 28960 16292
rect 28976 16348 29040 16352
rect 28976 16292 28980 16348
rect 28980 16292 29036 16348
rect 29036 16292 29040 16348
rect 28976 16288 29040 16292
rect 4425 15804 4489 15808
rect 4425 15748 4429 15804
rect 4429 15748 4485 15804
rect 4485 15748 4489 15804
rect 4425 15744 4489 15748
rect 4505 15804 4569 15808
rect 4505 15748 4509 15804
rect 4509 15748 4565 15804
rect 4565 15748 4569 15804
rect 4505 15744 4569 15748
rect 4585 15804 4649 15808
rect 4585 15748 4589 15804
rect 4589 15748 4645 15804
rect 4645 15748 4649 15804
rect 4585 15744 4649 15748
rect 4665 15804 4729 15808
rect 4665 15748 4669 15804
rect 4669 15748 4725 15804
rect 4725 15748 4729 15804
rect 4665 15744 4729 15748
rect 11371 15804 11435 15808
rect 11371 15748 11375 15804
rect 11375 15748 11431 15804
rect 11431 15748 11435 15804
rect 11371 15744 11435 15748
rect 11451 15804 11515 15808
rect 11451 15748 11455 15804
rect 11455 15748 11511 15804
rect 11511 15748 11515 15804
rect 11451 15744 11515 15748
rect 11531 15804 11595 15808
rect 11531 15748 11535 15804
rect 11535 15748 11591 15804
rect 11591 15748 11595 15804
rect 11531 15744 11595 15748
rect 11611 15804 11675 15808
rect 11611 15748 11615 15804
rect 11615 15748 11671 15804
rect 11671 15748 11675 15804
rect 11611 15744 11675 15748
rect 18317 15804 18381 15808
rect 18317 15748 18321 15804
rect 18321 15748 18377 15804
rect 18377 15748 18381 15804
rect 18317 15744 18381 15748
rect 18397 15804 18461 15808
rect 18397 15748 18401 15804
rect 18401 15748 18457 15804
rect 18457 15748 18461 15804
rect 18397 15744 18461 15748
rect 18477 15804 18541 15808
rect 18477 15748 18481 15804
rect 18481 15748 18537 15804
rect 18537 15748 18541 15804
rect 18477 15744 18541 15748
rect 18557 15804 18621 15808
rect 18557 15748 18561 15804
rect 18561 15748 18617 15804
rect 18617 15748 18621 15804
rect 18557 15744 18621 15748
rect 25263 15804 25327 15808
rect 25263 15748 25267 15804
rect 25267 15748 25323 15804
rect 25323 15748 25327 15804
rect 25263 15744 25327 15748
rect 25343 15804 25407 15808
rect 25343 15748 25347 15804
rect 25347 15748 25403 15804
rect 25403 15748 25407 15804
rect 25343 15744 25407 15748
rect 25423 15804 25487 15808
rect 25423 15748 25427 15804
rect 25427 15748 25483 15804
rect 25483 15748 25487 15804
rect 25423 15744 25487 15748
rect 25503 15804 25567 15808
rect 25503 15748 25507 15804
rect 25507 15748 25563 15804
rect 25563 15748 25567 15804
rect 25503 15744 25567 15748
rect 7898 15260 7962 15264
rect 7898 15204 7902 15260
rect 7902 15204 7958 15260
rect 7958 15204 7962 15260
rect 7898 15200 7962 15204
rect 7978 15260 8042 15264
rect 7978 15204 7982 15260
rect 7982 15204 8038 15260
rect 8038 15204 8042 15260
rect 7978 15200 8042 15204
rect 8058 15260 8122 15264
rect 8058 15204 8062 15260
rect 8062 15204 8118 15260
rect 8118 15204 8122 15260
rect 8058 15200 8122 15204
rect 8138 15260 8202 15264
rect 8138 15204 8142 15260
rect 8142 15204 8198 15260
rect 8198 15204 8202 15260
rect 8138 15200 8202 15204
rect 14844 15260 14908 15264
rect 14844 15204 14848 15260
rect 14848 15204 14904 15260
rect 14904 15204 14908 15260
rect 14844 15200 14908 15204
rect 14924 15260 14988 15264
rect 14924 15204 14928 15260
rect 14928 15204 14984 15260
rect 14984 15204 14988 15260
rect 14924 15200 14988 15204
rect 15004 15260 15068 15264
rect 15004 15204 15008 15260
rect 15008 15204 15064 15260
rect 15064 15204 15068 15260
rect 15004 15200 15068 15204
rect 15084 15260 15148 15264
rect 15084 15204 15088 15260
rect 15088 15204 15144 15260
rect 15144 15204 15148 15260
rect 15084 15200 15148 15204
rect 21790 15260 21854 15264
rect 21790 15204 21794 15260
rect 21794 15204 21850 15260
rect 21850 15204 21854 15260
rect 21790 15200 21854 15204
rect 21870 15260 21934 15264
rect 21870 15204 21874 15260
rect 21874 15204 21930 15260
rect 21930 15204 21934 15260
rect 21870 15200 21934 15204
rect 21950 15260 22014 15264
rect 21950 15204 21954 15260
rect 21954 15204 22010 15260
rect 22010 15204 22014 15260
rect 21950 15200 22014 15204
rect 22030 15260 22094 15264
rect 22030 15204 22034 15260
rect 22034 15204 22090 15260
rect 22090 15204 22094 15260
rect 22030 15200 22094 15204
rect 28736 15260 28800 15264
rect 28736 15204 28740 15260
rect 28740 15204 28796 15260
rect 28796 15204 28800 15260
rect 28736 15200 28800 15204
rect 28816 15260 28880 15264
rect 28816 15204 28820 15260
rect 28820 15204 28876 15260
rect 28876 15204 28880 15260
rect 28816 15200 28880 15204
rect 28896 15260 28960 15264
rect 28896 15204 28900 15260
rect 28900 15204 28956 15260
rect 28956 15204 28960 15260
rect 28896 15200 28960 15204
rect 28976 15260 29040 15264
rect 28976 15204 28980 15260
rect 28980 15204 29036 15260
rect 29036 15204 29040 15260
rect 28976 15200 29040 15204
rect 4425 14716 4489 14720
rect 4425 14660 4429 14716
rect 4429 14660 4485 14716
rect 4485 14660 4489 14716
rect 4425 14656 4489 14660
rect 4505 14716 4569 14720
rect 4505 14660 4509 14716
rect 4509 14660 4565 14716
rect 4565 14660 4569 14716
rect 4505 14656 4569 14660
rect 4585 14716 4649 14720
rect 4585 14660 4589 14716
rect 4589 14660 4645 14716
rect 4645 14660 4649 14716
rect 4585 14656 4649 14660
rect 4665 14716 4729 14720
rect 4665 14660 4669 14716
rect 4669 14660 4725 14716
rect 4725 14660 4729 14716
rect 4665 14656 4729 14660
rect 11371 14716 11435 14720
rect 11371 14660 11375 14716
rect 11375 14660 11431 14716
rect 11431 14660 11435 14716
rect 11371 14656 11435 14660
rect 11451 14716 11515 14720
rect 11451 14660 11455 14716
rect 11455 14660 11511 14716
rect 11511 14660 11515 14716
rect 11451 14656 11515 14660
rect 11531 14716 11595 14720
rect 11531 14660 11535 14716
rect 11535 14660 11591 14716
rect 11591 14660 11595 14716
rect 11531 14656 11595 14660
rect 11611 14716 11675 14720
rect 11611 14660 11615 14716
rect 11615 14660 11671 14716
rect 11671 14660 11675 14716
rect 11611 14656 11675 14660
rect 18317 14716 18381 14720
rect 18317 14660 18321 14716
rect 18321 14660 18377 14716
rect 18377 14660 18381 14716
rect 18317 14656 18381 14660
rect 18397 14716 18461 14720
rect 18397 14660 18401 14716
rect 18401 14660 18457 14716
rect 18457 14660 18461 14716
rect 18397 14656 18461 14660
rect 18477 14716 18541 14720
rect 18477 14660 18481 14716
rect 18481 14660 18537 14716
rect 18537 14660 18541 14716
rect 18477 14656 18541 14660
rect 18557 14716 18621 14720
rect 18557 14660 18561 14716
rect 18561 14660 18617 14716
rect 18617 14660 18621 14716
rect 18557 14656 18621 14660
rect 25263 14716 25327 14720
rect 25263 14660 25267 14716
rect 25267 14660 25323 14716
rect 25323 14660 25327 14716
rect 25263 14656 25327 14660
rect 25343 14716 25407 14720
rect 25343 14660 25347 14716
rect 25347 14660 25403 14716
rect 25403 14660 25407 14716
rect 25343 14656 25407 14660
rect 25423 14716 25487 14720
rect 25423 14660 25427 14716
rect 25427 14660 25483 14716
rect 25483 14660 25487 14716
rect 25423 14656 25487 14660
rect 25503 14716 25567 14720
rect 25503 14660 25507 14716
rect 25507 14660 25563 14716
rect 25563 14660 25567 14716
rect 25503 14656 25567 14660
rect 7898 14172 7962 14176
rect 7898 14116 7902 14172
rect 7902 14116 7958 14172
rect 7958 14116 7962 14172
rect 7898 14112 7962 14116
rect 7978 14172 8042 14176
rect 7978 14116 7982 14172
rect 7982 14116 8038 14172
rect 8038 14116 8042 14172
rect 7978 14112 8042 14116
rect 8058 14172 8122 14176
rect 8058 14116 8062 14172
rect 8062 14116 8118 14172
rect 8118 14116 8122 14172
rect 8058 14112 8122 14116
rect 8138 14172 8202 14176
rect 8138 14116 8142 14172
rect 8142 14116 8198 14172
rect 8198 14116 8202 14172
rect 8138 14112 8202 14116
rect 14844 14172 14908 14176
rect 14844 14116 14848 14172
rect 14848 14116 14904 14172
rect 14904 14116 14908 14172
rect 14844 14112 14908 14116
rect 14924 14172 14988 14176
rect 14924 14116 14928 14172
rect 14928 14116 14984 14172
rect 14984 14116 14988 14172
rect 14924 14112 14988 14116
rect 15004 14172 15068 14176
rect 15004 14116 15008 14172
rect 15008 14116 15064 14172
rect 15064 14116 15068 14172
rect 15004 14112 15068 14116
rect 15084 14172 15148 14176
rect 15084 14116 15088 14172
rect 15088 14116 15144 14172
rect 15144 14116 15148 14172
rect 15084 14112 15148 14116
rect 21790 14172 21854 14176
rect 21790 14116 21794 14172
rect 21794 14116 21850 14172
rect 21850 14116 21854 14172
rect 21790 14112 21854 14116
rect 21870 14172 21934 14176
rect 21870 14116 21874 14172
rect 21874 14116 21930 14172
rect 21930 14116 21934 14172
rect 21870 14112 21934 14116
rect 21950 14172 22014 14176
rect 21950 14116 21954 14172
rect 21954 14116 22010 14172
rect 22010 14116 22014 14172
rect 21950 14112 22014 14116
rect 22030 14172 22094 14176
rect 22030 14116 22034 14172
rect 22034 14116 22090 14172
rect 22090 14116 22094 14172
rect 22030 14112 22094 14116
rect 28736 14172 28800 14176
rect 28736 14116 28740 14172
rect 28740 14116 28796 14172
rect 28796 14116 28800 14172
rect 28736 14112 28800 14116
rect 28816 14172 28880 14176
rect 28816 14116 28820 14172
rect 28820 14116 28876 14172
rect 28876 14116 28880 14172
rect 28816 14112 28880 14116
rect 28896 14172 28960 14176
rect 28896 14116 28900 14172
rect 28900 14116 28956 14172
rect 28956 14116 28960 14172
rect 28896 14112 28960 14116
rect 28976 14172 29040 14176
rect 28976 14116 28980 14172
rect 28980 14116 29036 14172
rect 29036 14116 29040 14172
rect 28976 14112 29040 14116
rect 4425 13628 4489 13632
rect 4425 13572 4429 13628
rect 4429 13572 4485 13628
rect 4485 13572 4489 13628
rect 4425 13568 4489 13572
rect 4505 13628 4569 13632
rect 4505 13572 4509 13628
rect 4509 13572 4565 13628
rect 4565 13572 4569 13628
rect 4505 13568 4569 13572
rect 4585 13628 4649 13632
rect 4585 13572 4589 13628
rect 4589 13572 4645 13628
rect 4645 13572 4649 13628
rect 4585 13568 4649 13572
rect 4665 13628 4729 13632
rect 4665 13572 4669 13628
rect 4669 13572 4725 13628
rect 4725 13572 4729 13628
rect 4665 13568 4729 13572
rect 11371 13628 11435 13632
rect 11371 13572 11375 13628
rect 11375 13572 11431 13628
rect 11431 13572 11435 13628
rect 11371 13568 11435 13572
rect 11451 13628 11515 13632
rect 11451 13572 11455 13628
rect 11455 13572 11511 13628
rect 11511 13572 11515 13628
rect 11451 13568 11515 13572
rect 11531 13628 11595 13632
rect 11531 13572 11535 13628
rect 11535 13572 11591 13628
rect 11591 13572 11595 13628
rect 11531 13568 11595 13572
rect 11611 13628 11675 13632
rect 11611 13572 11615 13628
rect 11615 13572 11671 13628
rect 11671 13572 11675 13628
rect 11611 13568 11675 13572
rect 18317 13628 18381 13632
rect 18317 13572 18321 13628
rect 18321 13572 18377 13628
rect 18377 13572 18381 13628
rect 18317 13568 18381 13572
rect 18397 13628 18461 13632
rect 18397 13572 18401 13628
rect 18401 13572 18457 13628
rect 18457 13572 18461 13628
rect 18397 13568 18461 13572
rect 18477 13628 18541 13632
rect 18477 13572 18481 13628
rect 18481 13572 18537 13628
rect 18537 13572 18541 13628
rect 18477 13568 18541 13572
rect 18557 13628 18621 13632
rect 18557 13572 18561 13628
rect 18561 13572 18617 13628
rect 18617 13572 18621 13628
rect 18557 13568 18621 13572
rect 25263 13628 25327 13632
rect 25263 13572 25267 13628
rect 25267 13572 25323 13628
rect 25323 13572 25327 13628
rect 25263 13568 25327 13572
rect 25343 13628 25407 13632
rect 25343 13572 25347 13628
rect 25347 13572 25403 13628
rect 25403 13572 25407 13628
rect 25343 13568 25407 13572
rect 25423 13628 25487 13632
rect 25423 13572 25427 13628
rect 25427 13572 25483 13628
rect 25483 13572 25487 13628
rect 25423 13568 25487 13572
rect 25503 13628 25567 13632
rect 25503 13572 25507 13628
rect 25507 13572 25563 13628
rect 25563 13572 25567 13628
rect 25503 13568 25567 13572
rect 7898 13084 7962 13088
rect 7898 13028 7902 13084
rect 7902 13028 7958 13084
rect 7958 13028 7962 13084
rect 7898 13024 7962 13028
rect 7978 13084 8042 13088
rect 7978 13028 7982 13084
rect 7982 13028 8038 13084
rect 8038 13028 8042 13084
rect 7978 13024 8042 13028
rect 8058 13084 8122 13088
rect 8058 13028 8062 13084
rect 8062 13028 8118 13084
rect 8118 13028 8122 13084
rect 8058 13024 8122 13028
rect 8138 13084 8202 13088
rect 8138 13028 8142 13084
rect 8142 13028 8198 13084
rect 8198 13028 8202 13084
rect 8138 13024 8202 13028
rect 14844 13084 14908 13088
rect 14844 13028 14848 13084
rect 14848 13028 14904 13084
rect 14904 13028 14908 13084
rect 14844 13024 14908 13028
rect 14924 13084 14988 13088
rect 14924 13028 14928 13084
rect 14928 13028 14984 13084
rect 14984 13028 14988 13084
rect 14924 13024 14988 13028
rect 15004 13084 15068 13088
rect 15004 13028 15008 13084
rect 15008 13028 15064 13084
rect 15064 13028 15068 13084
rect 15004 13024 15068 13028
rect 15084 13084 15148 13088
rect 15084 13028 15088 13084
rect 15088 13028 15144 13084
rect 15144 13028 15148 13084
rect 15084 13024 15148 13028
rect 21790 13084 21854 13088
rect 21790 13028 21794 13084
rect 21794 13028 21850 13084
rect 21850 13028 21854 13084
rect 21790 13024 21854 13028
rect 21870 13084 21934 13088
rect 21870 13028 21874 13084
rect 21874 13028 21930 13084
rect 21930 13028 21934 13084
rect 21870 13024 21934 13028
rect 21950 13084 22014 13088
rect 21950 13028 21954 13084
rect 21954 13028 22010 13084
rect 22010 13028 22014 13084
rect 21950 13024 22014 13028
rect 22030 13084 22094 13088
rect 22030 13028 22034 13084
rect 22034 13028 22090 13084
rect 22090 13028 22094 13084
rect 22030 13024 22094 13028
rect 28736 13084 28800 13088
rect 28736 13028 28740 13084
rect 28740 13028 28796 13084
rect 28796 13028 28800 13084
rect 28736 13024 28800 13028
rect 28816 13084 28880 13088
rect 28816 13028 28820 13084
rect 28820 13028 28876 13084
rect 28876 13028 28880 13084
rect 28816 13024 28880 13028
rect 28896 13084 28960 13088
rect 28896 13028 28900 13084
rect 28900 13028 28956 13084
rect 28956 13028 28960 13084
rect 28896 13024 28960 13028
rect 28976 13084 29040 13088
rect 28976 13028 28980 13084
rect 28980 13028 29036 13084
rect 29036 13028 29040 13084
rect 28976 13024 29040 13028
rect 4425 12540 4489 12544
rect 4425 12484 4429 12540
rect 4429 12484 4485 12540
rect 4485 12484 4489 12540
rect 4425 12480 4489 12484
rect 4505 12540 4569 12544
rect 4505 12484 4509 12540
rect 4509 12484 4565 12540
rect 4565 12484 4569 12540
rect 4505 12480 4569 12484
rect 4585 12540 4649 12544
rect 4585 12484 4589 12540
rect 4589 12484 4645 12540
rect 4645 12484 4649 12540
rect 4585 12480 4649 12484
rect 4665 12540 4729 12544
rect 4665 12484 4669 12540
rect 4669 12484 4725 12540
rect 4725 12484 4729 12540
rect 4665 12480 4729 12484
rect 11371 12540 11435 12544
rect 11371 12484 11375 12540
rect 11375 12484 11431 12540
rect 11431 12484 11435 12540
rect 11371 12480 11435 12484
rect 11451 12540 11515 12544
rect 11451 12484 11455 12540
rect 11455 12484 11511 12540
rect 11511 12484 11515 12540
rect 11451 12480 11515 12484
rect 11531 12540 11595 12544
rect 11531 12484 11535 12540
rect 11535 12484 11591 12540
rect 11591 12484 11595 12540
rect 11531 12480 11595 12484
rect 11611 12540 11675 12544
rect 11611 12484 11615 12540
rect 11615 12484 11671 12540
rect 11671 12484 11675 12540
rect 11611 12480 11675 12484
rect 18317 12540 18381 12544
rect 18317 12484 18321 12540
rect 18321 12484 18377 12540
rect 18377 12484 18381 12540
rect 18317 12480 18381 12484
rect 18397 12540 18461 12544
rect 18397 12484 18401 12540
rect 18401 12484 18457 12540
rect 18457 12484 18461 12540
rect 18397 12480 18461 12484
rect 18477 12540 18541 12544
rect 18477 12484 18481 12540
rect 18481 12484 18537 12540
rect 18537 12484 18541 12540
rect 18477 12480 18541 12484
rect 18557 12540 18621 12544
rect 18557 12484 18561 12540
rect 18561 12484 18617 12540
rect 18617 12484 18621 12540
rect 18557 12480 18621 12484
rect 25263 12540 25327 12544
rect 25263 12484 25267 12540
rect 25267 12484 25323 12540
rect 25323 12484 25327 12540
rect 25263 12480 25327 12484
rect 25343 12540 25407 12544
rect 25343 12484 25347 12540
rect 25347 12484 25403 12540
rect 25403 12484 25407 12540
rect 25343 12480 25407 12484
rect 25423 12540 25487 12544
rect 25423 12484 25427 12540
rect 25427 12484 25483 12540
rect 25483 12484 25487 12540
rect 25423 12480 25487 12484
rect 25503 12540 25567 12544
rect 25503 12484 25507 12540
rect 25507 12484 25563 12540
rect 25563 12484 25567 12540
rect 25503 12480 25567 12484
rect 7898 11996 7962 12000
rect 7898 11940 7902 11996
rect 7902 11940 7958 11996
rect 7958 11940 7962 11996
rect 7898 11936 7962 11940
rect 7978 11996 8042 12000
rect 7978 11940 7982 11996
rect 7982 11940 8038 11996
rect 8038 11940 8042 11996
rect 7978 11936 8042 11940
rect 8058 11996 8122 12000
rect 8058 11940 8062 11996
rect 8062 11940 8118 11996
rect 8118 11940 8122 11996
rect 8058 11936 8122 11940
rect 8138 11996 8202 12000
rect 8138 11940 8142 11996
rect 8142 11940 8198 11996
rect 8198 11940 8202 11996
rect 8138 11936 8202 11940
rect 14844 11996 14908 12000
rect 14844 11940 14848 11996
rect 14848 11940 14904 11996
rect 14904 11940 14908 11996
rect 14844 11936 14908 11940
rect 14924 11996 14988 12000
rect 14924 11940 14928 11996
rect 14928 11940 14984 11996
rect 14984 11940 14988 11996
rect 14924 11936 14988 11940
rect 15004 11996 15068 12000
rect 15004 11940 15008 11996
rect 15008 11940 15064 11996
rect 15064 11940 15068 11996
rect 15004 11936 15068 11940
rect 15084 11996 15148 12000
rect 15084 11940 15088 11996
rect 15088 11940 15144 11996
rect 15144 11940 15148 11996
rect 15084 11936 15148 11940
rect 21790 11996 21854 12000
rect 21790 11940 21794 11996
rect 21794 11940 21850 11996
rect 21850 11940 21854 11996
rect 21790 11936 21854 11940
rect 21870 11996 21934 12000
rect 21870 11940 21874 11996
rect 21874 11940 21930 11996
rect 21930 11940 21934 11996
rect 21870 11936 21934 11940
rect 21950 11996 22014 12000
rect 21950 11940 21954 11996
rect 21954 11940 22010 11996
rect 22010 11940 22014 11996
rect 21950 11936 22014 11940
rect 22030 11996 22094 12000
rect 22030 11940 22034 11996
rect 22034 11940 22090 11996
rect 22090 11940 22094 11996
rect 22030 11936 22094 11940
rect 28736 11996 28800 12000
rect 28736 11940 28740 11996
rect 28740 11940 28796 11996
rect 28796 11940 28800 11996
rect 28736 11936 28800 11940
rect 28816 11996 28880 12000
rect 28816 11940 28820 11996
rect 28820 11940 28876 11996
rect 28876 11940 28880 11996
rect 28816 11936 28880 11940
rect 28896 11996 28960 12000
rect 28896 11940 28900 11996
rect 28900 11940 28956 11996
rect 28956 11940 28960 11996
rect 28896 11936 28960 11940
rect 28976 11996 29040 12000
rect 28976 11940 28980 11996
rect 28980 11940 29036 11996
rect 29036 11940 29040 11996
rect 28976 11936 29040 11940
rect 18828 11928 18892 11932
rect 18828 11872 18878 11928
rect 18878 11872 18892 11928
rect 18828 11868 18892 11872
rect 4425 11452 4489 11456
rect 4425 11396 4429 11452
rect 4429 11396 4485 11452
rect 4485 11396 4489 11452
rect 4425 11392 4489 11396
rect 4505 11452 4569 11456
rect 4505 11396 4509 11452
rect 4509 11396 4565 11452
rect 4565 11396 4569 11452
rect 4505 11392 4569 11396
rect 4585 11452 4649 11456
rect 4585 11396 4589 11452
rect 4589 11396 4645 11452
rect 4645 11396 4649 11452
rect 4585 11392 4649 11396
rect 4665 11452 4729 11456
rect 4665 11396 4669 11452
rect 4669 11396 4725 11452
rect 4725 11396 4729 11452
rect 4665 11392 4729 11396
rect 11371 11452 11435 11456
rect 11371 11396 11375 11452
rect 11375 11396 11431 11452
rect 11431 11396 11435 11452
rect 11371 11392 11435 11396
rect 11451 11452 11515 11456
rect 11451 11396 11455 11452
rect 11455 11396 11511 11452
rect 11511 11396 11515 11452
rect 11451 11392 11515 11396
rect 11531 11452 11595 11456
rect 11531 11396 11535 11452
rect 11535 11396 11591 11452
rect 11591 11396 11595 11452
rect 11531 11392 11595 11396
rect 11611 11452 11675 11456
rect 11611 11396 11615 11452
rect 11615 11396 11671 11452
rect 11671 11396 11675 11452
rect 11611 11392 11675 11396
rect 18317 11452 18381 11456
rect 18317 11396 18321 11452
rect 18321 11396 18377 11452
rect 18377 11396 18381 11452
rect 18317 11392 18381 11396
rect 18397 11452 18461 11456
rect 18397 11396 18401 11452
rect 18401 11396 18457 11452
rect 18457 11396 18461 11452
rect 18397 11392 18461 11396
rect 18477 11452 18541 11456
rect 18477 11396 18481 11452
rect 18481 11396 18537 11452
rect 18537 11396 18541 11452
rect 18477 11392 18541 11396
rect 18557 11452 18621 11456
rect 18557 11396 18561 11452
rect 18561 11396 18617 11452
rect 18617 11396 18621 11452
rect 18557 11392 18621 11396
rect 25263 11452 25327 11456
rect 25263 11396 25267 11452
rect 25267 11396 25323 11452
rect 25323 11396 25327 11452
rect 25263 11392 25327 11396
rect 25343 11452 25407 11456
rect 25343 11396 25347 11452
rect 25347 11396 25403 11452
rect 25403 11396 25407 11452
rect 25343 11392 25407 11396
rect 25423 11452 25487 11456
rect 25423 11396 25427 11452
rect 25427 11396 25483 11452
rect 25483 11396 25487 11452
rect 25423 11392 25487 11396
rect 25503 11452 25567 11456
rect 25503 11396 25507 11452
rect 25507 11396 25563 11452
rect 25563 11396 25567 11452
rect 25503 11392 25567 11396
rect 7898 10908 7962 10912
rect 7898 10852 7902 10908
rect 7902 10852 7958 10908
rect 7958 10852 7962 10908
rect 7898 10848 7962 10852
rect 7978 10908 8042 10912
rect 7978 10852 7982 10908
rect 7982 10852 8038 10908
rect 8038 10852 8042 10908
rect 7978 10848 8042 10852
rect 8058 10908 8122 10912
rect 8058 10852 8062 10908
rect 8062 10852 8118 10908
rect 8118 10852 8122 10908
rect 8058 10848 8122 10852
rect 8138 10908 8202 10912
rect 8138 10852 8142 10908
rect 8142 10852 8198 10908
rect 8198 10852 8202 10908
rect 8138 10848 8202 10852
rect 14844 10908 14908 10912
rect 14844 10852 14848 10908
rect 14848 10852 14904 10908
rect 14904 10852 14908 10908
rect 14844 10848 14908 10852
rect 14924 10908 14988 10912
rect 14924 10852 14928 10908
rect 14928 10852 14984 10908
rect 14984 10852 14988 10908
rect 14924 10848 14988 10852
rect 15004 10908 15068 10912
rect 15004 10852 15008 10908
rect 15008 10852 15064 10908
rect 15064 10852 15068 10908
rect 15004 10848 15068 10852
rect 15084 10908 15148 10912
rect 15084 10852 15088 10908
rect 15088 10852 15144 10908
rect 15144 10852 15148 10908
rect 15084 10848 15148 10852
rect 21790 10908 21854 10912
rect 21790 10852 21794 10908
rect 21794 10852 21850 10908
rect 21850 10852 21854 10908
rect 21790 10848 21854 10852
rect 21870 10908 21934 10912
rect 21870 10852 21874 10908
rect 21874 10852 21930 10908
rect 21930 10852 21934 10908
rect 21870 10848 21934 10852
rect 21950 10908 22014 10912
rect 21950 10852 21954 10908
rect 21954 10852 22010 10908
rect 22010 10852 22014 10908
rect 21950 10848 22014 10852
rect 22030 10908 22094 10912
rect 22030 10852 22034 10908
rect 22034 10852 22090 10908
rect 22090 10852 22094 10908
rect 22030 10848 22094 10852
rect 28736 10908 28800 10912
rect 28736 10852 28740 10908
rect 28740 10852 28796 10908
rect 28796 10852 28800 10908
rect 28736 10848 28800 10852
rect 28816 10908 28880 10912
rect 28816 10852 28820 10908
rect 28820 10852 28876 10908
rect 28876 10852 28880 10908
rect 28816 10848 28880 10852
rect 28896 10908 28960 10912
rect 28896 10852 28900 10908
rect 28900 10852 28956 10908
rect 28956 10852 28960 10908
rect 28896 10848 28960 10852
rect 28976 10908 29040 10912
rect 28976 10852 28980 10908
rect 28980 10852 29036 10908
rect 29036 10852 29040 10908
rect 28976 10848 29040 10852
rect 4425 10364 4489 10368
rect 4425 10308 4429 10364
rect 4429 10308 4485 10364
rect 4485 10308 4489 10364
rect 4425 10304 4489 10308
rect 4505 10364 4569 10368
rect 4505 10308 4509 10364
rect 4509 10308 4565 10364
rect 4565 10308 4569 10364
rect 4505 10304 4569 10308
rect 4585 10364 4649 10368
rect 4585 10308 4589 10364
rect 4589 10308 4645 10364
rect 4645 10308 4649 10364
rect 4585 10304 4649 10308
rect 4665 10364 4729 10368
rect 4665 10308 4669 10364
rect 4669 10308 4725 10364
rect 4725 10308 4729 10364
rect 4665 10304 4729 10308
rect 11371 10364 11435 10368
rect 11371 10308 11375 10364
rect 11375 10308 11431 10364
rect 11431 10308 11435 10364
rect 11371 10304 11435 10308
rect 11451 10364 11515 10368
rect 11451 10308 11455 10364
rect 11455 10308 11511 10364
rect 11511 10308 11515 10364
rect 11451 10304 11515 10308
rect 11531 10364 11595 10368
rect 11531 10308 11535 10364
rect 11535 10308 11591 10364
rect 11591 10308 11595 10364
rect 11531 10304 11595 10308
rect 11611 10364 11675 10368
rect 11611 10308 11615 10364
rect 11615 10308 11671 10364
rect 11671 10308 11675 10364
rect 11611 10304 11675 10308
rect 18317 10364 18381 10368
rect 18317 10308 18321 10364
rect 18321 10308 18377 10364
rect 18377 10308 18381 10364
rect 18317 10304 18381 10308
rect 18397 10364 18461 10368
rect 18397 10308 18401 10364
rect 18401 10308 18457 10364
rect 18457 10308 18461 10364
rect 18397 10304 18461 10308
rect 18477 10364 18541 10368
rect 18477 10308 18481 10364
rect 18481 10308 18537 10364
rect 18537 10308 18541 10364
rect 18477 10304 18541 10308
rect 18557 10364 18621 10368
rect 18557 10308 18561 10364
rect 18561 10308 18617 10364
rect 18617 10308 18621 10364
rect 18557 10304 18621 10308
rect 25263 10364 25327 10368
rect 25263 10308 25267 10364
rect 25267 10308 25323 10364
rect 25323 10308 25327 10364
rect 25263 10304 25327 10308
rect 25343 10364 25407 10368
rect 25343 10308 25347 10364
rect 25347 10308 25403 10364
rect 25403 10308 25407 10364
rect 25343 10304 25407 10308
rect 25423 10364 25487 10368
rect 25423 10308 25427 10364
rect 25427 10308 25483 10364
rect 25483 10308 25487 10364
rect 25423 10304 25487 10308
rect 25503 10364 25567 10368
rect 25503 10308 25507 10364
rect 25507 10308 25563 10364
rect 25563 10308 25567 10364
rect 25503 10304 25567 10308
rect 7898 9820 7962 9824
rect 7898 9764 7902 9820
rect 7902 9764 7958 9820
rect 7958 9764 7962 9820
rect 7898 9760 7962 9764
rect 7978 9820 8042 9824
rect 7978 9764 7982 9820
rect 7982 9764 8038 9820
rect 8038 9764 8042 9820
rect 7978 9760 8042 9764
rect 8058 9820 8122 9824
rect 8058 9764 8062 9820
rect 8062 9764 8118 9820
rect 8118 9764 8122 9820
rect 8058 9760 8122 9764
rect 8138 9820 8202 9824
rect 8138 9764 8142 9820
rect 8142 9764 8198 9820
rect 8198 9764 8202 9820
rect 8138 9760 8202 9764
rect 14844 9820 14908 9824
rect 14844 9764 14848 9820
rect 14848 9764 14904 9820
rect 14904 9764 14908 9820
rect 14844 9760 14908 9764
rect 14924 9820 14988 9824
rect 14924 9764 14928 9820
rect 14928 9764 14984 9820
rect 14984 9764 14988 9820
rect 14924 9760 14988 9764
rect 15004 9820 15068 9824
rect 15004 9764 15008 9820
rect 15008 9764 15064 9820
rect 15064 9764 15068 9820
rect 15004 9760 15068 9764
rect 15084 9820 15148 9824
rect 15084 9764 15088 9820
rect 15088 9764 15144 9820
rect 15144 9764 15148 9820
rect 15084 9760 15148 9764
rect 21790 9820 21854 9824
rect 21790 9764 21794 9820
rect 21794 9764 21850 9820
rect 21850 9764 21854 9820
rect 21790 9760 21854 9764
rect 21870 9820 21934 9824
rect 21870 9764 21874 9820
rect 21874 9764 21930 9820
rect 21930 9764 21934 9820
rect 21870 9760 21934 9764
rect 21950 9820 22014 9824
rect 21950 9764 21954 9820
rect 21954 9764 22010 9820
rect 22010 9764 22014 9820
rect 21950 9760 22014 9764
rect 22030 9820 22094 9824
rect 22030 9764 22034 9820
rect 22034 9764 22090 9820
rect 22090 9764 22094 9820
rect 22030 9760 22094 9764
rect 28736 9820 28800 9824
rect 28736 9764 28740 9820
rect 28740 9764 28796 9820
rect 28796 9764 28800 9820
rect 28736 9760 28800 9764
rect 28816 9820 28880 9824
rect 28816 9764 28820 9820
rect 28820 9764 28876 9820
rect 28876 9764 28880 9820
rect 28816 9760 28880 9764
rect 28896 9820 28960 9824
rect 28896 9764 28900 9820
rect 28900 9764 28956 9820
rect 28956 9764 28960 9820
rect 28896 9760 28960 9764
rect 28976 9820 29040 9824
rect 28976 9764 28980 9820
rect 28980 9764 29036 9820
rect 29036 9764 29040 9820
rect 28976 9760 29040 9764
rect 4425 9276 4489 9280
rect 4425 9220 4429 9276
rect 4429 9220 4485 9276
rect 4485 9220 4489 9276
rect 4425 9216 4489 9220
rect 4505 9276 4569 9280
rect 4505 9220 4509 9276
rect 4509 9220 4565 9276
rect 4565 9220 4569 9276
rect 4505 9216 4569 9220
rect 4585 9276 4649 9280
rect 4585 9220 4589 9276
rect 4589 9220 4645 9276
rect 4645 9220 4649 9276
rect 4585 9216 4649 9220
rect 4665 9276 4729 9280
rect 4665 9220 4669 9276
rect 4669 9220 4725 9276
rect 4725 9220 4729 9276
rect 4665 9216 4729 9220
rect 11371 9276 11435 9280
rect 11371 9220 11375 9276
rect 11375 9220 11431 9276
rect 11431 9220 11435 9276
rect 11371 9216 11435 9220
rect 11451 9276 11515 9280
rect 11451 9220 11455 9276
rect 11455 9220 11511 9276
rect 11511 9220 11515 9276
rect 11451 9216 11515 9220
rect 11531 9276 11595 9280
rect 11531 9220 11535 9276
rect 11535 9220 11591 9276
rect 11591 9220 11595 9276
rect 11531 9216 11595 9220
rect 11611 9276 11675 9280
rect 11611 9220 11615 9276
rect 11615 9220 11671 9276
rect 11671 9220 11675 9276
rect 11611 9216 11675 9220
rect 18317 9276 18381 9280
rect 18317 9220 18321 9276
rect 18321 9220 18377 9276
rect 18377 9220 18381 9276
rect 18317 9216 18381 9220
rect 18397 9276 18461 9280
rect 18397 9220 18401 9276
rect 18401 9220 18457 9276
rect 18457 9220 18461 9276
rect 18397 9216 18461 9220
rect 18477 9276 18541 9280
rect 18477 9220 18481 9276
rect 18481 9220 18537 9276
rect 18537 9220 18541 9276
rect 18477 9216 18541 9220
rect 18557 9276 18621 9280
rect 18557 9220 18561 9276
rect 18561 9220 18617 9276
rect 18617 9220 18621 9276
rect 18557 9216 18621 9220
rect 25263 9276 25327 9280
rect 25263 9220 25267 9276
rect 25267 9220 25323 9276
rect 25323 9220 25327 9276
rect 25263 9216 25327 9220
rect 25343 9276 25407 9280
rect 25343 9220 25347 9276
rect 25347 9220 25403 9276
rect 25403 9220 25407 9276
rect 25343 9216 25407 9220
rect 25423 9276 25487 9280
rect 25423 9220 25427 9276
rect 25427 9220 25483 9276
rect 25483 9220 25487 9276
rect 25423 9216 25487 9220
rect 25503 9276 25567 9280
rect 25503 9220 25507 9276
rect 25507 9220 25563 9276
rect 25563 9220 25567 9276
rect 25503 9216 25567 9220
rect 7898 8732 7962 8736
rect 7898 8676 7902 8732
rect 7902 8676 7958 8732
rect 7958 8676 7962 8732
rect 7898 8672 7962 8676
rect 7978 8732 8042 8736
rect 7978 8676 7982 8732
rect 7982 8676 8038 8732
rect 8038 8676 8042 8732
rect 7978 8672 8042 8676
rect 8058 8732 8122 8736
rect 8058 8676 8062 8732
rect 8062 8676 8118 8732
rect 8118 8676 8122 8732
rect 8058 8672 8122 8676
rect 8138 8732 8202 8736
rect 8138 8676 8142 8732
rect 8142 8676 8198 8732
rect 8198 8676 8202 8732
rect 8138 8672 8202 8676
rect 14844 8732 14908 8736
rect 14844 8676 14848 8732
rect 14848 8676 14904 8732
rect 14904 8676 14908 8732
rect 14844 8672 14908 8676
rect 14924 8732 14988 8736
rect 14924 8676 14928 8732
rect 14928 8676 14984 8732
rect 14984 8676 14988 8732
rect 14924 8672 14988 8676
rect 15004 8732 15068 8736
rect 15004 8676 15008 8732
rect 15008 8676 15064 8732
rect 15064 8676 15068 8732
rect 15004 8672 15068 8676
rect 15084 8732 15148 8736
rect 15084 8676 15088 8732
rect 15088 8676 15144 8732
rect 15144 8676 15148 8732
rect 15084 8672 15148 8676
rect 21790 8732 21854 8736
rect 21790 8676 21794 8732
rect 21794 8676 21850 8732
rect 21850 8676 21854 8732
rect 21790 8672 21854 8676
rect 21870 8732 21934 8736
rect 21870 8676 21874 8732
rect 21874 8676 21930 8732
rect 21930 8676 21934 8732
rect 21870 8672 21934 8676
rect 21950 8732 22014 8736
rect 21950 8676 21954 8732
rect 21954 8676 22010 8732
rect 22010 8676 22014 8732
rect 21950 8672 22014 8676
rect 22030 8732 22094 8736
rect 22030 8676 22034 8732
rect 22034 8676 22090 8732
rect 22090 8676 22094 8732
rect 22030 8672 22094 8676
rect 28736 8732 28800 8736
rect 28736 8676 28740 8732
rect 28740 8676 28796 8732
rect 28796 8676 28800 8732
rect 28736 8672 28800 8676
rect 28816 8732 28880 8736
rect 28816 8676 28820 8732
rect 28820 8676 28876 8732
rect 28876 8676 28880 8732
rect 28816 8672 28880 8676
rect 28896 8732 28960 8736
rect 28896 8676 28900 8732
rect 28900 8676 28956 8732
rect 28956 8676 28960 8732
rect 28896 8672 28960 8676
rect 28976 8732 29040 8736
rect 28976 8676 28980 8732
rect 28980 8676 29036 8732
rect 29036 8676 29040 8732
rect 28976 8672 29040 8676
rect 4425 8188 4489 8192
rect 4425 8132 4429 8188
rect 4429 8132 4485 8188
rect 4485 8132 4489 8188
rect 4425 8128 4489 8132
rect 4505 8188 4569 8192
rect 4505 8132 4509 8188
rect 4509 8132 4565 8188
rect 4565 8132 4569 8188
rect 4505 8128 4569 8132
rect 4585 8188 4649 8192
rect 4585 8132 4589 8188
rect 4589 8132 4645 8188
rect 4645 8132 4649 8188
rect 4585 8128 4649 8132
rect 4665 8188 4729 8192
rect 4665 8132 4669 8188
rect 4669 8132 4725 8188
rect 4725 8132 4729 8188
rect 4665 8128 4729 8132
rect 11371 8188 11435 8192
rect 11371 8132 11375 8188
rect 11375 8132 11431 8188
rect 11431 8132 11435 8188
rect 11371 8128 11435 8132
rect 11451 8188 11515 8192
rect 11451 8132 11455 8188
rect 11455 8132 11511 8188
rect 11511 8132 11515 8188
rect 11451 8128 11515 8132
rect 11531 8188 11595 8192
rect 11531 8132 11535 8188
rect 11535 8132 11591 8188
rect 11591 8132 11595 8188
rect 11531 8128 11595 8132
rect 11611 8188 11675 8192
rect 11611 8132 11615 8188
rect 11615 8132 11671 8188
rect 11671 8132 11675 8188
rect 11611 8128 11675 8132
rect 18317 8188 18381 8192
rect 18317 8132 18321 8188
rect 18321 8132 18377 8188
rect 18377 8132 18381 8188
rect 18317 8128 18381 8132
rect 18397 8188 18461 8192
rect 18397 8132 18401 8188
rect 18401 8132 18457 8188
rect 18457 8132 18461 8188
rect 18397 8128 18461 8132
rect 18477 8188 18541 8192
rect 18477 8132 18481 8188
rect 18481 8132 18537 8188
rect 18537 8132 18541 8188
rect 18477 8128 18541 8132
rect 18557 8188 18621 8192
rect 18557 8132 18561 8188
rect 18561 8132 18617 8188
rect 18617 8132 18621 8188
rect 18557 8128 18621 8132
rect 25263 8188 25327 8192
rect 25263 8132 25267 8188
rect 25267 8132 25323 8188
rect 25323 8132 25327 8188
rect 25263 8128 25327 8132
rect 25343 8188 25407 8192
rect 25343 8132 25347 8188
rect 25347 8132 25403 8188
rect 25403 8132 25407 8188
rect 25343 8128 25407 8132
rect 25423 8188 25487 8192
rect 25423 8132 25427 8188
rect 25427 8132 25483 8188
rect 25483 8132 25487 8188
rect 25423 8128 25487 8132
rect 25503 8188 25567 8192
rect 25503 8132 25507 8188
rect 25507 8132 25563 8188
rect 25563 8132 25567 8188
rect 25503 8128 25567 8132
rect 7898 7644 7962 7648
rect 7898 7588 7902 7644
rect 7902 7588 7958 7644
rect 7958 7588 7962 7644
rect 7898 7584 7962 7588
rect 7978 7644 8042 7648
rect 7978 7588 7982 7644
rect 7982 7588 8038 7644
rect 8038 7588 8042 7644
rect 7978 7584 8042 7588
rect 8058 7644 8122 7648
rect 8058 7588 8062 7644
rect 8062 7588 8118 7644
rect 8118 7588 8122 7644
rect 8058 7584 8122 7588
rect 8138 7644 8202 7648
rect 8138 7588 8142 7644
rect 8142 7588 8198 7644
rect 8198 7588 8202 7644
rect 8138 7584 8202 7588
rect 14844 7644 14908 7648
rect 14844 7588 14848 7644
rect 14848 7588 14904 7644
rect 14904 7588 14908 7644
rect 14844 7584 14908 7588
rect 14924 7644 14988 7648
rect 14924 7588 14928 7644
rect 14928 7588 14984 7644
rect 14984 7588 14988 7644
rect 14924 7584 14988 7588
rect 15004 7644 15068 7648
rect 15004 7588 15008 7644
rect 15008 7588 15064 7644
rect 15064 7588 15068 7644
rect 15004 7584 15068 7588
rect 15084 7644 15148 7648
rect 15084 7588 15088 7644
rect 15088 7588 15144 7644
rect 15144 7588 15148 7644
rect 15084 7584 15148 7588
rect 21790 7644 21854 7648
rect 21790 7588 21794 7644
rect 21794 7588 21850 7644
rect 21850 7588 21854 7644
rect 21790 7584 21854 7588
rect 21870 7644 21934 7648
rect 21870 7588 21874 7644
rect 21874 7588 21930 7644
rect 21930 7588 21934 7644
rect 21870 7584 21934 7588
rect 21950 7644 22014 7648
rect 21950 7588 21954 7644
rect 21954 7588 22010 7644
rect 22010 7588 22014 7644
rect 21950 7584 22014 7588
rect 22030 7644 22094 7648
rect 22030 7588 22034 7644
rect 22034 7588 22090 7644
rect 22090 7588 22094 7644
rect 22030 7584 22094 7588
rect 28736 7644 28800 7648
rect 28736 7588 28740 7644
rect 28740 7588 28796 7644
rect 28796 7588 28800 7644
rect 28736 7584 28800 7588
rect 28816 7644 28880 7648
rect 28816 7588 28820 7644
rect 28820 7588 28876 7644
rect 28876 7588 28880 7644
rect 28816 7584 28880 7588
rect 28896 7644 28960 7648
rect 28896 7588 28900 7644
rect 28900 7588 28956 7644
rect 28956 7588 28960 7644
rect 28896 7584 28960 7588
rect 28976 7644 29040 7648
rect 28976 7588 28980 7644
rect 28980 7588 29036 7644
rect 29036 7588 29040 7644
rect 28976 7584 29040 7588
rect 4425 7100 4489 7104
rect 4425 7044 4429 7100
rect 4429 7044 4485 7100
rect 4485 7044 4489 7100
rect 4425 7040 4489 7044
rect 4505 7100 4569 7104
rect 4505 7044 4509 7100
rect 4509 7044 4565 7100
rect 4565 7044 4569 7100
rect 4505 7040 4569 7044
rect 4585 7100 4649 7104
rect 4585 7044 4589 7100
rect 4589 7044 4645 7100
rect 4645 7044 4649 7100
rect 4585 7040 4649 7044
rect 4665 7100 4729 7104
rect 4665 7044 4669 7100
rect 4669 7044 4725 7100
rect 4725 7044 4729 7100
rect 4665 7040 4729 7044
rect 11371 7100 11435 7104
rect 11371 7044 11375 7100
rect 11375 7044 11431 7100
rect 11431 7044 11435 7100
rect 11371 7040 11435 7044
rect 11451 7100 11515 7104
rect 11451 7044 11455 7100
rect 11455 7044 11511 7100
rect 11511 7044 11515 7100
rect 11451 7040 11515 7044
rect 11531 7100 11595 7104
rect 11531 7044 11535 7100
rect 11535 7044 11591 7100
rect 11591 7044 11595 7100
rect 11531 7040 11595 7044
rect 11611 7100 11675 7104
rect 11611 7044 11615 7100
rect 11615 7044 11671 7100
rect 11671 7044 11675 7100
rect 11611 7040 11675 7044
rect 18317 7100 18381 7104
rect 18317 7044 18321 7100
rect 18321 7044 18377 7100
rect 18377 7044 18381 7100
rect 18317 7040 18381 7044
rect 18397 7100 18461 7104
rect 18397 7044 18401 7100
rect 18401 7044 18457 7100
rect 18457 7044 18461 7100
rect 18397 7040 18461 7044
rect 18477 7100 18541 7104
rect 18477 7044 18481 7100
rect 18481 7044 18537 7100
rect 18537 7044 18541 7100
rect 18477 7040 18541 7044
rect 18557 7100 18621 7104
rect 18557 7044 18561 7100
rect 18561 7044 18617 7100
rect 18617 7044 18621 7100
rect 18557 7040 18621 7044
rect 25263 7100 25327 7104
rect 25263 7044 25267 7100
rect 25267 7044 25323 7100
rect 25323 7044 25327 7100
rect 25263 7040 25327 7044
rect 25343 7100 25407 7104
rect 25343 7044 25347 7100
rect 25347 7044 25403 7100
rect 25403 7044 25407 7100
rect 25343 7040 25407 7044
rect 25423 7100 25487 7104
rect 25423 7044 25427 7100
rect 25427 7044 25483 7100
rect 25483 7044 25487 7100
rect 25423 7040 25487 7044
rect 25503 7100 25567 7104
rect 25503 7044 25507 7100
rect 25507 7044 25563 7100
rect 25563 7044 25567 7100
rect 25503 7040 25567 7044
rect 7898 6556 7962 6560
rect 7898 6500 7902 6556
rect 7902 6500 7958 6556
rect 7958 6500 7962 6556
rect 7898 6496 7962 6500
rect 7978 6556 8042 6560
rect 7978 6500 7982 6556
rect 7982 6500 8038 6556
rect 8038 6500 8042 6556
rect 7978 6496 8042 6500
rect 8058 6556 8122 6560
rect 8058 6500 8062 6556
rect 8062 6500 8118 6556
rect 8118 6500 8122 6556
rect 8058 6496 8122 6500
rect 8138 6556 8202 6560
rect 8138 6500 8142 6556
rect 8142 6500 8198 6556
rect 8198 6500 8202 6556
rect 8138 6496 8202 6500
rect 14844 6556 14908 6560
rect 14844 6500 14848 6556
rect 14848 6500 14904 6556
rect 14904 6500 14908 6556
rect 14844 6496 14908 6500
rect 14924 6556 14988 6560
rect 14924 6500 14928 6556
rect 14928 6500 14984 6556
rect 14984 6500 14988 6556
rect 14924 6496 14988 6500
rect 15004 6556 15068 6560
rect 15004 6500 15008 6556
rect 15008 6500 15064 6556
rect 15064 6500 15068 6556
rect 15004 6496 15068 6500
rect 15084 6556 15148 6560
rect 15084 6500 15088 6556
rect 15088 6500 15144 6556
rect 15144 6500 15148 6556
rect 15084 6496 15148 6500
rect 21790 6556 21854 6560
rect 21790 6500 21794 6556
rect 21794 6500 21850 6556
rect 21850 6500 21854 6556
rect 21790 6496 21854 6500
rect 21870 6556 21934 6560
rect 21870 6500 21874 6556
rect 21874 6500 21930 6556
rect 21930 6500 21934 6556
rect 21870 6496 21934 6500
rect 21950 6556 22014 6560
rect 21950 6500 21954 6556
rect 21954 6500 22010 6556
rect 22010 6500 22014 6556
rect 21950 6496 22014 6500
rect 22030 6556 22094 6560
rect 22030 6500 22034 6556
rect 22034 6500 22090 6556
rect 22090 6500 22094 6556
rect 22030 6496 22094 6500
rect 28736 6556 28800 6560
rect 28736 6500 28740 6556
rect 28740 6500 28796 6556
rect 28796 6500 28800 6556
rect 28736 6496 28800 6500
rect 28816 6556 28880 6560
rect 28816 6500 28820 6556
rect 28820 6500 28876 6556
rect 28876 6500 28880 6556
rect 28816 6496 28880 6500
rect 28896 6556 28960 6560
rect 28896 6500 28900 6556
rect 28900 6500 28956 6556
rect 28956 6500 28960 6556
rect 28896 6496 28960 6500
rect 28976 6556 29040 6560
rect 28976 6500 28980 6556
rect 28980 6500 29036 6556
rect 29036 6500 29040 6556
rect 28976 6496 29040 6500
rect 4425 6012 4489 6016
rect 4425 5956 4429 6012
rect 4429 5956 4485 6012
rect 4485 5956 4489 6012
rect 4425 5952 4489 5956
rect 4505 6012 4569 6016
rect 4505 5956 4509 6012
rect 4509 5956 4565 6012
rect 4565 5956 4569 6012
rect 4505 5952 4569 5956
rect 4585 6012 4649 6016
rect 4585 5956 4589 6012
rect 4589 5956 4645 6012
rect 4645 5956 4649 6012
rect 4585 5952 4649 5956
rect 4665 6012 4729 6016
rect 4665 5956 4669 6012
rect 4669 5956 4725 6012
rect 4725 5956 4729 6012
rect 4665 5952 4729 5956
rect 11371 6012 11435 6016
rect 11371 5956 11375 6012
rect 11375 5956 11431 6012
rect 11431 5956 11435 6012
rect 11371 5952 11435 5956
rect 11451 6012 11515 6016
rect 11451 5956 11455 6012
rect 11455 5956 11511 6012
rect 11511 5956 11515 6012
rect 11451 5952 11515 5956
rect 11531 6012 11595 6016
rect 11531 5956 11535 6012
rect 11535 5956 11591 6012
rect 11591 5956 11595 6012
rect 11531 5952 11595 5956
rect 11611 6012 11675 6016
rect 11611 5956 11615 6012
rect 11615 5956 11671 6012
rect 11671 5956 11675 6012
rect 11611 5952 11675 5956
rect 18317 6012 18381 6016
rect 18317 5956 18321 6012
rect 18321 5956 18377 6012
rect 18377 5956 18381 6012
rect 18317 5952 18381 5956
rect 18397 6012 18461 6016
rect 18397 5956 18401 6012
rect 18401 5956 18457 6012
rect 18457 5956 18461 6012
rect 18397 5952 18461 5956
rect 18477 6012 18541 6016
rect 18477 5956 18481 6012
rect 18481 5956 18537 6012
rect 18537 5956 18541 6012
rect 18477 5952 18541 5956
rect 18557 6012 18621 6016
rect 18557 5956 18561 6012
rect 18561 5956 18617 6012
rect 18617 5956 18621 6012
rect 18557 5952 18621 5956
rect 25263 6012 25327 6016
rect 25263 5956 25267 6012
rect 25267 5956 25323 6012
rect 25323 5956 25327 6012
rect 25263 5952 25327 5956
rect 25343 6012 25407 6016
rect 25343 5956 25347 6012
rect 25347 5956 25403 6012
rect 25403 5956 25407 6012
rect 25343 5952 25407 5956
rect 25423 6012 25487 6016
rect 25423 5956 25427 6012
rect 25427 5956 25483 6012
rect 25483 5956 25487 6012
rect 25423 5952 25487 5956
rect 25503 6012 25567 6016
rect 25503 5956 25507 6012
rect 25507 5956 25563 6012
rect 25563 5956 25567 6012
rect 25503 5952 25567 5956
rect 7898 5468 7962 5472
rect 7898 5412 7902 5468
rect 7902 5412 7958 5468
rect 7958 5412 7962 5468
rect 7898 5408 7962 5412
rect 7978 5468 8042 5472
rect 7978 5412 7982 5468
rect 7982 5412 8038 5468
rect 8038 5412 8042 5468
rect 7978 5408 8042 5412
rect 8058 5468 8122 5472
rect 8058 5412 8062 5468
rect 8062 5412 8118 5468
rect 8118 5412 8122 5468
rect 8058 5408 8122 5412
rect 8138 5468 8202 5472
rect 8138 5412 8142 5468
rect 8142 5412 8198 5468
rect 8198 5412 8202 5468
rect 8138 5408 8202 5412
rect 14844 5468 14908 5472
rect 14844 5412 14848 5468
rect 14848 5412 14904 5468
rect 14904 5412 14908 5468
rect 14844 5408 14908 5412
rect 14924 5468 14988 5472
rect 14924 5412 14928 5468
rect 14928 5412 14984 5468
rect 14984 5412 14988 5468
rect 14924 5408 14988 5412
rect 15004 5468 15068 5472
rect 15004 5412 15008 5468
rect 15008 5412 15064 5468
rect 15064 5412 15068 5468
rect 15004 5408 15068 5412
rect 15084 5468 15148 5472
rect 15084 5412 15088 5468
rect 15088 5412 15144 5468
rect 15144 5412 15148 5468
rect 15084 5408 15148 5412
rect 21790 5468 21854 5472
rect 21790 5412 21794 5468
rect 21794 5412 21850 5468
rect 21850 5412 21854 5468
rect 21790 5408 21854 5412
rect 21870 5468 21934 5472
rect 21870 5412 21874 5468
rect 21874 5412 21930 5468
rect 21930 5412 21934 5468
rect 21870 5408 21934 5412
rect 21950 5468 22014 5472
rect 21950 5412 21954 5468
rect 21954 5412 22010 5468
rect 22010 5412 22014 5468
rect 21950 5408 22014 5412
rect 22030 5468 22094 5472
rect 22030 5412 22034 5468
rect 22034 5412 22090 5468
rect 22090 5412 22094 5468
rect 22030 5408 22094 5412
rect 28736 5468 28800 5472
rect 28736 5412 28740 5468
rect 28740 5412 28796 5468
rect 28796 5412 28800 5468
rect 28736 5408 28800 5412
rect 28816 5468 28880 5472
rect 28816 5412 28820 5468
rect 28820 5412 28876 5468
rect 28876 5412 28880 5468
rect 28816 5408 28880 5412
rect 28896 5468 28960 5472
rect 28896 5412 28900 5468
rect 28900 5412 28956 5468
rect 28956 5412 28960 5468
rect 28896 5408 28960 5412
rect 28976 5468 29040 5472
rect 28976 5412 28980 5468
rect 28980 5412 29036 5468
rect 29036 5412 29040 5468
rect 28976 5408 29040 5412
rect 4425 4924 4489 4928
rect 4425 4868 4429 4924
rect 4429 4868 4485 4924
rect 4485 4868 4489 4924
rect 4425 4864 4489 4868
rect 4505 4924 4569 4928
rect 4505 4868 4509 4924
rect 4509 4868 4565 4924
rect 4565 4868 4569 4924
rect 4505 4864 4569 4868
rect 4585 4924 4649 4928
rect 4585 4868 4589 4924
rect 4589 4868 4645 4924
rect 4645 4868 4649 4924
rect 4585 4864 4649 4868
rect 4665 4924 4729 4928
rect 4665 4868 4669 4924
rect 4669 4868 4725 4924
rect 4725 4868 4729 4924
rect 4665 4864 4729 4868
rect 11371 4924 11435 4928
rect 11371 4868 11375 4924
rect 11375 4868 11431 4924
rect 11431 4868 11435 4924
rect 11371 4864 11435 4868
rect 11451 4924 11515 4928
rect 11451 4868 11455 4924
rect 11455 4868 11511 4924
rect 11511 4868 11515 4924
rect 11451 4864 11515 4868
rect 11531 4924 11595 4928
rect 11531 4868 11535 4924
rect 11535 4868 11591 4924
rect 11591 4868 11595 4924
rect 11531 4864 11595 4868
rect 11611 4924 11675 4928
rect 11611 4868 11615 4924
rect 11615 4868 11671 4924
rect 11671 4868 11675 4924
rect 11611 4864 11675 4868
rect 18317 4924 18381 4928
rect 18317 4868 18321 4924
rect 18321 4868 18377 4924
rect 18377 4868 18381 4924
rect 18317 4864 18381 4868
rect 18397 4924 18461 4928
rect 18397 4868 18401 4924
rect 18401 4868 18457 4924
rect 18457 4868 18461 4924
rect 18397 4864 18461 4868
rect 18477 4924 18541 4928
rect 18477 4868 18481 4924
rect 18481 4868 18537 4924
rect 18537 4868 18541 4924
rect 18477 4864 18541 4868
rect 18557 4924 18621 4928
rect 18557 4868 18561 4924
rect 18561 4868 18617 4924
rect 18617 4868 18621 4924
rect 18557 4864 18621 4868
rect 25263 4924 25327 4928
rect 25263 4868 25267 4924
rect 25267 4868 25323 4924
rect 25323 4868 25327 4924
rect 25263 4864 25327 4868
rect 25343 4924 25407 4928
rect 25343 4868 25347 4924
rect 25347 4868 25403 4924
rect 25403 4868 25407 4924
rect 25343 4864 25407 4868
rect 25423 4924 25487 4928
rect 25423 4868 25427 4924
rect 25427 4868 25483 4924
rect 25483 4868 25487 4924
rect 25423 4864 25487 4868
rect 25503 4924 25567 4928
rect 25503 4868 25507 4924
rect 25507 4868 25563 4924
rect 25563 4868 25567 4924
rect 25503 4864 25567 4868
rect 7898 4380 7962 4384
rect 7898 4324 7902 4380
rect 7902 4324 7958 4380
rect 7958 4324 7962 4380
rect 7898 4320 7962 4324
rect 7978 4380 8042 4384
rect 7978 4324 7982 4380
rect 7982 4324 8038 4380
rect 8038 4324 8042 4380
rect 7978 4320 8042 4324
rect 8058 4380 8122 4384
rect 8058 4324 8062 4380
rect 8062 4324 8118 4380
rect 8118 4324 8122 4380
rect 8058 4320 8122 4324
rect 8138 4380 8202 4384
rect 8138 4324 8142 4380
rect 8142 4324 8198 4380
rect 8198 4324 8202 4380
rect 8138 4320 8202 4324
rect 14844 4380 14908 4384
rect 14844 4324 14848 4380
rect 14848 4324 14904 4380
rect 14904 4324 14908 4380
rect 14844 4320 14908 4324
rect 14924 4380 14988 4384
rect 14924 4324 14928 4380
rect 14928 4324 14984 4380
rect 14984 4324 14988 4380
rect 14924 4320 14988 4324
rect 15004 4380 15068 4384
rect 15004 4324 15008 4380
rect 15008 4324 15064 4380
rect 15064 4324 15068 4380
rect 15004 4320 15068 4324
rect 15084 4380 15148 4384
rect 15084 4324 15088 4380
rect 15088 4324 15144 4380
rect 15144 4324 15148 4380
rect 15084 4320 15148 4324
rect 21790 4380 21854 4384
rect 21790 4324 21794 4380
rect 21794 4324 21850 4380
rect 21850 4324 21854 4380
rect 21790 4320 21854 4324
rect 21870 4380 21934 4384
rect 21870 4324 21874 4380
rect 21874 4324 21930 4380
rect 21930 4324 21934 4380
rect 21870 4320 21934 4324
rect 21950 4380 22014 4384
rect 21950 4324 21954 4380
rect 21954 4324 22010 4380
rect 22010 4324 22014 4380
rect 21950 4320 22014 4324
rect 22030 4380 22094 4384
rect 22030 4324 22034 4380
rect 22034 4324 22090 4380
rect 22090 4324 22094 4380
rect 22030 4320 22094 4324
rect 28736 4380 28800 4384
rect 28736 4324 28740 4380
rect 28740 4324 28796 4380
rect 28796 4324 28800 4380
rect 28736 4320 28800 4324
rect 28816 4380 28880 4384
rect 28816 4324 28820 4380
rect 28820 4324 28876 4380
rect 28876 4324 28880 4380
rect 28816 4320 28880 4324
rect 28896 4380 28960 4384
rect 28896 4324 28900 4380
rect 28900 4324 28956 4380
rect 28956 4324 28960 4380
rect 28896 4320 28960 4324
rect 28976 4380 29040 4384
rect 28976 4324 28980 4380
rect 28980 4324 29036 4380
rect 29036 4324 29040 4380
rect 28976 4320 29040 4324
rect 4425 3836 4489 3840
rect 4425 3780 4429 3836
rect 4429 3780 4485 3836
rect 4485 3780 4489 3836
rect 4425 3776 4489 3780
rect 4505 3836 4569 3840
rect 4505 3780 4509 3836
rect 4509 3780 4565 3836
rect 4565 3780 4569 3836
rect 4505 3776 4569 3780
rect 4585 3836 4649 3840
rect 4585 3780 4589 3836
rect 4589 3780 4645 3836
rect 4645 3780 4649 3836
rect 4585 3776 4649 3780
rect 4665 3836 4729 3840
rect 4665 3780 4669 3836
rect 4669 3780 4725 3836
rect 4725 3780 4729 3836
rect 4665 3776 4729 3780
rect 11371 3836 11435 3840
rect 11371 3780 11375 3836
rect 11375 3780 11431 3836
rect 11431 3780 11435 3836
rect 11371 3776 11435 3780
rect 11451 3836 11515 3840
rect 11451 3780 11455 3836
rect 11455 3780 11511 3836
rect 11511 3780 11515 3836
rect 11451 3776 11515 3780
rect 11531 3836 11595 3840
rect 11531 3780 11535 3836
rect 11535 3780 11591 3836
rect 11591 3780 11595 3836
rect 11531 3776 11595 3780
rect 11611 3836 11675 3840
rect 11611 3780 11615 3836
rect 11615 3780 11671 3836
rect 11671 3780 11675 3836
rect 11611 3776 11675 3780
rect 18317 3836 18381 3840
rect 18317 3780 18321 3836
rect 18321 3780 18377 3836
rect 18377 3780 18381 3836
rect 18317 3776 18381 3780
rect 18397 3836 18461 3840
rect 18397 3780 18401 3836
rect 18401 3780 18457 3836
rect 18457 3780 18461 3836
rect 18397 3776 18461 3780
rect 18477 3836 18541 3840
rect 18477 3780 18481 3836
rect 18481 3780 18537 3836
rect 18537 3780 18541 3836
rect 18477 3776 18541 3780
rect 18557 3836 18621 3840
rect 18557 3780 18561 3836
rect 18561 3780 18617 3836
rect 18617 3780 18621 3836
rect 18557 3776 18621 3780
rect 25263 3836 25327 3840
rect 25263 3780 25267 3836
rect 25267 3780 25323 3836
rect 25323 3780 25327 3836
rect 25263 3776 25327 3780
rect 25343 3836 25407 3840
rect 25343 3780 25347 3836
rect 25347 3780 25403 3836
rect 25403 3780 25407 3836
rect 25343 3776 25407 3780
rect 25423 3836 25487 3840
rect 25423 3780 25427 3836
rect 25427 3780 25483 3836
rect 25483 3780 25487 3836
rect 25423 3776 25487 3780
rect 25503 3836 25567 3840
rect 25503 3780 25507 3836
rect 25507 3780 25563 3836
rect 25563 3780 25567 3836
rect 25503 3776 25567 3780
rect 7898 3292 7962 3296
rect 7898 3236 7902 3292
rect 7902 3236 7958 3292
rect 7958 3236 7962 3292
rect 7898 3232 7962 3236
rect 7978 3292 8042 3296
rect 7978 3236 7982 3292
rect 7982 3236 8038 3292
rect 8038 3236 8042 3292
rect 7978 3232 8042 3236
rect 8058 3292 8122 3296
rect 8058 3236 8062 3292
rect 8062 3236 8118 3292
rect 8118 3236 8122 3292
rect 8058 3232 8122 3236
rect 8138 3292 8202 3296
rect 8138 3236 8142 3292
rect 8142 3236 8198 3292
rect 8198 3236 8202 3292
rect 8138 3232 8202 3236
rect 14844 3292 14908 3296
rect 14844 3236 14848 3292
rect 14848 3236 14904 3292
rect 14904 3236 14908 3292
rect 14844 3232 14908 3236
rect 14924 3292 14988 3296
rect 14924 3236 14928 3292
rect 14928 3236 14984 3292
rect 14984 3236 14988 3292
rect 14924 3232 14988 3236
rect 15004 3292 15068 3296
rect 15004 3236 15008 3292
rect 15008 3236 15064 3292
rect 15064 3236 15068 3292
rect 15004 3232 15068 3236
rect 15084 3292 15148 3296
rect 15084 3236 15088 3292
rect 15088 3236 15144 3292
rect 15144 3236 15148 3292
rect 15084 3232 15148 3236
rect 21790 3292 21854 3296
rect 21790 3236 21794 3292
rect 21794 3236 21850 3292
rect 21850 3236 21854 3292
rect 21790 3232 21854 3236
rect 21870 3292 21934 3296
rect 21870 3236 21874 3292
rect 21874 3236 21930 3292
rect 21930 3236 21934 3292
rect 21870 3232 21934 3236
rect 21950 3292 22014 3296
rect 21950 3236 21954 3292
rect 21954 3236 22010 3292
rect 22010 3236 22014 3292
rect 21950 3232 22014 3236
rect 22030 3292 22094 3296
rect 22030 3236 22034 3292
rect 22034 3236 22090 3292
rect 22090 3236 22094 3292
rect 22030 3232 22094 3236
rect 28736 3292 28800 3296
rect 28736 3236 28740 3292
rect 28740 3236 28796 3292
rect 28796 3236 28800 3292
rect 28736 3232 28800 3236
rect 28816 3292 28880 3296
rect 28816 3236 28820 3292
rect 28820 3236 28876 3292
rect 28876 3236 28880 3292
rect 28816 3232 28880 3236
rect 28896 3292 28960 3296
rect 28896 3236 28900 3292
rect 28900 3236 28956 3292
rect 28956 3236 28960 3292
rect 28896 3232 28960 3236
rect 28976 3292 29040 3296
rect 28976 3236 28980 3292
rect 28980 3236 29036 3292
rect 29036 3236 29040 3292
rect 28976 3232 29040 3236
rect 4425 2748 4489 2752
rect 4425 2692 4429 2748
rect 4429 2692 4485 2748
rect 4485 2692 4489 2748
rect 4425 2688 4489 2692
rect 4505 2748 4569 2752
rect 4505 2692 4509 2748
rect 4509 2692 4565 2748
rect 4565 2692 4569 2748
rect 4505 2688 4569 2692
rect 4585 2748 4649 2752
rect 4585 2692 4589 2748
rect 4589 2692 4645 2748
rect 4645 2692 4649 2748
rect 4585 2688 4649 2692
rect 4665 2748 4729 2752
rect 4665 2692 4669 2748
rect 4669 2692 4725 2748
rect 4725 2692 4729 2748
rect 4665 2688 4729 2692
rect 11371 2748 11435 2752
rect 11371 2692 11375 2748
rect 11375 2692 11431 2748
rect 11431 2692 11435 2748
rect 11371 2688 11435 2692
rect 11451 2748 11515 2752
rect 11451 2692 11455 2748
rect 11455 2692 11511 2748
rect 11511 2692 11515 2748
rect 11451 2688 11515 2692
rect 11531 2748 11595 2752
rect 11531 2692 11535 2748
rect 11535 2692 11591 2748
rect 11591 2692 11595 2748
rect 11531 2688 11595 2692
rect 11611 2748 11675 2752
rect 11611 2692 11615 2748
rect 11615 2692 11671 2748
rect 11671 2692 11675 2748
rect 11611 2688 11675 2692
rect 18317 2748 18381 2752
rect 18317 2692 18321 2748
rect 18321 2692 18377 2748
rect 18377 2692 18381 2748
rect 18317 2688 18381 2692
rect 18397 2748 18461 2752
rect 18397 2692 18401 2748
rect 18401 2692 18457 2748
rect 18457 2692 18461 2748
rect 18397 2688 18461 2692
rect 18477 2748 18541 2752
rect 18477 2692 18481 2748
rect 18481 2692 18537 2748
rect 18537 2692 18541 2748
rect 18477 2688 18541 2692
rect 18557 2748 18621 2752
rect 18557 2692 18561 2748
rect 18561 2692 18617 2748
rect 18617 2692 18621 2748
rect 18557 2688 18621 2692
rect 25263 2748 25327 2752
rect 25263 2692 25267 2748
rect 25267 2692 25323 2748
rect 25323 2692 25327 2748
rect 25263 2688 25327 2692
rect 25343 2748 25407 2752
rect 25343 2692 25347 2748
rect 25347 2692 25403 2748
rect 25403 2692 25407 2748
rect 25343 2688 25407 2692
rect 25423 2748 25487 2752
rect 25423 2692 25427 2748
rect 25427 2692 25483 2748
rect 25483 2692 25487 2748
rect 25423 2688 25487 2692
rect 25503 2748 25567 2752
rect 25503 2692 25507 2748
rect 25507 2692 25563 2748
rect 25563 2692 25567 2748
rect 25503 2688 25567 2692
rect 7898 2204 7962 2208
rect 7898 2148 7902 2204
rect 7902 2148 7958 2204
rect 7958 2148 7962 2204
rect 7898 2144 7962 2148
rect 7978 2204 8042 2208
rect 7978 2148 7982 2204
rect 7982 2148 8038 2204
rect 8038 2148 8042 2204
rect 7978 2144 8042 2148
rect 8058 2204 8122 2208
rect 8058 2148 8062 2204
rect 8062 2148 8118 2204
rect 8118 2148 8122 2204
rect 8058 2144 8122 2148
rect 8138 2204 8202 2208
rect 8138 2148 8142 2204
rect 8142 2148 8198 2204
rect 8198 2148 8202 2204
rect 8138 2144 8202 2148
rect 14844 2204 14908 2208
rect 14844 2148 14848 2204
rect 14848 2148 14904 2204
rect 14904 2148 14908 2204
rect 14844 2144 14908 2148
rect 14924 2204 14988 2208
rect 14924 2148 14928 2204
rect 14928 2148 14984 2204
rect 14984 2148 14988 2204
rect 14924 2144 14988 2148
rect 15004 2204 15068 2208
rect 15004 2148 15008 2204
rect 15008 2148 15064 2204
rect 15064 2148 15068 2204
rect 15004 2144 15068 2148
rect 15084 2204 15148 2208
rect 15084 2148 15088 2204
rect 15088 2148 15144 2204
rect 15144 2148 15148 2204
rect 15084 2144 15148 2148
rect 21790 2204 21854 2208
rect 21790 2148 21794 2204
rect 21794 2148 21850 2204
rect 21850 2148 21854 2204
rect 21790 2144 21854 2148
rect 21870 2204 21934 2208
rect 21870 2148 21874 2204
rect 21874 2148 21930 2204
rect 21930 2148 21934 2204
rect 21870 2144 21934 2148
rect 21950 2204 22014 2208
rect 21950 2148 21954 2204
rect 21954 2148 22010 2204
rect 22010 2148 22014 2204
rect 21950 2144 22014 2148
rect 22030 2204 22094 2208
rect 22030 2148 22034 2204
rect 22034 2148 22090 2204
rect 22090 2148 22094 2204
rect 22030 2144 22094 2148
rect 28736 2204 28800 2208
rect 28736 2148 28740 2204
rect 28740 2148 28796 2204
rect 28796 2148 28800 2204
rect 28736 2144 28800 2148
rect 28816 2204 28880 2208
rect 28816 2148 28820 2204
rect 28820 2148 28876 2204
rect 28876 2148 28880 2204
rect 28816 2144 28880 2148
rect 28896 2204 28960 2208
rect 28896 2148 28900 2204
rect 28900 2148 28956 2204
rect 28956 2148 28960 2204
rect 28896 2144 28960 2148
rect 28976 2204 29040 2208
rect 28976 2148 28980 2204
rect 28980 2148 29036 2204
rect 29036 2148 29040 2204
rect 28976 2144 29040 2148
<< metal4 >>
rect 4417 47360 4737 47376
rect 4417 47296 4425 47360
rect 4489 47296 4505 47360
rect 4569 47296 4585 47360
rect 4649 47296 4665 47360
rect 4729 47296 4737 47360
rect 4417 46272 4737 47296
rect 4417 46208 4425 46272
rect 4489 46208 4505 46272
rect 4569 46208 4585 46272
rect 4649 46208 4665 46272
rect 4729 46208 4737 46272
rect 4417 45184 4737 46208
rect 4417 45120 4425 45184
rect 4489 45120 4505 45184
rect 4569 45120 4585 45184
rect 4649 45120 4665 45184
rect 4729 45120 4737 45184
rect 4417 44096 4737 45120
rect 4417 44032 4425 44096
rect 4489 44032 4505 44096
rect 4569 44032 4585 44096
rect 4649 44032 4665 44096
rect 4729 44032 4737 44096
rect 4417 43008 4737 44032
rect 4417 42944 4425 43008
rect 4489 42944 4505 43008
rect 4569 42944 4585 43008
rect 4649 42944 4665 43008
rect 4729 42944 4737 43008
rect 4417 41920 4737 42944
rect 4417 41856 4425 41920
rect 4489 41856 4505 41920
rect 4569 41856 4585 41920
rect 4649 41856 4665 41920
rect 4729 41856 4737 41920
rect 4417 40832 4737 41856
rect 4417 40768 4425 40832
rect 4489 40768 4505 40832
rect 4569 40768 4585 40832
rect 4649 40768 4665 40832
rect 4729 40768 4737 40832
rect 4417 39744 4737 40768
rect 4417 39680 4425 39744
rect 4489 39680 4505 39744
rect 4569 39680 4585 39744
rect 4649 39680 4665 39744
rect 4729 39680 4737 39744
rect 4417 38656 4737 39680
rect 4417 38592 4425 38656
rect 4489 38592 4505 38656
rect 4569 38592 4585 38656
rect 4649 38592 4665 38656
rect 4729 38592 4737 38656
rect 4417 37568 4737 38592
rect 4417 37504 4425 37568
rect 4489 37504 4505 37568
rect 4569 37504 4585 37568
rect 4649 37504 4665 37568
rect 4729 37504 4737 37568
rect 4417 36480 4737 37504
rect 4417 36416 4425 36480
rect 4489 36416 4505 36480
rect 4569 36416 4585 36480
rect 4649 36416 4665 36480
rect 4729 36416 4737 36480
rect 4417 35392 4737 36416
rect 4417 35328 4425 35392
rect 4489 35328 4505 35392
rect 4569 35328 4585 35392
rect 4649 35328 4665 35392
rect 4729 35328 4737 35392
rect 4417 34304 4737 35328
rect 4417 34240 4425 34304
rect 4489 34240 4505 34304
rect 4569 34240 4585 34304
rect 4649 34240 4665 34304
rect 4729 34240 4737 34304
rect 4417 33216 4737 34240
rect 4417 33152 4425 33216
rect 4489 33152 4505 33216
rect 4569 33152 4585 33216
rect 4649 33152 4665 33216
rect 4729 33152 4737 33216
rect 4417 32128 4737 33152
rect 4417 32064 4425 32128
rect 4489 32064 4505 32128
rect 4569 32064 4585 32128
rect 4649 32064 4665 32128
rect 4729 32064 4737 32128
rect 4417 31040 4737 32064
rect 4417 30976 4425 31040
rect 4489 30976 4505 31040
rect 4569 30976 4585 31040
rect 4649 30976 4665 31040
rect 4729 30976 4737 31040
rect 4417 29952 4737 30976
rect 4417 29888 4425 29952
rect 4489 29888 4505 29952
rect 4569 29888 4585 29952
rect 4649 29888 4665 29952
rect 4729 29888 4737 29952
rect 4417 28864 4737 29888
rect 4417 28800 4425 28864
rect 4489 28800 4505 28864
rect 4569 28800 4585 28864
rect 4649 28800 4665 28864
rect 4729 28800 4737 28864
rect 4417 27776 4737 28800
rect 4417 27712 4425 27776
rect 4489 27712 4505 27776
rect 4569 27712 4585 27776
rect 4649 27712 4665 27776
rect 4729 27712 4737 27776
rect 4417 26688 4737 27712
rect 4417 26624 4425 26688
rect 4489 26624 4505 26688
rect 4569 26624 4585 26688
rect 4649 26624 4665 26688
rect 4729 26624 4737 26688
rect 4417 25600 4737 26624
rect 4417 25536 4425 25600
rect 4489 25536 4505 25600
rect 4569 25536 4585 25600
rect 4649 25536 4665 25600
rect 4729 25536 4737 25600
rect 4417 24512 4737 25536
rect 4417 24448 4425 24512
rect 4489 24448 4505 24512
rect 4569 24448 4585 24512
rect 4649 24448 4665 24512
rect 4729 24448 4737 24512
rect 4417 23424 4737 24448
rect 4417 23360 4425 23424
rect 4489 23360 4505 23424
rect 4569 23360 4585 23424
rect 4649 23360 4665 23424
rect 4729 23360 4737 23424
rect 4417 22336 4737 23360
rect 4417 22272 4425 22336
rect 4489 22272 4505 22336
rect 4569 22272 4585 22336
rect 4649 22272 4665 22336
rect 4729 22272 4737 22336
rect 4417 21248 4737 22272
rect 4417 21184 4425 21248
rect 4489 21184 4505 21248
rect 4569 21184 4585 21248
rect 4649 21184 4665 21248
rect 4729 21184 4737 21248
rect 4417 20160 4737 21184
rect 4417 20096 4425 20160
rect 4489 20096 4505 20160
rect 4569 20096 4585 20160
rect 4649 20096 4665 20160
rect 4729 20096 4737 20160
rect 4417 19072 4737 20096
rect 4417 19008 4425 19072
rect 4489 19008 4505 19072
rect 4569 19008 4585 19072
rect 4649 19008 4665 19072
rect 4729 19008 4737 19072
rect 4417 17984 4737 19008
rect 4417 17920 4425 17984
rect 4489 17920 4505 17984
rect 4569 17920 4585 17984
rect 4649 17920 4665 17984
rect 4729 17920 4737 17984
rect 4417 16896 4737 17920
rect 4417 16832 4425 16896
rect 4489 16832 4505 16896
rect 4569 16832 4585 16896
rect 4649 16832 4665 16896
rect 4729 16832 4737 16896
rect 4417 15808 4737 16832
rect 4417 15744 4425 15808
rect 4489 15744 4505 15808
rect 4569 15744 4585 15808
rect 4649 15744 4665 15808
rect 4729 15744 4737 15808
rect 4417 14720 4737 15744
rect 4417 14656 4425 14720
rect 4489 14656 4505 14720
rect 4569 14656 4585 14720
rect 4649 14656 4665 14720
rect 4729 14656 4737 14720
rect 4417 13632 4737 14656
rect 4417 13568 4425 13632
rect 4489 13568 4505 13632
rect 4569 13568 4585 13632
rect 4649 13568 4665 13632
rect 4729 13568 4737 13632
rect 4417 12544 4737 13568
rect 4417 12480 4425 12544
rect 4489 12480 4505 12544
rect 4569 12480 4585 12544
rect 4649 12480 4665 12544
rect 4729 12480 4737 12544
rect 4417 11456 4737 12480
rect 4417 11392 4425 11456
rect 4489 11392 4505 11456
rect 4569 11392 4585 11456
rect 4649 11392 4665 11456
rect 4729 11392 4737 11456
rect 4417 10368 4737 11392
rect 4417 10304 4425 10368
rect 4489 10304 4505 10368
rect 4569 10304 4585 10368
rect 4649 10304 4665 10368
rect 4729 10304 4737 10368
rect 4417 9280 4737 10304
rect 4417 9216 4425 9280
rect 4489 9216 4505 9280
rect 4569 9216 4585 9280
rect 4649 9216 4665 9280
rect 4729 9216 4737 9280
rect 4417 8192 4737 9216
rect 4417 8128 4425 8192
rect 4489 8128 4505 8192
rect 4569 8128 4585 8192
rect 4649 8128 4665 8192
rect 4729 8128 4737 8192
rect 4417 7104 4737 8128
rect 4417 7040 4425 7104
rect 4489 7040 4505 7104
rect 4569 7040 4585 7104
rect 4649 7040 4665 7104
rect 4729 7040 4737 7104
rect 4417 6016 4737 7040
rect 4417 5952 4425 6016
rect 4489 5952 4505 6016
rect 4569 5952 4585 6016
rect 4649 5952 4665 6016
rect 4729 5952 4737 6016
rect 4417 4928 4737 5952
rect 4417 4864 4425 4928
rect 4489 4864 4505 4928
rect 4569 4864 4585 4928
rect 4649 4864 4665 4928
rect 4729 4864 4737 4928
rect 4417 3840 4737 4864
rect 4417 3776 4425 3840
rect 4489 3776 4505 3840
rect 4569 3776 4585 3840
rect 4649 3776 4665 3840
rect 4729 3776 4737 3840
rect 4417 2752 4737 3776
rect 4417 2688 4425 2752
rect 4489 2688 4505 2752
rect 4569 2688 4585 2752
rect 4649 2688 4665 2752
rect 4729 2688 4737 2752
rect 4417 2128 4737 2688
rect 7890 46816 8210 47376
rect 7890 46752 7898 46816
rect 7962 46752 7978 46816
rect 8042 46752 8058 46816
rect 8122 46752 8138 46816
rect 8202 46752 8210 46816
rect 7890 45728 8210 46752
rect 7890 45664 7898 45728
rect 7962 45664 7978 45728
rect 8042 45664 8058 45728
rect 8122 45664 8138 45728
rect 8202 45664 8210 45728
rect 7890 44640 8210 45664
rect 7890 44576 7898 44640
rect 7962 44576 7978 44640
rect 8042 44576 8058 44640
rect 8122 44576 8138 44640
rect 8202 44576 8210 44640
rect 7890 43552 8210 44576
rect 7890 43488 7898 43552
rect 7962 43488 7978 43552
rect 8042 43488 8058 43552
rect 8122 43488 8138 43552
rect 8202 43488 8210 43552
rect 7890 42464 8210 43488
rect 7890 42400 7898 42464
rect 7962 42400 7978 42464
rect 8042 42400 8058 42464
rect 8122 42400 8138 42464
rect 8202 42400 8210 42464
rect 7890 41376 8210 42400
rect 7890 41312 7898 41376
rect 7962 41312 7978 41376
rect 8042 41312 8058 41376
rect 8122 41312 8138 41376
rect 8202 41312 8210 41376
rect 7890 40288 8210 41312
rect 7890 40224 7898 40288
rect 7962 40224 7978 40288
rect 8042 40224 8058 40288
rect 8122 40224 8138 40288
rect 8202 40224 8210 40288
rect 7890 39200 8210 40224
rect 7890 39136 7898 39200
rect 7962 39136 7978 39200
rect 8042 39136 8058 39200
rect 8122 39136 8138 39200
rect 8202 39136 8210 39200
rect 7890 38112 8210 39136
rect 7890 38048 7898 38112
rect 7962 38048 7978 38112
rect 8042 38048 8058 38112
rect 8122 38048 8138 38112
rect 8202 38048 8210 38112
rect 7890 37024 8210 38048
rect 7890 36960 7898 37024
rect 7962 36960 7978 37024
rect 8042 36960 8058 37024
rect 8122 36960 8138 37024
rect 8202 36960 8210 37024
rect 7890 35936 8210 36960
rect 7890 35872 7898 35936
rect 7962 35872 7978 35936
rect 8042 35872 8058 35936
rect 8122 35872 8138 35936
rect 8202 35872 8210 35936
rect 7890 34848 8210 35872
rect 7890 34784 7898 34848
rect 7962 34784 7978 34848
rect 8042 34784 8058 34848
rect 8122 34784 8138 34848
rect 8202 34784 8210 34848
rect 7890 33760 8210 34784
rect 7890 33696 7898 33760
rect 7962 33696 7978 33760
rect 8042 33696 8058 33760
rect 8122 33696 8138 33760
rect 8202 33696 8210 33760
rect 7890 32672 8210 33696
rect 7890 32608 7898 32672
rect 7962 32608 7978 32672
rect 8042 32608 8058 32672
rect 8122 32608 8138 32672
rect 8202 32608 8210 32672
rect 7890 31584 8210 32608
rect 7890 31520 7898 31584
rect 7962 31520 7978 31584
rect 8042 31520 8058 31584
rect 8122 31520 8138 31584
rect 8202 31520 8210 31584
rect 7890 30496 8210 31520
rect 7890 30432 7898 30496
rect 7962 30432 7978 30496
rect 8042 30432 8058 30496
rect 8122 30432 8138 30496
rect 8202 30432 8210 30496
rect 7890 29408 8210 30432
rect 7890 29344 7898 29408
rect 7962 29344 7978 29408
rect 8042 29344 8058 29408
rect 8122 29344 8138 29408
rect 8202 29344 8210 29408
rect 7890 28320 8210 29344
rect 7890 28256 7898 28320
rect 7962 28256 7978 28320
rect 8042 28256 8058 28320
rect 8122 28256 8138 28320
rect 8202 28256 8210 28320
rect 7890 27232 8210 28256
rect 7890 27168 7898 27232
rect 7962 27168 7978 27232
rect 8042 27168 8058 27232
rect 8122 27168 8138 27232
rect 8202 27168 8210 27232
rect 7890 26144 8210 27168
rect 7890 26080 7898 26144
rect 7962 26080 7978 26144
rect 8042 26080 8058 26144
rect 8122 26080 8138 26144
rect 8202 26080 8210 26144
rect 7890 25056 8210 26080
rect 7890 24992 7898 25056
rect 7962 24992 7978 25056
rect 8042 24992 8058 25056
rect 8122 24992 8138 25056
rect 8202 24992 8210 25056
rect 7890 23968 8210 24992
rect 7890 23904 7898 23968
rect 7962 23904 7978 23968
rect 8042 23904 8058 23968
rect 8122 23904 8138 23968
rect 8202 23904 8210 23968
rect 7890 22880 8210 23904
rect 7890 22816 7898 22880
rect 7962 22816 7978 22880
rect 8042 22816 8058 22880
rect 8122 22816 8138 22880
rect 8202 22816 8210 22880
rect 7890 21792 8210 22816
rect 7890 21728 7898 21792
rect 7962 21728 7978 21792
rect 8042 21728 8058 21792
rect 8122 21728 8138 21792
rect 8202 21728 8210 21792
rect 7890 20704 8210 21728
rect 7890 20640 7898 20704
rect 7962 20640 7978 20704
rect 8042 20640 8058 20704
rect 8122 20640 8138 20704
rect 8202 20640 8210 20704
rect 7890 19616 8210 20640
rect 7890 19552 7898 19616
rect 7962 19552 7978 19616
rect 8042 19552 8058 19616
rect 8122 19552 8138 19616
rect 8202 19552 8210 19616
rect 7890 18528 8210 19552
rect 7890 18464 7898 18528
rect 7962 18464 7978 18528
rect 8042 18464 8058 18528
rect 8122 18464 8138 18528
rect 8202 18464 8210 18528
rect 7890 17440 8210 18464
rect 7890 17376 7898 17440
rect 7962 17376 7978 17440
rect 8042 17376 8058 17440
rect 8122 17376 8138 17440
rect 8202 17376 8210 17440
rect 7890 16352 8210 17376
rect 7890 16288 7898 16352
rect 7962 16288 7978 16352
rect 8042 16288 8058 16352
rect 8122 16288 8138 16352
rect 8202 16288 8210 16352
rect 7890 15264 8210 16288
rect 7890 15200 7898 15264
rect 7962 15200 7978 15264
rect 8042 15200 8058 15264
rect 8122 15200 8138 15264
rect 8202 15200 8210 15264
rect 7890 14176 8210 15200
rect 7890 14112 7898 14176
rect 7962 14112 7978 14176
rect 8042 14112 8058 14176
rect 8122 14112 8138 14176
rect 8202 14112 8210 14176
rect 7890 13088 8210 14112
rect 7890 13024 7898 13088
rect 7962 13024 7978 13088
rect 8042 13024 8058 13088
rect 8122 13024 8138 13088
rect 8202 13024 8210 13088
rect 7890 12000 8210 13024
rect 7890 11936 7898 12000
rect 7962 11936 7978 12000
rect 8042 11936 8058 12000
rect 8122 11936 8138 12000
rect 8202 11936 8210 12000
rect 7890 10912 8210 11936
rect 7890 10848 7898 10912
rect 7962 10848 7978 10912
rect 8042 10848 8058 10912
rect 8122 10848 8138 10912
rect 8202 10848 8210 10912
rect 7890 9824 8210 10848
rect 7890 9760 7898 9824
rect 7962 9760 7978 9824
rect 8042 9760 8058 9824
rect 8122 9760 8138 9824
rect 8202 9760 8210 9824
rect 7890 8736 8210 9760
rect 7890 8672 7898 8736
rect 7962 8672 7978 8736
rect 8042 8672 8058 8736
rect 8122 8672 8138 8736
rect 8202 8672 8210 8736
rect 7890 7648 8210 8672
rect 7890 7584 7898 7648
rect 7962 7584 7978 7648
rect 8042 7584 8058 7648
rect 8122 7584 8138 7648
rect 8202 7584 8210 7648
rect 7890 6560 8210 7584
rect 7890 6496 7898 6560
rect 7962 6496 7978 6560
rect 8042 6496 8058 6560
rect 8122 6496 8138 6560
rect 8202 6496 8210 6560
rect 7890 5472 8210 6496
rect 7890 5408 7898 5472
rect 7962 5408 7978 5472
rect 8042 5408 8058 5472
rect 8122 5408 8138 5472
rect 8202 5408 8210 5472
rect 7890 4384 8210 5408
rect 7890 4320 7898 4384
rect 7962 4320 7978 4384
rect 8042 4320 8058 4384
rect 8122 4320 8138 4384
rect 8202 4320 8210 4384
rect 7890 3296 8210 4320
rect 7890 3232 7898 3296
rect 7962 3232 7978 3296
rect 8042 3232 8058 3296
rect 8122 3232 8138 3296
rect 8202 3232 8210 3296
rect 7890 2208 8210 3232
rect 7890 2144 7898 2208
rect 7962 2144 7978 2208
rect 8042 2144 8058 2208
rect 8122 2144 8138 2208
rect 8202 2144 8210 2208
rect 7890 2128 8210 2144
rect 11363 47360 11683 47376
rect 11363 47296 11371 47360
rect 11435 47296 11451 47360
rect 11515 47296 11531 47360
rect 11595 47296 11611 47360
rect 11675 47296 11683 47360
rect 11363 46272 11683 47296
rect 11363 46208 11371 46272
rect 11435 46208 11451 46272
rect 11515 46208 11531 46272
rect 11595 46208 11611 46272
rect 11675 46208 11683 46272
rect 11363 45184 11683 46208
rect 11363 45120 11371 45184
rect 11435 45120 11451 45184
rect 11515 45120 11531 45184
rect 11595 45120 11611 45184
rect 11675 45120 11683 45184
rect 11363 44096 11683 45120
rect 11363 44032 11371 44096
rect 11435 44032 11451 44096
rect 11515 44032 11531 44096
rect 11595 44032 11611 44096
rect 11675 44032 11683 44096
rect 11363 43008 11683 44032
rect 11363 42944 11371 43008
rect 11435 42944 11451 43008
rect 11515 42944 11531 43008
rect 11595 42944 11611 43008
rect 11675 42944 11683 43008
rect 11363 41920 11683 42944
rect 11363 41856 11371 41920
rect 11435 41856 11451 41920
rect 11515 41856 11531 41920
rect 11595 41856 11611 41920
rect 11675 41856 11683 41920
rect 11363 40832 11683 41856
rect 11363 40768 11371 40832
rect 11435 40768 11451 40832
rect 11515 40768 11531 40832
rect 11595 40768 11611 40832
rect 11675 40768 11683 40832
rect 11363 39744 11683 40768
rect 11363 39680 11371 39744
rect 11435 39680 11451 39744
rect 11515 39680 11531 39744
rect 11595 39680 11611 39744
rect 11675 39680 11683 39744
rect 11363 38656 11683 39680
rect 11363 38592 11371 38656
rect 11435 38592 11451 38656
rect 11515 38592 11531 38656
rect 11595 38592 11611 38656
rect 11675 38592 11683 38656
rect 11363 37568 11683 38592
rect 11363 37504 11371 37568
rect 11435 37504 11451 37568
rect 11515 37504 11531 37568
rect 11595 37504 11611 37568
rect 11675 37504 11683 37568
rect 11363 36480 11683 37504
rect 11363 36416 11371 36480
rect 11435 36416 11451 36480
rect 11515 36416 11531 36480
rect 11595 36416 11611 36480
rect 11675 36416 11683 36480
rect 11363 35392 11683 36416
rect 11363 35328 11371 35392
rect 11435 35328 11451 35392
rect 11515 35328 11531 35392
rect 11595 35328 11611 35392
rect 11675 35328 11683 35392
rect 11363 34304 11683 35328
rect 11363 34240 11371 34304
rect 11435 34240 11451 34304
rect 11515 34240 11531 34304
rect 11595 34240 11611 34304
rect 11675 34240 11683 34304
rect 11363 33216 11683 34240
rect 11363 33152 11371 33216
rect 11435 33152 11451 33216
rect 11515 33152 11531 33216
rect 11595 33152 11611 33216
rect 11675 33152 11683 33216
rect 11363 32128 11683 33152
rect 11363 32064 11371 32128
rect 11435 32064 11451 32128
rect 11515 32064 11531 32128
rect 11595 32064 11611 32128
rect 11675 32064 11683 32128
rect 11363 31040 11683 32064
rect 11363 30976 11371 31040
rect 11435 30976 11451 31040
rect 11515 30976 11531 31040
rect 11595 30976 11611 31040
rect 11675 30976 11683 31040
rect 11363 29952 11683 30976
rect 11363 29888 11371 29952
rect 11435 29888 11451 29952
rect 11515 29888 11531 29952
rect 11595 29888 11611 29952
rect 11675 29888 11683 29952
rect 11363 28864 11683 29888
rect 11363 28800 11371 28864
rect 11435 28800 11451 28864
rect 11515 28800 11531 28864
rect 11595 28800 11611 28864
rect 11675 28800 11683 28864
rect 11363 27776 11683 28800
rect 11363 27712 11371 27776
rect 11435 27712 11451 27776
rect 11515 27712 11531 27776
rect 11595 27712 11611 27776
rect 11675 27712 11683 27776
rect 11363 26688 11683 27712
rect 11363 26624 11371 26688
rect 11435 26624 11451 26688
rect 11515 26624 11531 26688
rect 11595 26624 11611 26688
rect 11675 26624 11683 26688
rect 11363 25600 11683 26624
rect 11363 25536 11371 25600
rect 11435 25536 11451 25600
rect 11515 25536 11531 25600
rect 11595 25536 11611 25600
rect 11675 25536 11683 25600
rect 11363 24512 11683 25536
rect 11363 24448 11371 24512
rect 11435 24448 11451 24512
rect 11515 24448 11531 24512
rect 11595 24448 11611 24512
rect 11675 24448 11683 24512
rect 11363 23424 11683 24448
rect 11363 23360 11371 23424
rect 11435 23360 11451 23424
rect 11515 23360 11531 23424
rect 11595 23360 11611 23424
rect 11675 23360 11683 23424
rect 11363 22336 11683 23360
rect 11363 22272 11371 22336
rect 11435 22272 11451 22336
rect 11515 22272 11531 22336
rect 11595 22272 11611 22336
rect 11675 22272 11683 22336
rect 11363 21248 11683 22272
rect 11363 21184 11371 21248
rect 11435 21184 11451 21248
rect 11515 21184 11531 21248
rect 11595 21184 11611 21248
rect 11675 21184 11683 21248
rect 11363 20160 11683 21184
rect 11363 20096 11371 20160
rect 11435 20096 11451 20160
rect 11515 20096 11531 20160
rect 11595 20096 11611 20160
rect 11675 20096 11683 20160
rect 11363 19072 11683 20096
rect 11363 19008 11371 19072
rect 11435 19008 11451 19072
rect 11515 19008 11531 19072
rect 11595 19008 11611 19072
rect 11675 19008 11683 19072
rect 11363 17984 11683 19008
rect 11363 17920 11371 17984
rect 11435 17920 11451 17984
rect 11515 17920 11531 17984
rect 11595 17920 11611 17984
rect 11675 17920 11683 17984
rect 11363 16896 11683 17920
rect 11363 16832 11371 16896
rect 11435 16832 11451 16896
rect 11515 16832 11531 16896
rect 11595 16832 11611 16896
rect 11675 16832 11683 16896
rect 11363 15808 11683 16832
rect 11363 15744 11371 15808
rect 11435 15744 11451 15808
rect 11515 15744 11531 15808
rect 11595 15744 11611 15808
rect 11675 15744 11683 15808
rect 11363 14720 11683 15744
rect 11363 14656 11371 14720
rect 11435 14656 11451 14720
rect 11515 14656 11531 14720
rect 11595 14656 11611 14720
rect 11675 14656 11683 14720
rect 11363 13632 11683 14656
rect 11363 13568 11371 13632
rect 11435 13568 11451 13632
rect 11515 13568 11531 13632
rect 11595 13568 11611 13632
rect 11675 13568 11683 13632
rect 11363 12544 11683 13568
rect 11363 12480 11371 12544
rect 11435 12480 11451 12544
rect 11515 12480 11531 12544
rect 11595 12480 11611 12544
rect 11675 12480 11683 12544
rect 11363 11456 11683 12480
rect 11363 11392 11371 11456
rect 11435 11392 11451 11456
rect 11515 11392 11531 11456
rect 11595 11392 11611 11456
rect 11675 11392 11683 11456
rect 11363 10368 11683 11392
rect 11363 10304 11371 10368
rect 11435 10304 11451 10368
rect 11515 10304 11531 10368
rect 11595 10304 11611 10368
rect 11675 10304 11683 10368
rect 11363 9280 11683 10304
rect 11363 9216 11371 9280
rect 11435 9216 11451 9280
rect 11515 9216 11531 9280
rect 11595 9216 11611 9280
rect 11675 9216 11683 9280
rect 11363 8192 11683 9216
rect 11363 8128 11371 8192
rect 11435 8128 11451 8192
rect 11515 8128 11531 8192
rect 11595 8128 11611 8192
rect 11675 8128 11683 8192
rect 11363 7104 11683 8128
rect 11363 7040 11371 7104
rect 11435 7040 11451 7104
rect 11515 7040 11531 7104
rect 11595 7040 11611 7104
rect 11675 7040 11683 7104
rect 11363 6016 11683 7040
rect 11363 5952 11371 6016
rect 11435 5952 11451 6016
rect 11515 5952 11531 6016
rect 11595 5952 11611 6016
rect 11675 5952 11683 6016
rect 11363 4928 11683 5952
rect 11363 4864 11371 4928
rect 11435 4864 11451 4928
rect 11515 4864 11531 4928
rect 11595 4864 11611 4928
rect 11675 4864 11683 4928
rect 11363 3840 11683 4864
rect 11363 3776 11371 3840
rect 11435 3776 11451 3840
rect 11515 3776 11531 3840
rect 11595 3776 11611 3840
rect 11675 3776 11683 3840
rect 11363 2752 11683 3776
rect 11363 2688 11371 2752
rect 11435 2688 11451 2752
rect 11515 2688 11531 2752
rect 11595 2688 11611 2752
rect 11675 2688 11683 2752
rect 11363 2128 11683 2688
rect 14836 46816 15156 47376
rect 14836 46752 14844 46816
rect 14908 46752 14924 46816
rect 14988 46752 15004 46816
rect 15068 46752 15084 46816
rect 15148 46752 15156 46816
rect 14836 45728 15156 46752
rect 14836 45664 14844 45728
rect 14908 45664 14924 45728
rect 14988 45664 15004 45728
rect 15068 45664 15084 45728
rect 15148 45664 15156 45728
rect 14836 44640 15156 45664
rect 14836 44576 14844 44640
rect 14908 44576 14924 44640
rect 14988 44576 15004 44640
rect 15068 44576 15084 44640
rect 15148 44576 15156 44640
rect 14836 43552 15156 44576
rect 14836 43488 14844 43552
rect 14908 43488 14924 43552
rect 14988 43488 15004 43552
rect 15068 43488 15084 43552
rect 15148 43488 15156 43552
rect 14836 42464 15156 43488
rect 14836 42400 14844 42464
rect 14908 42400 14924 42464
rect 14988 42400 15004 42464
rect 15068 42400 15084 42464
rect 15148 42400 15156 42464
rect 14836 41376 15156 42400
rect 14836 41312 14844 41376
rect 14908 41312 14924 41376
rect 14988 41312 15004 41376
rect 15068 41312 15084 41376
rect 15148 41312 15156 41376
rect 14836 40288 15156 41312
rect 14836 40224 14844 40288
rect 14908 40224 14924 40288
rect 14988 40224 15004 40288
rect 15068 40224 15084 40288
rect 15148 40224 15156 40288
rect 14836 39200 15156 40224
rect 14836 39136 14844 39200
rect 14908 39136 14924 39200
rect 14988 39136 15004 39200
rect 15068 39136 15084 39200
rect 15148 39136 15156 39200
rect 14836 38112 15156 39136
rect 14836 38048 14844 38112
rect 14908 38048 14924 38112
rect 14988 38048 15004 38112
rect 15068 38048 15084 38112
rect 15148 38048 15156 38112
rect 14836 37024 15156 38048
rect 14836 36960 14844 37024
rect 14908 36960 14924 37024
rect 14988 36960 15004 37024
rect 15068 36960 15084 37024
rect 15148 36960 15156 37024
rect 14836 35936 15156 36960
rect 14836 35872 14844 35936
rect 14908 35872 14924 35936
rect 14988 35872 15004 35936
rect 15068 35872 15084 35936
rect 15148 35872 15156 35936
rect 14836 34848 15156 35872
rect 14836 34784 14844 34848
rect 14908 34784 14924 34848
rect 14988 34784 15004 34848
rect 15068 34784 15084 34848
rect 15148 34784 15156 34848
rect 14836 33760 15156 34784
rect 14836 33696 14844 33760
rect 14908 33696 14924 33760
rect 14988 33696 15004 33760
rect 15068 33696 15084 33760
rect 15148 33696 15156 33760
rect 14836 32672 15156 33696
rect 14836 32608 14844 32672
rect 14908 32608 14924 32672
rect 14988 32608 15004 32672
rect 15068 32608 15084 32672
rect 15148 32608 15156 32672
rect 14836 31584 15156 32608
rect 14836 31520 14844 31584
rect 14908 31520 14924 31584
rect 14988 31520 15004 31584
rect 15068 31520 15084 31584
rect 15148 31520 15156 31584
rect 14836 30496 15156 31520
rect 14836 30432 14844 30496
rect 14908 30432 14924 30496
rect 14988 30432 15004 30496
rect 15068 30432 15084 30496
rect 15148 30432 15156 30496
rect 14836 29408 15156 30432
rect 14836 29344 14844 29408
rect 14908 29344 14924 29408
rect 14988 29344 15004 29408
rect 15068 29344 15084 29408
rect 15148 29344 15156 29408
rect 14836 28320 15156 29344
rect 14836 28256 14844 28320
rect 14908 28256 14924 28320
rect 14988 28256 15004 28320
rect 15068 28256 15084 28320
rect 15148 28256 15156 28320
rect 14836 27232 15156 28256
rect 14836 27168 14844 27232
rect 14908 27168 14924 27232
rect 14988 27168 15004 27232
rect 15068 27168 15084 27232
rect 15148 27168 15156 27232
rect 14836 26144 15156 27168
rect 14836 26080 14844 26144
rect 14908 26080 14924 26144
rect 14988 26080 15004 26144
rect 15068 26080 15084 26144
rect 15148 26080 15156 26144
rect 14836 25056 15156 26080
rect 14836 24992 14844 25056
rect 14908 24992 14924 25056
rect 14988 24992 15004 25056
rect 15068 24992 15084 25056
rect 15148 24992 15156 25056
rect 14836 23968 15156 24992
rect 14836 23904 14844 23968
rect 14908 23904 14924 23968
rect 14988 23904 15004 23968
rect 15068 23904 15084 23968
rect 15148 23904 15156 23968
rect 14836 22880 15156 23904
rect 14836 22816 14844 22880
rect 14908 22816 14924 22880
rect 14988 22816 15004 22880
rect 15068 22816 15084 22880
rect 15148 22816 15156 22880
rect 14836 21792 15156 22816
rect 14836 21728 14844 21792
rect 14908 21728 14924 21792
rect 14988 21728 15004 21792
rect 15068 21728 15084 21792
rect 15148 21728 15156 21792
rect 14836 20704 15156 21728
rect 14836 20640 14844 20704
rect 14908 20640 14924 20704
rect 14988 20640 15004 20704
rect 15068 20640 15084 20704
rect 15148 20640 15156 20704
rect 14836 19616 15156 20640
rect 14836 19552 14844 19616
rect 14908 19552 14924 19616
rect 14988 19552 15004 19616
rect 15068 19552 15084 19616
rect 15148 19552 15156 19616
rect 14836 18528 15156 19552
rect 14836 18464 14844 18528
rect 14908 18464 14924 18528
rect 14988 18464 15004 18528
rect 15068 18464 15084 18528
rect 15148 18464 15156 18528
rect 14836 17440 15156 18464
rect 14836 17376 14844 17440
rect 14908 17376 14924 17440
rect 14988 17376 15004 17440
rect 15068 17376 15084 17440
rect 15148 17376 15156 17440
rect 14836 16352 15156 17376
rect 14836 16288 14844 16352
rect 14908 16288 14924 16352
rect 14988 16288 15004 16352
rect 15068 16288 15084 16352
rect 15148 16288 15156 16352
rect 14836 15264 15156 16288
rect 14836 15200 14844 15264
rect 14908 15200 14924 15264
rect 14988 15200 15004 15264
rect 15068 15200 15084 15264
rect 15148 15200 15156 15264
rect 14836 14176 15156 15200
rect 14836 14112 14844 14176
rect 14908 14112 14924 14176
rect 14988 14112 15004 14176
rect 15068 14112 15084 14176
rect 15148 14112 15156 14176
rect 14836 13088 15156 14112
rect 14836 13024 14844 13088
rect 14908 13024 14924 13088
rect 14988 13024 15004 13088
rect 15068 13024 15084 13088
rect 15148 13024 15156 13088
rect 14836 12000 15156 13024
rect 14836 11936 14844 12000
rect 14908 11936 14924 12000
rect 14988 11936 15004 12000
rect 15068 11936 15084 12000
rect 15148 11936 15156 12000
rect 14836 10912 15156 11936
rect 14836 10848 14844 10912
rect 14908 10848 14924 10912
rect 14988 10848 15004 10912
rect 15068 10848 15084 10912
rect 15148 10848 15156 10912
rect 14836 9824 15156 10848
rect 14836 9760 14844 9824
rect 14908 9760 14924 9824
rect 14988 9760 15004 9824
rect 15068 9760 15084 9824
rect 15148 9760 15156 9824
rect 14836 8736 15156 9760
rect 14836 8672 14844 8736
rect 14908 8672 14924 8736
rect 14988 8672 15004 8736
rect 15068 8672 15084 8736
rect 15148 8672 15156 8736
rect 14836 7648 15156 8672
rect 14836 7584 14844 7648
rect 14908 7584 14924 7648
rect 14988 7584 15004 7648
rect 15068 7584 15084 7648
rect 15148 7584 15156 7648
rect 14836 6560 15156 7584
rect 14836 6496 14844 6560
rect 14908 6496 14924 6560
rect 14988 6496 15004 6560
rect 15068 6496 15084 6560
rect 15148 6496 15156 6560
rect 14836 5472 15156 6496
rect 14836 5408 14844 5472
rect 14908 5408 14924 5472
rect 14988 5408 15004 5472
rect 15068 5408 15084 5472
rect 15148 5408 15156 5472
rect 14836 4384 15156 5408
rect 14836 4320 14844 4384
rect 14908 4320 14924 4384
rect 14988 4320 15004 4384
rect 15068 4320 15084 4384
rect 15148 4320 15156 4384
rect 14836 3296 15156 4320
rect 14836 3232 14844 3296
rect 14908 3232 14924 3296
rect 14988 3232 15004 3296
rect 15068 3232 15084 3296
rect 15148 3232 15156 3296
rect 14836 2208 15156 3232
rect 14836 2144 14844 2208
rect 14908 2144 14924 2208
rect 14988 2144 15004 2208
rect 15068 2144 15084 2208
rect 15148 2144 15156 2208
rect 14836 2128 15156 2144
rect 18309 47360 18629 47376
rect 18309 47296 18317 47360
rect 18381 47296 18397 47360
rect 18461 47296 18477 47360
rect 18541 47296 18557 47360
rect 18621 47296 18629 47360
rect 18309 46272 18629 47296
rect 18309 46208 18317 46272
rect 18381 46208 18397 46272
rect 18461 46208 18477 46272
rect 18541 46208 18557 46272
rect 18621 46208 18629 46272
rect 18309 45184 18629 46208
rect 18309 45120 18317 45184
rect 18381 45120 18397 45184
rect 18461 45120 18477 45184
rect 18541 45120 18557 45184
rect 18621 45120 18629 45184
rect 18309 44096 18629 45120
rect 18309 44032 18317 44096
rect 18381 44032 18397 44096
rect 18461 44032 18477 44096
rect 18541 44032 18557 44096
rect 18621 44032 18629 44096
rect 18309 43008 18629 44032
rect 18309 42944 18317 43008
rect 18381 42944 18397 43008
rect 18461 42944 18477 43008
rect 18541 42944 18557 43008
rect 18621 42944 18629 43008
rect 18309 41920 18629 42944
rect 18309 41856 18317 41920
rect 18381 41856 18397 41920
rect 18461 41856 18477 41920
rect 18541 41856 18557 41920
rect 18621 41856 18629 41920
rect 18309 40832 18629 41856
rect 18309 40768 18317 40832
rect 18381 40768 18397 40832
rect 18461 40768 18477 40832
rect 18541 40768 18557 40832
rect 18621 40768 18629 40832
rect 18309 39744 18629 40768
rect 18309 39680 18317 39744
rect 18381 39680 18397 39744
rect 18461 39680 18477 39744
rect 18541 39680 18557 39744
rect 18621 39680 18629 39744
rect 18309 38656 18629 39680
rect 18309 38592 18317 38656
rect 18381 38592 18397 38656
rect 18461 38592 18477 38656
rect 18541 38592 18557 38656
rect 18621 38592 18629 38656
rect 18309 37568 18629 38592
rect 18309 37504 18317 37568
rect 18381 37504 18397 37568
rect 18461 37504 18477 37568
rect 18541 37504 18557 37568
rect 18621 37504 18629 37568
rect 18309 36480 18629 37504
rect 18309 36416 18317 36480
rect 18381 36416 18397 36480
rect 18461 36416 18477 36480
rect 18541 36416 18557 36480
rect 18621 36416 18629 36480
rect 18309 35392 18629 36416
rect 18309 35328 18317 35392
rect 18381 35328 18397 35392
rect 18461 35328 18477 35392
rect 18541 35328 18557 35392
rect 18621 35328 18629 35392
rect 18309 34304 18629 35328
rect 18309 34240 18317 34304
rect 18381 34240 18397 34304
rect 18461 34240 18477 34304
rect 18541 34240 18557 34304
rect 18621 34240 18629 34304
rect 18309 33216 18629 34240
rect 18309 33152 18317 33216
rect 18381 33152 18397 33216
rect 18461 33152 18477 33216
rect 18541 33152 18557 33216
rect 18621 33152 18629 33216
rect 18309 32128 18629 33152
rect 18309 32064 18317 32128
rect 18381 32064 18397 32128
rect 18461 32064 18477 32128
rect 18541 32064 18557 32128
rect 18621 32064 18629 32128
rect 18309 31040 18629 32064
rect 18309 30976 18317 31040
rect 18381 30976 18397 31040
rect 18461 30976 18477 31040
rect 18541 30976 18557 31040
rect 18621 30976 18629 31040
rect 18309 29952 18629 30976
rect 18309 29888 18317 29952
rect 18381 29888 18397 29952
rect 18461 29888 18477 29952
rect 18541 29888 18557 29952
rect 18621 29888 18629 29952
rect 18309 28864 18629 29888
rect 18309 28800 18317 28864
rect 18381 28800 18397 28864
rect 18461 28800 18477 28864
rect 18541 28800 18557 28864
rect 18621 28800 18629 28864
rect 18309 27776 18629 28800
rect 21782 46816 22102 47376
rect 21782 46752 21790 46816
rect 21854 46752 21870 46816
rect 21934 46752 21950 46816
rect 22014 46752 22030 46816
rect 22094 46752 22102 46816
rect 21782 45728 22102 46752
rect 21782 45664 21790 45728
rect 21854 45664 21870 45728
rect 21934 45664 21950 45728
rect 22014 45664 22030 45728
rect 22094 45664 22102 45728
rect 21782 44640 22102 45664
rect 21782 44576 21790 44640
rect 21854 44576 21870 44640
rect 21934 44576 21950 44640
rect 22014 44576 22030 44640
rect 22094 44576 22102 44640
rect 21782 43552 22102 44576
rect 21782 43488 21790 43552
rect 21854 43488 21870 43552
rect 21934 43488 21950 43552
rect 22014 43488 22030 43552
rect 22094 43488 22102 43552
rect 21782 42464 22102 43488
rect 21782 42400 21790 42464
rect 21854 42400 21870 42464
rect 21934 42400 21950 42464
rect 22014 42400 22030 42464
rect 22094 42400 22102 42464
rect 21782 41376 22102 42400
rect 21782 41312 21790 41376
rect 21854 41312 21870 41376
rect 21934 41312 21950 41376
rect 22014 41312 22030 41376
rect 22094 41312 22102 41376
rect 21782 40288 22102 41312
rect 21782 40224 21790 40288
rect 21854 40224 21870 40288
rect 21934 40224 21950 40288
rect 22014 40224 22030 40288
rect 22094 40224 22102 40288
rect 21782 39200 22102 40224
rect 21782 39136 21790 39200
rect 21854 39136 21870 39200
rect 21934 39136 21950 39200
rect 22014 39136 22030 39200
rect 22094 39136 22102 39200
rect 21782 38112 22102 39136
rect 21782 38048 21790 38112
rect 21854 38048 21870 38112
rect 21934 38048 21950 38112
rect 22014 38048 22030 38112
rect 22094 38048 22102 38112
rect 21782 37024 22102 38048
rect 21782 36960 21790 37024
rect 21854 36960 21870 37024
rect 21934 36960 21950 37024
rect 22014 36960 22030 37024
rect 22094 36960 22102 37024
rect 21782 35936 22102 36960
rect 21782 35872 21790 35936
rect 21854 35872 21870 35936
rect 21934 35872 21950 35936
rect 22014 35872 22030 35936
rect 22094 35872 22102 35936
rect 21782 34848 22102 35872
rect 21782 34784 21790 34848
rect 21854 34784 21870 34848
rect 21934 34784 21950 34848
rect 22014 34784 22030 34848
rect 22094 34784 22102 34848
rect 21782 33760 22102 34784
rect 21782 33696 21790 33760
rect 21854 33696 21870 33760
rect 21934 33696 21950 33760
rect 22014 33696 22030 33760
rect 22094 33696 22102 33760
rect 21782 32672 22102 33696
rect 21782 32608 21790 32672
rect 21854 32608 21870 32672
rect 21934 32608 21950 32672
rect 22014 32608 22030 32672
rect 22094 32608 22102 32672
rect 21782 31584 22102 32608
rect 21782 31520 21790 31584
rect 21854 31520 21870 31584
rect 21934 31520 21950 31584
rect 22014 31520 22030 31584
rect 22094 31520 22102 31584
rect 21782 30496 22102 31520
rect 21782 30432 21790 30496
rect 21854 30432 21870 30496
rect 21934 30432 21950 30496
rect 22014 30432 22030 30496
rect 22094 30432 22102 30496
rect 21782 29408 22102 30432
rect 21782 29344 21790 29408
rect 21854 29344 21870 29408
rect 21934 29344 21950 29408
rect 22014 29344 22030 29408
rect 22094 29344 22102 29408
rect 21782 28320 22102 29344
rect 21782 28256 21790 28320
rect 21854 28256 21870 28320
rect 21934 28256 21950 28320
rect 22014 28256 22030 28320
rect 22094 28256 22102 28320
rect 18827 27980 18893 27981
rect 18827 27916 18828 27980
rect 18892 27916 18893 27980
rect 18827 27915 18893 27916
rect 18309 27712 18317 27776
rect 18381 27712 18397 27776
rect 18461 27712 18477 27776
rect 18541 27712 18557 27776
rect 18621 27712 18629 27776
rect 18309 26688 18629 27712
rect 18309 26624 18317 26688
rect 18381 26624 18397 26688
rect 18461 26624 18477 26688
rect 18541 26624 18557 26688
rect 18621 26624 18629 26688
rect 18309 25600 18629 26624
rect 18309 25536 18317 25600
rect 18381 25536 18397 25600
rect 18461 25536 18477 25600
rect 18541 25536 18557 25600
rect 18621 25536 18629 25600
rect 18309 24512 18629 25536
rect 18309 24448 18317 24512
rect 18381 24448 18397 24512
rect 18461 24448 18477 24512
rect 18541 24448 18557 24512
rect 18621 24448 18629 24512
rect 18309 23424 18629 24448
rect 18309 23360 18317 23424
rect 18381 23360 18397 23424
rect 18461 23360 18477 23424
rect 18541 23360 18557 23424
rect 18621 23360 18629 23424
rect 18309 22336 18629 23360
rect 18309 22272 18317 22336
rect 18381 22272 18397 22336
rect 18461 22272 18477 22336
rect 18541 22272 18557 22336
rect 18621 22272 18629 22336
rect 18309 21248 18629 22272
rect 18309 21184 18317 21248
rect 18381 21184 18397 21248
rect 18461 21184 18477 21248
rect 18541 21184 18557 21248
rect 18621 21184 18629 21248
rect 18309 20160 18629 21184
rect 18309 20096 18317 20160
rect 18381 20096 18397 20160
rect 18461 20096 18477 20160
rect 18541 20096 18557 20160
rect 18621 20096 18629 20160
rect 18309 19072 18629 20096
rect 18309 19008 18317 19072
rect 18381 19008 18397 19072
rect 18461 19008 18477 19072
rect 18541 19008 18557 19072
rect 18621 19008 18629 19072
rect 18309 17984 18629 19008
rect 18309 17920 18317 17984
rect 18381 17920 18397 17984
rect 18461 17920 18477 17984
rect 18541 17920 18557 17984
rect 18621 17920 18629 17984
rect 18309 16896 18629 17920
rect 18309 16832 18317 16896
rect 18381 16832 18397 16896
rect 18461 16832 18477 16896
rect 18541 16832 18557 16896
rect 18621 16832 18629 16896
rect 18309 15808 18629 16832
rect 18309 15744 18317 15808
rect 18381 15744 18397 15808
rect 18461 15744 18477 15808
rect 18541 15744 18557 15808
rect 18621 15744 18629 15808
rect 18309 14720 18629 15744
rect 18309 14656 18317 14720
rect 18381 14656 18397 14720
rect 18461 14656 18477 14720
rect 18541 14656 18557 14720
rect 18621 14656 18629 14720
rect 18309 13632 18629 14656
rect 18309 13568 18317 13632
rect 18381 13568 18397 13632
rect 18461 13568 18477 13632
rect 18541 13568 18557 13632
rect 18621 13568 18629 13632
rect 18309 12544 18629 13568
rect 18309 12480 18317 12544
rect 18381 12480 18397 12544
rect 18461 12480 18477 12544
rect 18541 12480 18557 12544
rect 18621 12480 18629 12544
rect 18309 11456 18629 12480
rect 18830 11933 18890 27915
rect 21782 27232 22102 28256
rect 21782 27168 21790 27232
rect 21854 27168 21870 27232
rect 21934 27168 21950 27232
rect 22014 27168 22030 27232
rect 22094 27168 22102 27232
rect 21782 26144 22102 27168
rect 21782 26080 21790 26144
rect 21854 26080 21870 26144
rect 21934 26080 21950 26144
rect 22014 26080 22030 26144
rect 22094 26080 22102 26144
rect 21782 25056 22102 26080
rect 21782 24992 21790 25056
rect 21854 24992 21870 25056
rect 21934 24992 21950 25056
rect 22014 24992 22030 25056
rect 22094 24992 22102 25056
rect 21782 23968 22102 24992
rect 21782 23904 21790 23968
rect 21854 23904 21870 23968
rect 21934 23904 21950 23968
rect 22014 23904 22030 23968
rect 22094 23904 22102 23968
rect 21782 22880 22102 23904
rect 21782 22816 21790 22880
rect 21854 22816 21870 22880
rect 21934 22816 21950 22880
rect 22014 22816 22030 22880
rect 22094 22816 22102 22880
rect 21782 21792 22102 22816
rect 21782 21728 21790 21792
rect 21854 21728 21870 21792
rect 21934 21728 21950 21792
rect 22014 21728 22030 21792
rect 22094 21728 22102 21792
rect 21782 20704 22102 21728
rect 21782 20640 21790 20704
rect 21854 20640 21870 20704
rect 21934 20640 21950 20704
rect 22014 20640 22030 20704
rect 22094 20640 22102 20704
rect 21782 19616 22102 20640
rect 21782 19552 21790 19616
rect 21854 19552 21870 19616
rect 21934 19552 21950 19616
rect 22014 19552 22030 19616
rect 22094 19552 22102 19616
rect 21782 18528 22102 19552
rect 21782 18464 21790 18528
rect 21854 18464 21870 18528
rect 21934 18464 21950 18528
rect 22014 18464 22030 18528
rect 22094 18464 22102 18528
rect 21782 17440 22102 18464
rect 21782 17376 21790 17440
rect 21854 17376 21870 17440
rect 21934 17376 21950 17440
rect 22014 17376 22030 17440
rect 22094 17376 22102 17440
rect 21782 16352 22102 17376
rect 21782 16288 21790 16352
rect 21854 16288 21870 16352
rect 21934 16288 21950 16352
rect 22014 16288 22030 16352
rect 22094 16288 22102 16352
rect 21782 15264 22102 16288
rect 21782 15200 21790 15264
rect 21854 15200 21870 15264
rect 21934 15200 21950 15264
rect 22014 15200 22030 15264
rect 22094 15200 22102 15264
rect 21782 14176 22102 15200
rect 21782 14112 21790 14176
rect 21854 14112 21870 14176
rect 21934 14112 21950 14176
rect 22014 14112 22030 14176
rect 22094 14112 22102 14176
rect 21782 13088 22102 14112
rect 21782 13024 21790 13088
rect 21854 13024 21870 13088
rect 21934 13024 21950 13088
rect 22014 13024 22030 13088
rect 22094 13024 22102 13088
rect 21782 12000 22102 13024
rect 21782 11936 21790 12000
rect 21854 11936 21870 12000
rect 21934 11936 21950 12000
rect 22014 11936 22030 12000
rect 22094 11936 22102 12000
rect 18827 11932 18893 11933
rect 18827 11868 18828 11932
rect 18892 11868 18893 11932
rect 18827 11867 18893 11868
rect 18309 11392 18317 11456
rect 18381 11392 18397 11456
rect 18461 11392 18477 11456
rect 18541 11392 18557 11456
rect 18621 11392 18629 11456
rect 18309 10368 18629 11392
rect 18309 10304 18317 10368
rect 18381 10304 18397 10368
rect 18461 10304 18477 10368
rect 18541 10304 18557 10368
rect 18621 10304 18629 10368
rect 18309 9280 18629 10304
rect 18309 9216 18317 9280
rect 18381 9216 18397 9280
rect 18461 9216 18477 9280
rect 18541 9216 18557 9280
rect 18621 9216 18629 9280
rect 18309 8192 18629 9216
rect 18309 8128 18317 8192
rect 18381 8128 18397 8192
rect 18461 8128 18477 8192
rect 18541 8128 18557 8192
rect 18621 8128 18629 8192
rect 18309 7104 18629 8128
rect 18309 7040 18317 7104
rect 18381 7040 18397 7104
rect 18461 7040 18477 7104
rect 18541 7040 18557 7104
rect 18621 7040 18629 7104
rect 18309 6016 18629 7040
rect 18309 5952 18317 6016
rect 18381 5952 18397 6016
rect 18461 5952 18477 6016
rect 18541 5952 18557 6016
rect 18621 5952 18629 6016
rect 18309 4928 18629 5952
rect 18309 4864 18317 4928
rect 18381 4864 18397 4928
rect 18461 4864 18477 4928
rect 18541 4864 18557 4928
rect 18621 4864 18629 4928
rect 18309 3840 18629 4864
rect 18309 3776 18317 3840
rect 18381 3776 18397 3840
rect 18461 3776 18477 3840
rect 18541 3776 18557 3840
rect 18621 3776 18629 3840
rect 18309 2752 18629 3776
rect 18309 2688 18317 2752
rect 18381 2688 18397 2752
rect 18461 2688 18477 2752
rect 18541 2688 18557 2752
rect 18621 2688 18629 2752
rect 18309 2128 18629 2688
rect 21782 10912 22102 11936
rect 21782 10848 21790 10912
rect 21854 10848 21870 10912
rect 21934 10848 21950 10912
rect 22014 10848 22030 10912
rect 22094 10848 22102 10912
rect 21782 9824 22102 10848
rect 21782 9760 21790 9824
rect 21854 9760 21870 9824
rect 21934 9760 21950 9824
rect 22014 9760 22030 9824
rect 22094 9760 22102 9824
rect 21782 8736 22102 9760
rect 21782 8672 21790 8736
rect 21854 8672 21870 8736
rect 21934 8672 21950 8736
rect 22014 8672 22030 8736
rect 22094 8672 22102 8736
rect 21782 7648 22102 8672
rect 21782 7584 21790 7648
rect 21854 7584 21870 7648
rect 21934 7584 21950 7648
rect 22014 7584 22030 7648
rect 22094 7584 22102 7648
rect 21782 6560 22102 7584
rect 21782 6496 21790 6560
rect 21854 6496 21870 6560
rect 21934 6496 21950 6560
rect 22014 6496 22030 6560
rect 22094 6496 22102 6560
rect 21782 5472 22102 6496
rect 21782 5408 21790 5472
rect 21854 5408 21870 5472
rect 21934 5408 21950 5472
rect 22014 5408 22030 5472
rect 22094 5408 22102 5472
rect 21782 4384 22102 5408
rect 21782 4320 21790 4384
rect 21854 4320 21870 4384
rect 21934 4320 21950 4384
rect 22014 4320 22030 4384
rect 22094 4320 22102 4384
rect 21782 3296 22102 4320
rect 21782 3232 21790 3296
rect 21854 3232 21870 3296
rect 21934 3232 21950 3296
rect 22014 3232 22030 3296
rect 22094 3232 22102 3296
rect 21782 2208 22102 3232
rect 21782 2144 21790 2208
rect 21854 2144 21870 2208
rect 21934 2144 21950 2208
rect 22014 2144 22030 2208
rect 22094 2144 22102 2208
rect 21782 2128 22102 2144
rect 25255 47360 25575 47376
rect 25255 47296 25263 47360
rect 25327 47296 25343 47360
rect 25407 47296 25423 47360
rect 25487 47296 25503 47360
rect 25567 47296 25575 47360
rect 25255 46272 25575 47296
rect 25255 46208 25263 46272
rect 25327 46208 25343 46272
rect 25407 46208 25423 46272
rect 25487 46208 25503 46272
rect 25567 46208 25575 46272
rect 25255 45184 25575 46208
rect 25255 45120 25263 45184
rect 25327 45120 25343 45184
rect 25407 45120 25423 45184
rect 25487 45120 25503 45184
rect 25567 45120 25575 45184
rect 25255 44096 25575 45120
rect 25255 44032 25263 44096
rect 25327 44032 25343 44096
rect 25407 44032 25423 44096
rect 25487 44032 25503 44096
rect 25567 44032 25575 44096
rect 25255 43008 25575 44032
rect 25255 42944 25263 43008
rect 25327 42944 25343 43008
rect 25407 42944 25423 43008
rect 25487 42944 25503 43008
rect 25567 42944 25575 43008
rect 25255 41920 25575 42944
rect 25255 41856 25263 41920
rect 25327 41856 25343 41920
rect 25407 41856 25423 41920
rect 25487 41856 25503 41920
rect 25567 41856 25575 41920
rect 25255 40832 25575 41856
rect 25255 40768 25263 40832
rect 25327 40768 25343 40832
rect 25407 40768 25423 40832
rect 25487 40768 25503 40832
rect 25567 40768 25575 40832
rect 25255 39744 25575 40768
rect 25255 39680 25263 39744
rect 25327 39680 25343 39744
rect 25407 39680 25423 39744
rect 25487 39680 25503 39744
rect 25567 39680 25575 39744
rect 25255 38656 25575 39680
rect 25255 38592 25263 38656
rect 25327 38592 25343 38656
rect 25407 38592 25423 38656
rect 25487 38592 25503 38656
rect 25567 38592 25575 38656
rect 25255 37568 25575 38592
rect 25255 37504 25263 37568
rect 25327 37504 25343 37568
rect 25407 37504 25423 37568
rect 25487 37504 25503 37568
rect 25567 37504 25575 37568
rect 25255 36480 25575 37504
rect 25255 36416 25263 36480
rect 25327 36416 25343 36480
rect 25407 36416 25423 36480
rect 25487 36416 25503 36480
rect 25567 36416 25575 36480
rect 25255 35392 25575 36416
rect 25255 35328 25263 35392
rect 25327 35328 25343 35392
rect 25407 35328 25423 35392
rect 25487 35328 25503 35392
rect 25567 35328 25575 35392
rect 25255 34304 25575 35328
rect 25255 34240 25263 34304
rect 25327 34240 25343 34304
rect 25407 34240 25423 34304
rect 25487 34240 25503 34304
rect 25567 34240 25575 34304
rect 25255 33216 25575 34240
rect 25255 33152 25263 33216
rect 25327 33152 25343 33216
rect 25407 33152 25423 33216
rect 25487 33152 25503 33216
rect 25567 33152 25575 33216
rect 25255 32128 25575 33152
rect 25255 32064 25263 32128
rect 25327 32064 25343 32128
rect 25407 32064 25423 32128
rect 25487 32064 25503 32128
rect 25567 32064 25575 32128
rect 25255 31040 25575 32064
rect 25255 30976 25263 31040
rect 25327 30976 25343 31040
rect 25407 30976 25423 31040
rect 25487 30976 25503 31040
rect 25567 30976 25575 31040
rect 25255 29952 25575 30976
rect 25255 29888 25263 29952
rect 25327 29888 25343 29952
rect 25407 29888 25423 29952
rect 25487 29888 25503 29952
rect 25567 29888 25575 29952
rect 25255 28864 25575 29888
rect 25255 28800 25263 28864
rect 25327 28800 25343 28864
rect 25407 28800 25423 28864
rect 25487 28800 25503 28864
rect 25567 28800 25575 28864
rect 25255 27776 25575 28800
rect 25255 27712 25263 27776
rect 25327 27712 25343 27776
rect 25407 27712 25423 27776
rect 25487 27712 25503 27776
rect 25567 27712 25575 27776
rect 25255 26688 25575 27712
rect 25255 26624 25263 26688
rect 25327 26624 25343 26688
rect 25407 26624 25423 26688
rect 25487 26624 25503 26688
rect 25567 26624 25575 26688
rect 25255 25600 25575 26624
rect 25255 25536 25263 25600
rect 25327 25536 25343 25600
rect 25407 25536 25423 25600
rect 25487 25536 25503 25600
rect 25567 25536 25575 25600
rect 25255 24512 25575 25536
rect 25255 24448 25263 24512
rect 25327 24448 25343 24512
rect 25407 24448 25423 24512
rect 25487 24448 25503 24512
rect 25567 24448 25575 24512
rect 25255 23424 25575 24448
rect 25255 23360 25263 23424
rect 25327 23360 25343 23424
rect 25407 23360 25423 23424
rect 25487 23360 25503 23424
rect 25567 23360 25575 23424
rect 25255 22336 25575 23360
rect 25255 22272 25263 22336
rect 25327 22272 25343 22336
rect 25407 22272 25423 22336
rect 25487 22272 25503 22336
rect 25567 22272 25575 22336
rect 25255 21248 25575 22272
rect 25255 21184 25263 21248
rect 25327 21184 25343 21248
rect 25407 21184 25423 21248
rect 25487 21184 25503 21248
rect 25567 21184 25575 21248
rect 25255 20160 25575 21184
rect 25255 20096 25263 20160
rect 25327 20096 25343 20160
rect 25407 20096 25423 20160
rect 25487 20096 25503 20160
rect 25567 20096 25575 20160
rect 25255 19072 25575 20096
rect 25255 19008 25263 19072
rect 25327 19008 25343 19072
rect 25407 19008 25423 19072
rect 25487 19008 25503 19072
rect 25567 19008 25575 19072
rect 25255 17984 25575 19008
rect 25255 17920 25263 17984
rect 25327 17920 25343 17984
rect 25407 17920 25423 17984
rect 25487 17920 25503 17984
rect 25567 17920 25575 17984
rect 25255 16896 25575 17920
rect 25255 16832 25263 16896
rect 25327 16832 25343 16896
rect 25407 16832 25423 16896
rect 25487 16832 25503 16896
rect 25567 16832 25575 16896
rect 25255 15808 25575 16832
rect 25255 15744 25263 15808
rect 25327 15744 25343 15808
rect 25407 15744 25423 15808
rect 25487 15744 25503 15808
rect 25567 15744 25575 15808
rect 25255 14720 25575 15744
rect 25255 14656 25263 14720
rect 25327 14656 25343 14720
rect 25407 14656 25423 14720
rect 25487 14656 25503 14720
rect 25567 14656 25575 14720
rect 25255 13632 25575 14656
rect 25255 13568 25263 13632
rect 25327 13568 25343 13632
rect 25407 13568 25423 13632
rect 25487 13568 25503 13632
rect 25567 13568 25575 13632
rect 25255 12544 25575 13568
rect 25255 12480 25263 12544
rect 25327 12480 25343 12544
rect 25407 12480 25423 12544
rect 25487 12480 25503 12544
rect 25567 12480 25575 12544
rect 25255 11456 25575 12480
rect 25255 11392 25263 11456
rect 25327 11392 25343 11456
rect 25407 11392 25423 11456
rect 25487 11392 25503 11456
rect 25567 11392 25575 11456
rect 25255 10368 25575 11392
rect 25255 10304 25263 10368
rect 25327 10304 25343 10368
rect 25407 10304 25423 10368
rect 25487 10304 25503 10368
rect 25567 10304 25575 10368
rect 25255 9280 25575 10304
rect 25255 9216 25263 9280
rect 25327 9216 25343 9280
rect 25407 9216 25423 9280
rect 25487 9216 25503 9280
rect 25567 9216 25575 9280
rect 25255 8192 25575 9216
rect 25255 8128 25263 8192
rect 25327 8128 25343 8192
rect 25407 8128 25423 8192
rect 25487 8128 25503 8192
rect 25567 8128 25575 8192
rect 25255 7104 25575 8128
rect 25255 7040 25263 7104
rect 25327 7040 25343 7104
rect 25407 7040 25423 7104
rect 25487 7040 25503 7104
rect 25567 7040 25575 7104
rect 25255 6016 25575 7040
rect 25255 5952 25263 6016
rect 25327 5952 25343 6016
rect 25407 5952 25423 6016
rect 25487 5952 25503 6016
rect 25567 5952 25575 6016
rect 25255 4928 25575 5952
rect 25255 4864 25263 4928
rect 25327 4864 25343 4928
rect 25407 4864 25423 4928
rect 25487 4864 25503 4928
rect 25567 4864 25575 4928
rect 25255 3840 25575 4864
rect 25255 3776 25263 3840
rect 25327 3776 25343 3840
rect 25407 3776 25423 3840
rect 25487 3776 25503 3840
rect 25567 3776 25575 3840
rect 25255 2752 25575 3776
rect 25255 2688 25263 2752
rect 25327 2688 25343 2752
rect 25407 2688 25423 2752
rect 25487 2688 25503 2752
rect 25567 2688 25575 2752
rect 25255 2128 25575 2688
rect 28728 46816 29048 47376
rect 28728 46752 28736 46816
rect 28800 46752 28816 46816
rect 28880 46752 28896 46816
rect 28960 46752 28976 46816
rect 29040 46752 29048 46816
rect 28728 45728 29048 46752
rect 28728 45664 28736 45728
rect 28800 45664 28816 45728
rect 28880 45664 28896 45728
rect 28960 45664 28976 45728
rect 29040 45664 29048 45728
rect 28728 44640 29048 45664
rect 28728 44576 28736 44640
rect 28800 44576 28816 44640
rect 28880 44576 28896 44640
rect 28960 44576 28976 44640
rect 29040 44576 29048 44640
rect 28728 43552 29048 44576
rect 28728 43488 28736 43552
rect 28800 43488 28816 43552
rect 28880 43488 28896 43552
rect 28960 43488 28976 43552
rect 29040 43488 29048 43552
rect 28728 42464 29048 43488
rect 28728 42400 28736 42464
rect 28800 42400 28816 42464
rect 28880 42400 28896 42464
rect 28960 42400 28976 42464
rect 29040 42400 29048 42464
rect 28728 41376 29048 42400
rect 28728 41312 28736 41376
rect 28800 41312 28816 41376
rect 28880 41312 28896 41376
rect 28960 41312 28976 41376
rect 29040 41312 29048 41376
rect 28728 40288 29048 41312
rect 28728 40224 28736 40288
rect 28800 40224 28816 40288
rect 28880 40224 28896 40288
rect 28960 40224 28976 40288
rect 29040 40224 29048 40288
rect 28728 39200 29048 40224
rect 28728 39136 28736 39200
rect 28800 39136 28816 39200
rect 28880 39136 28896 39200
rect 28960 39136 28976 39200
rect 29040 39136 29048 39200
rect 28728 38112 29048 39136
rect 28728 38048 28736 38112
rect 28800 38048 28816 38112
rect 28880 38048 28896 38112
rect 28960 38048 28976 38112
rect 29040 38048 29048 38112
rect 28728 37024 29048 38048
rect 28728 36960 28736 37024
rect 28800 36960 28816 37024
rect 28880 36960 28896 37024
rect 28960 36960 28976 37024
rect 29040 36960 29048 37024
rect 28728 35936 29048 36960
rect 28728 35872 28736 35936
rect 28800 35872 28816 35936
rect 28880 35872 28896 35936
rect 28960 35872 28976 35936
rect 29040 35872 29048 35936
rect 28728 34848 29048 35872
rect 28728 34784 28736 34848
rect 28800 34784 28816 34848
rect 28880 34784 28896 34848
rect 28960 34784 28976 34848
rect 29040 34784 29048 34848
rect 28728 33760 29048 34784
rect 28728 33696 28736 33760
rect 28800 33696 28816 33760
rect 28880 33696 28896 33760
rect 28960 33696 28976 33760
rect 29040 33696 29048 33760
rect 28728 32672 29048 33696
rect 28728 32608 28736 32672
rect 28800 32608 28816 32672
rect 28880 32608 28896 32672
rect 28960 32608 28976 32672
rect 29040 32608 29048 32672
rect 28728 31584 29048 32608
rect 28728 31520 28736 31584
rect 28800 31520 28816 31584
rect 28880 31520 28896 31584
rect 28960 31520 28976 31584
rect 29040 31520 29048 31584
rect 28728 30496 29048 31520
rect 28728 30432 28736 30496
rect 28800 30432 28816 30496
rect 28880 30432 28896 30496
rect 28960 30432 28976 30496
rect 29040 30432 29048 30496
rect 28728 29408 29048 30432
rect 28728 29344 28736 29408
rect 28800 29344 28816 29408
rect 28880 29344 28896 29408
rect 28960 29344 28976 29408
rect 29040 29344 29048 29408
rect 28728 28320 29048 29344
rect 28728 28256 28736 28320
rect 28800 28256 28816 28320
rect 28880 28256 28896 28320
rect 28960 28256 28976 28320
rect 29040 28256 29048 28320
rect 28728 27232 29048 28256
rect 28728 27168 28736 27232
rect 28800 27168 28816 27232
rect 28880 27168 28896 27232
rect 28960 27168 28976 27232
rect 29040 27168 29048 27232
rect 28728 26144 29048 27168
rect 28728 26080 28736 26144
rect 28800 26080 28816 26144
rect 28880 26080 28896 26144
rect 28960 26080 28976 26144
rect 29040 26080 29048 26144
rect 28728 25056 29048 26080
rect 28728 24992 28736 25056
rect 28800 24992 28816 25056
rect 28880 24992 28896 25056
rect 28960 24992 28976 25056
rect 29040 24992 29048 25056
rect 28728 23968 29048 24992
rect 28728 23904 28736 23968
rect 28800 23904 28816 23968
rect 28880 23904 28896 23968
rect 28960 23904 28976 23968
rect 29040 23904 29048 23968
rect 28728 22880 29048 23904
rect 28728 22816 28736 22880
rect 28800 22816 28816 22880
rect 28880 22816 28896 22880
rect 28960 22816 28976 22880
rect 29040 22816 29048 22880
rect 28728 21792 29048 22816
rect 28728 21728 28736 21792
rect 28800 21728 28816 21792
rect 28880 21728 28896 21792
rect 28960 21728 28976 21792
rect 29040 21728 29048 21792
rect 28728 20704 29048 21728
rect 28728 20640 28736 20704
rect 28800 20640 28816 20704
rect 28880 20640 28896 20704
rect 28960 20640 28976 20704
rect 29040 20640 29048 20704
rect 28728 19616 29048 20640
rect 28728 19552 28736 19616
rect 28800 19552 28816 19616
rect 28880 19552 28896 19616
rect 28960 19552 28976 19616
rect 29040 19552 29048 19616
rect 28728 18528 29048 19552
rect 28728 18464 28736 18528
rect 28800 18464 28816 18528
rect 28880 18464 28896 18528
rect 28960 18464 28976 18528
rect 29040 18464 29048 18528
rect 28728 17440 29048 18464
rect 28728 17376 28736 17440
rect 28800 17376 28816 17440
rect 28880 17376 28896 17440
rect 28960 17376 28976 17440
rect 29040 17376 29048 17440
rect 28728 16352 29048 17376
rect 28728 16288 28736 16352
rect 28800 16288 28816 16352
rect 28880 16288 28896 16352
rect 28960 16288 28976 16352
rect 29040 16288 29048 16352
rect 28728 15264 29048 16288
rect 28728 15200 28736 15264
rect 28800 15200 28816 15264
rect 28880 15200 28896 15264
rect 28960 15200 28976 15264
rect 29040 15200 29048 15264
rect 28728 14176 29048 15200
rect 28728 14112 28736 14176
rect 28800 14112 28816 14176
rect 28880 14112 28896 14176
rect 28960 14112 28976 14176
rect 29040 14112 29048 14176
rect 28728 13088 29048 14112
rect 28728 13024 28736 13088
rect 28800 13024 28816 13088
rect 28880 13024 28896 13088
rect 28960 13024 28976 13088
rect 29040 13024 29048 13088
rect 28728 12000 29048 13024
rect 28728 11936 28736 12000
rect 28800 11936 28816 12000
rect 28880 11936 28896 12000
rect 28960 11936 28976 12000
rect 29040 11936 29048 12000
rect 28728 10912 29048 11936
rect 28728 10848 28736 10912
rect 28800 10848 28816 10912
rect 28880 10848 28896 10912
rect 28960 10848 28976 10912
rect 29040 10848 29048 10912
rect 28728 9824 29048 10848
rect 28728 9760 28736 9824
rect 28800 9760 28816 9824
rect 28880 9760 28896 9824
rect 28960 9760 28976 9824
rect 29040 9760 29048 9824
rect 28728 8736 29048 9760
rect 28728 8672 28736 8736
rect 28800 8672 28816 8736
rect 28880 8672 28896 8736
rect 28960 8672 28976 8736
rect 29040 8672 29048 8736
rect 28728 7648 29048 8672
rect 28728 7584 28736 7648
rect 28800 7584 28816 7648
rect 28880 7584 28896 7648
rect 28960 7584 28976 7648
rect 29040 7584 29048 7648
rect 28728 6560 29048 7584
rect 28728 6496 28736 6560
rect 28800 6496 28816 6560
rect 28880 6496 28896 6560
rect 28960 6496 28976 6560
rect 29040 6496 29048 6560
rect 28728 5472 29048 6496
rect 28728 5408 28736 5472
rect 28800 5408 28816 5472
rect 28880 5408 28896 5472
rect 28960 5408 28976 5472
rect 29040 5408 29048 5472
rect 28728 4384 29048 5408
rect 28728 4320 28736 4384
rect 28800 4320 28816 4384
rect 28880 4320 28896 4384
rect 28960 4320 28976 4384
rect 29040 4320 29048 4384
rect 28728 3296 29048 4320
rect 28728 3232 28736 3296
rect 28800 3232 28816 3296
rect 28880 3232 28896 3296
rect 28960 3232 28976 3296
rect 29040 3232 29048 3296
rect 28728 2208 29048 3232
rect 28728 2144 28736 2208
rect 28800 2144 28816 2208
rect 28880 2144 28896 2208
rect 28960 2144 28976 2208
rect 29040 2144 29048 2208
rect 28728 2128 29048 2144
use sky130_fd_sc_hd__fill_2  FILLER_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 1380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26
timestamp 1667941163
transform 1 0 3496 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29
timestamp 1667941163
transform 1 0 3772 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 4232 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42
timestamp 1667941163
transform 1 0 4968 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 5428 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54
timestamp 1667941163
transform 1 0 6072 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_69
timestamp 1667941163
transform 1 0 7452 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 7820 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_77 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 8188 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_83
timestamp 1667941163
transform 1 0 8740 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_85
timestamp 1667941163
transform 1 0 8924 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97
timestamp 1667941163
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_109 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113
timestamp 1667941163
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_125
timestamp 1667941163
transform 1 0 12604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_137
timestamp 1667941163
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_141
timestamp 1667941163
transform 1 0 14076 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_146
timestamp 1667941163
transform 1 0 14536 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_158
timestamp 1667941163
transform 1 0 15640 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_166
timestamp 1667941163
transform 1 0 16376 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_169
timestamp 1667941163
transform 1 0 16652 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_194
timestamp 1667941163
transform 1 0 18952 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_197
timestamp 1667941163
transform 1 0 19228 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_209
timestamp 1667941163
transform 1 0 20332 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_221
timestamp 1667941163
transform 1 0 21436 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_225
timestamp 1667941163
transform 1 0 21804 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_237
timestamp 1667941163
transform 1 0 22908 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_249
timestamp 1667941163
transform 1 0 24012 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_253
timestamp 1667941163
transform 1 0 24380 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_278
timestamp 1667941163
transform 1 0 26680 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_281
timestamp 1667941163
transform 1 0 26956 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_286
timestamp 1667941163
transform 1 0 27416 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_293
timestamp 1667941163
transform 1 0 28060 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_3
timestamp 1667941163
transform 1 0 1380 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_10
timestamp 1667941163
transform 1 0 2024 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_17
timestamp 1667941163
transform 1 0 2668 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_24
timestamp 1667941163
transform 1 0 3312 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_49
timestamp 1667941163
transform 1 0 5612 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1667941163
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_57
timestamp 1667941163
transform 1 0 6348 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_80
timestamp 1667941163
transform 1 0 8464 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_84
timestamp 1667941163
transform 1 0 8832 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_106
timestamp 1667941163
transform 1 0 10856 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_1_113
timestamp 1667941163
transform 1 0 11500 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_1_136
timestamp 1667941163
transform 1 0 13616 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_142
timestamp 1667941163
transform 1 0 14168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_164
timestamp 1667941163
transform 1 0 16192 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_169
timestamp 1667941163
transform 1 0 16652 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_192
timestamp 1667941163
transform 1 0 18768 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_196
timestamp 1667941163
transform 1 0 19136 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_218
timestamp 1667941163
transform 1 0 21160 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_1_225
timestamp 1667941163
transform 1 0 21804 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_248
timestamp 1667941163
transform 1 0 23920 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_273
timestamp 1667941163
transform 1 0 26220 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_279
timestamp 1667941163
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_281
timestamp 1667941163
transform 1 0 26956 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_286
timestamp 1667941163
transform 1 0 27416 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_293
timestamp 1667941163
transform 1 0 28060 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_2_3
timestamp 1667941163
transform 1 0 1380 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_26
timestamp 1667941163
transform 1 0 3496 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_2_29
timestamp 1667941163
transform 1 0 3772 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_35
timestamp 1667941163
transform 1 0 4324 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_39
timestamp 1667941163
transform 1 0 4692 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_64
timestamp 1667941163
transform 1 0 6992 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_72
timestamp 1667941163
transform 1 0 7728 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_76
timestamp 1667941163
transform 1 0 8096 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_85
timestamp 1667941163
transform 1 0 8924 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_90
timestamp 1667941163
transform 1 0 9384 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_97
timestamp 1667941163
transform 1 0 10028 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_106
timestamp 1667941163
transform 1 0 10856 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_113
timestamp 1667941163
transform 1 0 11500 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_138
timestamp 1667941163
transform 1 0 13800 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_141
timestamp 1667941163
transform 1 0 14076 0 1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_2_147
timestamp 1667941163
transform 1 0 14628 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_159
timestamp 1667941163
transform 1 0 15732 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_166
timestamp 1667941163
transform 1 0 16376 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_173
timestamp 1667941163
transform 1 0 17020 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_180
timestamp 1667941163
transform 1 0 17664 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_187
timestamp 1667941163
transform 1 0 18308 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 1667941163
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_197
timestamp 1667941163
transform 1 0 19228 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_202
timestamp 1667941163
transform 1 0 19688 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_209
timestamp 1667941163
transform 1 0 20332 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_217
timestamp 1667941163
transform 1 0 21068 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_223
timestamp 1667941163
transform 1 0 21620 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_230
timestamp 1667941163
transform 1 0 22264 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_242
timestamp 1667941163
transform 1 0 23368 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_246
timestamp 1667941163
transform 1 0 23736 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_250
timestamp 1667941163
transform 1 0 24104 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_253
timestamp 1667941163
transform 1 0 24380 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_258
timestamp 1667941163
transform 1 0 24840 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_266
timestamp 1667941163
transform 1 0 25576 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_288
timestamp 1667941163
transform 1 0 27600 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_295
timestamp 1667941163
transform 1 0 28244 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_3_3
timestamp 1667941163
transform 1 0 1380 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_27
timestamp 1667941163
transform 1 0 3588 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_52
timestamp 1667941163
transform 1 0 5888 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_57
timestamp 1667941163
transform 1 0 6348 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_62
timestamp 1667941163
transform 1 0 6808 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_70
timestamp 1667941163
transform 1 0 7544 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_93
timestamp 1667941163
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp 1667941163
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1667941163
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_113
timestamp 1667941163
transform 1 0 11500 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_117
timestamp 1667941163
transform 1 0 11868 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_121
timestamp 1667941163
transform 1 0 12236 0 -1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_3_148
timestamp 1667941163
transform 1 0 14720 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_160
timestamp 1667941163
transform 1 0 15824 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_3_169
timestamp 1667941163
transform 1 0 16652 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_173
timestamp 1667941163
transform 1 0 17020 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_177
timestamp 1667941163
transform 1 0 17388 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_189
timestamp 1667941163
transform 1 0 18492 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_201
timestamp 1667941163
transform 1 0 19596 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_209
timestamp 1667941163
transform 1 0 20332 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_214
timestamp 1667941163
transform 1 0 20792 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_222
timestamp 1667941163
transform 1 0 21528 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_225
timestamp 1667941163
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_237
timestamp 1667941163
transform 1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_249
timestamp 1667941163
transform 1 0 24012 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_278
timestamp 1667941163
transform 1 0 26680 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_281
timestamp 1667941163
transform 1 0 26956 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_286
timestamp 1667941163
transform 1 0 27416 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_290
timestamp 1667941163
transform 1 0 27784 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_294
timestamp 1667941163
transform 1 0 28152 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_298
timestamp 1667941163
transform 1 0 28520 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_3
timestamp 1667941163
transform 1 0 1380 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_7
timestamp 1667941163
transform 1 0 1748 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_11
timestamp 1667941163
transform 1 0 2116 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_19
timestamp 1667941163
transform 1 0 2852 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_23
timestamp 1667941163
transform 1 0 3220 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1667941163
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_29
timestamp 1667941163
transform 1 0 3772 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_34
timestamp 1667941163
transform 1 0 4232 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_41
timestamp 1667941163
transform 1 0 4876 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_48
timestamp 1667941163
transform 1 0 5520 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_52
timestamp 1667941163
transform 1 0 5888 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_56
timestamp 1667941163
transform 1 0 6256 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_68
timestamp 1667941163
transform 1 0 7360 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_80
timestamp 1667941163
transform 1 0 8464 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1667941163
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_97
timestamp 1667941163
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_109
timestamp 1667941163
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_121
timestamp 1667941163
transform 1 0 12236 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_127
timestamp 1667941163
transform 1 0 12788 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_131
timestamp 1667941163
transform 1 0 13156 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1667941163
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_141
timestamp 1667941163
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_153
timestamp 1667941163
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_165
timestamp 1667941163
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_177
timestamp 1667941163
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_189
timestamp 1667941163
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 1667941163
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_197
timestamp 1667941163
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_209
timestamp 1667941163
transform 1 0 20332 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_231
timestamp 1667941163
transform 1 0 22356 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_243
timestamp 1667941163
transform 1 0 23460 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_251
timestamp 1667941163
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_253
timestamp 1667941163
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_265
timestamp 1667941163
transform 1 0 25484 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_271
timestamp 1667941163
transform 1 0 26036 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_275
timestamp 1667941163
transform 1 0 26404 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_297
timestamp 1667941163
transform 1 0 28428 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_3
timestamp 1667941163
transform 1 0 1380 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_7
timestamp 1667941163
transform 1 0 1748 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_11
timestamp 1667941163
transform 1 0 2116 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_5_40
timestamp 1667941163
transform 1 0 4784 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_47
timestamp 1667941163
transform 1 0 5428 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1667941163
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1667941163
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1667941163
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_81
timestamp 1667941163
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_93
timestamp 1667941163
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 1667941163
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1667941163
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_113
timestamp 1667941163
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_125
timestamp 1667941163
transform 1 0 12604 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_130
timestamp 1667941163
transform 1 0 13064 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_142
timestamp 1667941163
transform 1 0 14168 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_154
timestamp 1667941163
transform 1 0 15272 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_166
timestamp 1667941163
transform 1 0 16376 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_169
timestamp 1667941163
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_181
timestamp 1667941163
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_193
timestamp 1667941163
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_205
timestamp 1667941163
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_217
timestamp 1667941163
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_223
timestamp 1667941163
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_225
timestamp 1667941163
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_237
timestamp 1667941163
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_249
timestamp 1667941163
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_261
timestamp 1667941163
transform 1 0 25116 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_273
timestamp 1667941163
transform 1 0 26220 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_279
timestamp 1667941163
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_281
timestamp 1667941163
transform 1 0 26956 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_289
timestamp 1667941163
transform 1 0 27692 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_294
timestamp 1667941163
transform 1 0 28152 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_298
timestamp 1667941163
transform 1 0 28520 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_3
timestamp 1667941163
transform 1 0 1380 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_26
timestamp 1667941163
transform 1 0 3496 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_29
timestamp 1667941163
transform 1 0 3772 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_6_35
timestamp 1667941163
transform 1 0 4324 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_47
timestamp 1667941163
transform 1 0 5428 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_59
timestamp 1667941163
transform 1 0 6532 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_71
timestamp 1667941163
transform 1 0 7636 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1667941163
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1667941163
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_97
timestamp 1667941163
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_109
timestamp 1667941163
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_121
timestamp 1667941163
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1667941163
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1667941163
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_141
timestamp 1667941163
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_153
timestamp 1667941163
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_165
timestamp 1667941163
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_177
timestamp 1667941163
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_189
timestamp 1667941163
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1667941163
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_197
timestamp 1667941163
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_209
timestamp 1667941163
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_221
timestamp 1667941163
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_233
timestamp 1667941163
transform 1 0 22540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_245
timestamp 1667941163
transform 1 0 23644 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp 1667941163
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_253
timestamp 1667941163
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_265
timestamp 1667941163
transform 1 0 25484 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_6_273
timestamp 1667941163
transform 1 0 26220 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_297
timestamp 1667941163
transform 1 0 28428 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_3
timestamp 1667941163
transform 1 0 1380 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_27
timestamp 1667941163
transform 1 0 3588 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_52
timestamp 1667941163
transform 1 0 5888 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1667941163
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_69
timestamp 1667941163
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_81
timestamp 1667941163
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_93
timestamp 1667941163
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 1667941163
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1667941163
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_113
timestamp 1667941163
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_125
timestamp 1667941163
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_137
timestamp 1667941163
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_149
timestamp 1667941163
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_161
timestamp 1667941163
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1667941163
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_169
timestamp 1667941163
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_181
timestamp 1667941163
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_193
timestamp 1667941163
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_205
timestamp 1667941163
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_217
timestamp 1667941163
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp 1667941163
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_225
timestamp 1667941163
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_237
timestamp 1667941163
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_249
timestamp 1667941163
transform 1 0 24012 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_261
timestamp 1667941163
transform 1 0 25116 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_273
timestamp 1667941163
transform 1 0 26220 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_279
timestamp 1667941163
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_281
timestamp 1667941163
transform 1 0 26956 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_286
timestamp 1667941163
transform 1 0 27416 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_293
timestamp 1667941163
transform 1 0 28060 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_8_3
timestamp 1667941163
transform 1 0 1380 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_8
timestamp 1667941163
transform 1 0 1840 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_15
timestamp 1667941163
transform 1 0 2484 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_22
timestamp 1667941163
transform 1 0 3128 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_8_29
timestamp 1667941163
transform 1 0 3772 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_36
timestamp 1667941163
transform 1 0 4416 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_44
timestamp 1667941163
transform 1 0 5152 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_49
timestamp 1667941163
transform 1 0 5612 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_74
timestamp 1667941163
transform 1 0 7912 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_82
timestamp 1667941163
transform 1 0 8648 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_85
timestamp 1667941163
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_97
timestamp 1667941163
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_109
timestamp 1667941163
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_121
timestamp 1667941163
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_133
timestamp 1667941163
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1667941163
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_141
timestamp 1667941163
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_153
timestamp 1667941163
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_165
timestamp 1667941163
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_177
timestamp 1667941163
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_189
timestamp 1667941163
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1667941163
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_197
timestamp 1667941163
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_209
timestamp 1667941163
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_221
timestamp 1667941163
transform 1 0 21436 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_233
timestamp 1667941163
transform 1 0 22540 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_245
timestamp 1667941163
transform 1 0 23644 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_251
timestamp 1667941163
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_253
timestamp 1667941163
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_265
timestamp 1667941163
transform 1 0 25484 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_272
timestamp 1667941163
transform 1 0 26128 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_297
timestamp 1667941163
transform 1 0 28428 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_3
timestamp 1667941163
transform 1 0 1380 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_10
timestamp 1667941163
transform 1 0 2024 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_18
timestamp 1667941163
transform 1 0 2760 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_42
timestamp 1667941163
transform 1 0 4968 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_54
timestamp 1667941163
transform 1 0 6072 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 1667941163
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_69
timestamp 1667941163
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_81
timestamp 1667941163
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_93
timestamp 1667941163
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_105
timestamp 1667941163
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1667941163
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_113
timestamp 1667941163
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_125
timestamp 1667941163
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_137
timestamp 1667941163
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_149
timestamp 1667941163
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_161
timestamp 1667941163
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1667941163
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_169
timestamp 1667941163
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_181
timestamp 1667941163
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_193
timestamp 1667941163
transform 1 0 18860 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_205
timestamp 1667941163
transform 1 0 19964 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_217
timestamp 1667941163
transform 1 0 21068 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_223
timestamp 1667941163
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_225
timestamp 1667941163
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_237
timestamp 1667941163
transform 1 0 22908 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_249
timestamp 1667941163
transform 1 0 24012 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_278
timestamp 1667941163
transform 1 0 26680 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_281
timestamp 1667941163
transform 1 0 26956 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_286
timestamp 1667941163
transform 1 0 27416 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_293
timestamp 1667941163
transform 1 0 28060 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_10_3
timestamp 1667941163
transform 1 0 1380 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_9
timestamp 1667941163
transform 1 0 1932 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_16
timestamp 1667941163
transform 1 0 2576 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_10_25
timestamp 1667941163
transform 1 0 3404 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_29
timestamp 1667941163
transform 1 0 3772 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_34
timestamp 1667941163
transform 1 0 4232 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_46
timestamp 1667941163
transform 1 0 5336 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_58
timestamp 1667941163
transform 1 0 6440 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_70
timestamp 1667941163
transform 1 0 7544 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_10_82
timestamp 1667941163
transform 1 0 8648 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_85
timestamp 1667941163
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_97
timestamp 1667941163
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_109
timestamp 1667941163
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_121
timestamp 1667941163
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_133
timestamp 1667941163
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1667941163
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_141
timestamp 1667941163
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_153
timestamp 1667941163
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_165
timestamp 1667941163
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_177
timestamp 1667941163
transform 1 0 17388 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_189
timestamp 1667941163
transform 1 0 18492 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_195
timestamp 1667941163
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_197
timestamp 1667941163
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_209
timestamp 1667941163
transform 1 0 20332 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_221
timestamp 1667941163
transform 1 0 21436 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_233
timestamp 1667941163
transform 1 0 22540 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_245
timestamp 1667941163
transform 1 0 23644 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_251
timestamp 1667941163
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_253
timestamp 1667941163
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_265
timestamp 1667941163
transform 1 0 25484 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_272
timestamp 1667941163
transform 1 0 26128 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_297
timestamp 1667941163
transform 1 0 28428 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_3
timestamp 1667941163
transform 1 0 1380 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_10
timestamp 1667941163
transform 1 0 2024 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_11_35
timestamp 1667941163
transform 1 0 4324 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_47
timestamp 1667941163
transform 1 0 5428 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1667941163
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_57
timestamp 1667941163
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_69
timestamp 1667941163
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_81
timestamp 1667941163
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_93
timestamp 1667941163
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_105
timestamp 1667941163
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1667941163
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_113
timestamp 1667941163
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_125
timestamp 1667941163
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_137
timestamp 1667941163
transform 1 0 13708 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_149
timestamp 1667941163
transform 1 0 14812 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_161
timestamp 1667941163
transform 1 0 15916 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp 1667941163
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_169
timestamp 1667941163
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_181
timestamp 1667941163
transform 1 0 17756 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_193
timestamp 1667941163
transform 1 0 18860 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_205
timestamp 1667941163
transform 1 0 19964 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_217
timestamp 1667941163
transform 1 0 21068 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_223
timestamp 1667941163
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_225
timestamp 1667941163
transform 1 0 21804 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_237
timestamp 1667941163
transform 1 0 22908 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_249
timestamp 1667941163
transform 1 0 24012 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_261
timestamp 1667941163
transform 1 0 25116 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_273
timestamp 1667941163
transform 1 0 26220 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_278
timestamp 1667941163
transform 1 0 26680 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_281
timestamp 1667941163
transform 1 0 26956 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_286
timestamp 1667941163
transform 1 0 27416 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_293
timestamp 1667941163
transform 1 0 28060 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_12_3
timestamp 1667941163
transform 1 0 1380 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_26
timestamp 1667941163
transform 1 0 3496 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_29
timestamp 1667941163
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_41
timestamp 1667941163
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_53
timestamp 1667941163
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_65
timestamp 1667941163
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 1667941163
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1667941163
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_85
timestamp 1667941163
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_97
timestamp 1667941163
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_109
timestamp 1667941163
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_121
timestamp 1667941163
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_133
timestamp 1667941163
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1667941163
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_141
timestamp 1667941163
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_153
timestamp 1667941163
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_165
timestamp 1667941163
transform 1 0 16284 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_177
timestamp 1667941163
transform 1 0 17388 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_189
timestamp 1667941163
transform 1 0 18492 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_195
timestamp 1667941163
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_197
timestamp 1667941163
transform 1 0 19228 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_209
timestamp 1667941163
transform 1 0 20332 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_221
timestamp 1667941163
transform 1 0 21436 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_233
timestamp 1667941163
transform 1 0 22540 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_245
timestamp 1667941163
transform 1 0 23644 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_251
timestamp 1667941163
transform 1 0 24196 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_253
timestamp 1667941163
transform 1 0 24380 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_265
timestamp 1667941163
transform 1 0 25484 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_12_273
timestamp 1667941163
transform 1 0 26220 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_297
timestamp 1667941163
transform 1 0 28428 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_3
timestamp 1667941163
transform 1 0 1380 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_27
timestamp 1667941163
transform 1 0 3588 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_34
timestamp 1667941163
transform 1 0 4232 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_46
timestamp 1667941163
transform 1 0 5336 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_54
timestamp 1667941163
transform 1 0 6072 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_57
timestamp 1667941163
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_69
timestamp 1667941163
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_81
timestamp 1667941163
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_93
timestamp 1667941163
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_105
timestamp 1667941163
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1667941163
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_113
timestamp 1667941163
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_125
timestamp 1667941163
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_137
timestamp 1667941163
transform 1 0 13708 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_149
timestamp 1667941163
transform 1 0 14812 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_161
timestamp 1667941163
transform 1 0 15916 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 1667941163
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_169
timestamp 1667941163
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_181
timestamp 1667941163
transform 1 0 17756 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_193
timestamp 1667941163
transform 1 0 18860 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_205
timestamp 1667941163
transform 1 0 19964 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_209
timestamp 1667941163
transform 1 0 20332 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_213
timestamp 1667941163
transform 1 0 20700 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_221
timestamp 1667941163
transform 1 0 21436 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_225
timestamp 1667941163
transform 1 0 21804 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_237
timestamp 1667941163
transform 1 0 22908 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_249
timestamp 1667941163
transform 1 0 24012 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_261
timestamp 1667941163
transform 1 0 25116 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_273
timestamp 1667941163
transform 1 0 26220 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_279
timestamp 1667941163
transform 1 0 26772 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_281
timestamp 1667941163
transform 1 0 26956 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_13_292
timestamp 1667941163
transform 1 0 27968 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_298
timestamp 1667941163
transform 1 0 28520 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_14_3
timestamp 1667941163
transform 1 0 1380 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_14_9
timestamp 1667941163
transform 1 0 1932 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_17
timestamp 1667941163
transform 1 0 2668 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_14_22
timestamp 1667941163
transform 1 0 3128 0 1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_14_29
timestamp 1667941163
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_41
timestamp 1667941163
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_53
timestamp 1667941163
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_65
timestamp 1667941163
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp 1667941163
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1667941163
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_85
timestamp 1667941163
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_97
timestamp 1667941163
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_109
timestamp 1667941163
transform 1 0 11132 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_121
timestamp 1667941163
transform 1 0 12236 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_133
timestamp 1667941163
transform 1 0 13340 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1667941163
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_141
timestamp 1667941163
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_153
timestamp 1667941163
transform 1 0 15180 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_165
timestamp 1667941163
transform 1 0 16284 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_177
timestamp 1667941163
transform 1 0 17388 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_187
timestamp 1667941163
transform 1 0 18308 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_195
timestamp 1667941163
transform 1 0 19044 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_197
timestamp 1667941163
transform 1 0 19228 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_204
timestamp 1667941163
transform 1 0 19872 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_216
timestamp 1667941163
transform 1 0 20976 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_228
timestamp 1667941163
transform 1 0 22080 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_240
timestamp 1667941163
transform 1 0 23184 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_253
timestamp 1667941163
transform 1 0 24380 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_265
timestamp 1667941163
transform 1 0 25484 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_273
timestamp 1667941163
transform 1 0 26220 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_297
timestamp 1667941163
transform 1 0 28428 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3
timestamp 1667941163
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_15
timestamp 1667941163
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_27
timestamp 1667941163
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_39
timestamp 1667941163
transform 1 0 4692 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_51
timestamp 1667941163
transform 1 0 5796 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1667941163
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_57
timestamp 1667941163
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_69
timestamp 1667941163
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_81
timestamp 1667941163
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_93
timestamp 1667941163
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_105
timestamp 1667941163
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1667941163
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_113
timestamp 1667941163
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_125
timestamp 1667941163
transform 1 0 12604 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_137
timestamp 1667941163
transform 1 0 13708 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_149
timestamp 1667941163
transform 1 0 14812 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_161
timestamp 1667941163
transform 1 0 15916 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_167
timestamp 1667941163
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_169
timestamp 1667941163
transform 1 0 16652 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_177
timestamp 1667941163
transform 1 0 17388 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_187
timestamp 1667941163
transform 1 0 18308 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_198
timestamp 1667941163
transform 1 0 19320 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_209
timestamp 1667941163
transform 1 0 20332 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_15_221
timestamp 1667941163
transform 1 0 21436 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_15_225
timestamp 1667941163
transform 1 0 21804 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_237
timestamp 1667941163
transform 1 0 22908 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_249
timestamp 1667941163
transform 1 0 24012 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_261
timestamp 1667941163
transform 1 0 25116 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_273
timestamp 1667941163
transform 1 0 26220 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_279
timestamp 1667941163
transform 1 0 26772 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_281
timestamp 1667941163
transform 1 0 26956 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_286
timestamp 1667941163
transform 1 0 27416 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_293
timestamp 1667941163
transform 1 0 28060 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_16_3
timestamp 1667941163
transform 1 0 1380 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_10
timestamp 1667941163
transform 1 0 2024 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_22
timestamp 1667941163
transform 1 0 3128 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_16_29
timestamp 1667941163
transform 1 0 3772 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_43
timestamp 1667941163
transform 1 0 5060 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_55
timestamp 1667941163
transform 1 0 6164 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_67
timestamp 1667941163
transform 1 0 7268 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_79
timestamp 1667941163
transform 1 0 8372 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1667941163
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_85
timestamp 1667941163
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_97
timestamp 1667941163
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_109
timestamp 1667941163
transform 1 0 11132 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_121
timestamp 1667941163
transform 1 0 12236 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_133
timestamp 1667941163
transform 1 0 13340 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 1667941163
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_141
timestamp 1667941163
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_153
timestamp 1667941163
transform 1 0 15180 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_165
timestamp 1667941163
transform 1 0 16284 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_16_177
timestamp 1667941163
transform 1 0 17388 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_16_183
timestamp 1667941163
transform 1 0 17940 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_16_194
timestamp 1667941163
transform 1 0 18952 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_197
timestamp 1667941163
transform 1 0 19228 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_209
timestamp 1667941163
transform 1 0 20332 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_221
timestamp 1667941163
transform 1 0 21436 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_233
timestamp 1667941163
transform 1 0 22540 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_245
timestamp 1667941163
transform 1 0 23644 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_251
timestamp 1667941163
transform 1 0 24196 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_253
timestamp 1667941163
transform 1 0 24380 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_265
timestamp 1667941163
transform 1 0 25484 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_16_273
timestamp 1667941163
transform 1 0 26220 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_297
timestamp 1667941163
transform 1 0 28428 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_3
timestamp 1667941163
transform 1 0 1380 0 -1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_17_27
timestamp 1667941163
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_39
timestamp 1667941163
transform 1 0 4692 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_51
timestamp 1667941163
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1667941163
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_57
timestamp 1667941163
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_69
timestamp 1667941163
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_81
timestamp 1667941163
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_93
timestamp 1667941163
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_105
timestamp 1667941163
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1667941163
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_113
timestamp 1667941163
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_125
timestamp 1667941163
transform 1 0 12604 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_137
timestamp 1667941163
transform 1 0 13708 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_149
timestamp 1667941163
transform 1 0 14812 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_161
timestamp 1667941163
transform 1 0 15916 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_167
timestamp 1667941163
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_169
timestamp 1667941163
transform 1 0 16652 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_17_180
timestamp 1667941163
transform 1 0 17664 0 -1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_17_195
timestamp 1667941163
transform 1 0 19044 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_207
timestamp 1667941163
transform 1 0 20148 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_219
timestamp 1667941163
transform 1 0 21252 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_223
timestamp 1667941163
transform 1 0 21620 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_225
timestamp 1667941163
transform 1 0 21804 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_237
timestamp 1667941163
transform 1 0 22908 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_249
timestamp 1667941163
transform 1 0 24012 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_261
timestamp 1667941163
transform 1 0 25116 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_273
timestamp 1667941163
transform 1 0 26220 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_279
timestamp 1667941163
transform 1 0 26772 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_281
timestamp 1667941163
transform 1 0 26956 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_286
timestamp 1667941163
transform 1 0 27416 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_17_298
timestamp 1667941163
transform 1 0 28520 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_18_3
timestamp 1667941163
transform 1 0 1380 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_18_9
timestamp 1667941163
transform 1 0 1932 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_21
timestamp 1667941163
transform 1 0 3036 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1667941163
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_29
timestamp 1667941163
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_41
timestamp 1667941163
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_53
timestamp 1667941163
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_65
timestamp 1667941163
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_77
timestamp 1667941163
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1667941163
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_85
timestamp 1667941163
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_97
timestamp 1667941163
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_109
timestamp 1667941163
transform 1 0 11132 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_121
timestamp 1667941163
transform 1 0 12236 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_133
timestamp 1667941163
transform 1 0 13340 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_139
timestamp 1667941163
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_141
timestamp 1667941163
transform 1 0 14076 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_153
timestamp 1667941163
transform 1 0 15180 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_18_165
timestamp 1667941163
transform 1 0 16284 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_172
timestamp 1667941163
transform 1 0 16928 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_179
timestamp 1667941163
transform 1 0 17572 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_191
timestamp 1667941163
transform 1 0 18676 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_195
timestamp 1667941163
transform 1 0 19044 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_197
timestamp 1667941163
transform 1 0 19228 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_209
timestamp 1667941163
transform 1 0 20332 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_215
timestamp 1667941163
transform 1 0 20884 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_220
timestamp 1667941163
transform 1 0 21344 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_224
timestamp 1667941163
transform 1 0 21712 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_228
timestamp 1667941163
transform 1 0 22080 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_240
timestamp 1667941163
transform 1 0 23184 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_253
timestamp 1667941163
transform 1 0 24380 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_265
timestamp 1667941163
transform 1 0 25484 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_273
timestamp 1667941163
transform 1 0 26220 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_297
timestamp 1667941163
transform 1 0 28428 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_3
timestamp 1667941163
transform 1 0 1380 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_7
timestamp 1667941163
transform 1 0 1748 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_11
timestamp 1667941163
transform 1 0 2116 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_23
timestamp 1667941163
transform 1 0 3220 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_35
timestamp 1667941163
transform 1 0 4324 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_47
timestamp 1667941163
transform 1 0 5428 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1667941163
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_57
timestamp 1667941163
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_69
timestamp 1667941163
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_81
timestamp 1667941163
transform 1 0 8556 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_93
timestamp 1667941163
transform 1 0 9660 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_105
timestamp 1667941163
transform 1 0 10764 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1667941163
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_113
timestamp 1667941163
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_125
timestamp 1667941163
transform 1 0 12604 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_137
timestamp 1667941163
transform 1 0 13708 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_149
timestamp 1667941163
transform 1 0 14812 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_161
timestamp 1667941163
transform 1 0 15916 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_167
timestamp 1667941163
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_169
timestamp 1667941163
transform 1 0 16652 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_177
timestamp 1667941163
transform 1 0 17388 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_185
timestamp 1667941163
transform 1 0 18124 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_192
timestamp 1667941163
transform 1 0 18768 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_199
timestamp 1667941163
transform 1 0 19412 0 -1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_19_212
timestamp 1667941163
transform 1 0 20608 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_225
timestamp 1667941163
transform 1 0 21804 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_19_238
timestamp 1667941163
transform 1 0 23000 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_247
timestamp 1667941163
transform 1 0 23828 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_259
timestamp 1667941163
transform 1 0 24932 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_267
timestamp 1667941163
transform 1 0 25668 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_278
timestamp 1667941163
transform 1 0 26680 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_281
timestamp 1667941163
transform 1 0 26956 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_287
timestamp 1667941163
transform 1 0 27508 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_294
timestamp 1667941163
transform 1 0 28152 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_298
timestamp 1667941163
transform 1 0 28520 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_3
timestamp 1667941163
transform 1 0 1380 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_26
timestamp 1667941163
transform 1 0 3496 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_29
timestamp 1667941163
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_41
timestamp 1667941163
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_53
timestamp 1667941163
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_65
timestamp 1667941163
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_77
timestamp 1667941163
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1667941163
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_85
timestamp 1667941163
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_97
timestamp 1667941163
transform 1 0 10028 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_109
timestamp 1667941163
transform 1 0 11132 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_121
timestamp 1667941163
transform 1 0 12236 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_133
timestamp 1667941163
transform 1 0 13340 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_139
timestamp 1667941163
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_141
timestamp 1667941163
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_153
timestamp 1667941163
transform 1 0 15180 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_165
timestamp 1667941163
transform 1 0 16284 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_177
timestamp 1667941163
transform 1 0 17388 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_20_190
timestamp 1667941163
transform 1 0 18584 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_20_197
timestamp 1667941163
transform 1 0 19228 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_203
timestamp 1667941163
transform 1 0 19780 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_213
timestamp 1667941163
transform 1 0 20700 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_226
timestamp 1667941163
transform 1 0 21896 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_238
timestamp 1667941163
transform 1 0 23000 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_20_249
timestamp 1667941163
transform 1 0 24012 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_253
timestamp 1667941163
transform 1 0 24380 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_20_260
timestamp 1667941163
transform 1 0 25024 0 1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_20_271
timestamp 1667941163
transform 1 0 26036 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_283
timestamp 1667941163
transform 1 0 27140 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_295
timestamp 1667941163
transform 1 0 28244 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_3
timestamp 1667941163
transform 1 0 1380 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_21_14
timestamp 1667941163
transform 1 0 2392 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_21
timestamp 1667941163
transform 1 0 3036 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_28
timestamp 1667941163
transform 1 0 3680 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_40
timestamp 1667941163
transform 1 0 4784 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_52
timestamp 1667941163
transform 1 0 5888 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_57
timestamp 1667941163
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_69
timestamp 1667941163
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_81
timestamp 1667941163
transform 1 0 8556 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_93
timestamp 1667941163
transform 1 0 9660 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_105
timestamp 1667941163
transform 1 0 10764 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 1667941163
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_113
timestamp 1667941163
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_125
timestamp 1667941163
transform 1 0 12604 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_137
timestamp 1667941163
transform 1 0 13708 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_149
timestamp 1667941163
transform 1 0 14812 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_161
timestamp 1667941163
transform 1 0 15916 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_166
timestamp 1667941163
transform 1 0 16376 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_169
timestamp 1667941163
transform 1 0 16652 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_177
timestamp 1667941163
transform 1 0 17388 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_181
timestamp 1667941163
transform 1 0 17756 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_185
timestamp 1667941163
transform 1 0 18124 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_192
timestamp 1667941163
transform 1 0 18768 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_198
timestamp 1667941163
transform 1 0 19320 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_204
timestamp 1667941163
transform 1 0 19872 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_211
timestamp 1667941163
transform 1 0 20516 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_21_223
timestamp 1667941163
transform 1 0 21620 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_225
timestamp 1667941163
transform 1 0 21804 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_233
timestamp 1667941163
transform 1 0 22540 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_242
timestamp 1667941163
transform 1 0 23368 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_251
timestamp 1667941163
transform 1 0 24196 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_258
timestamp 1667941163
transform 1 0 24840 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_21_269
timestamp 1667941163
transform 1 0 25852 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_277
timestamp 1667941163
transform 1 0 26588 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_21_281
timestamp 1667941163
transform 1 0 26956 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_289
timestamp 1667941163
transform 1 0 27692 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_294
timestamp 1667941163
transform 1 0 28152 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_298
timestamp 1667941163
transform 1 0 28520 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_3
timestamp 1667941163
transform 1 0 1380 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_26
timestamp 1667941163
transform 1 0 3496 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_29
timestamp 1667941163
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_41
timestamp 1667941163
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_53
timestamp 1667941163
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_65
timestamp 1667941163
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_77
timestamp 1667941163
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1667941163
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_85
timestamp 1667941163
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_97
timestamp 1667941163
transform 1 0 10028 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_109
timestamp 1667941163
transform 1 0 11132 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_121
timestamp 1667941163
transform 1 0 12236 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_133
timestamp 1667941163
transform 1 0 13340 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_139
timestamp 1667941163
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_141
timestamp 1667941163
transform 1 0 14076 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_153
timestamp 1667941163
transform 1 0 15180 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_161
timestamp 1667941163
transform 1 0 15916 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_167
timestamp 1667941163
transform 1 0 16468 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_176
timestamp 1667941163
transform 1 0 17296 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_22_183
timestamp 1667941163
transform 1 0 17940 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_195
timestamp 1667941163
transform 1 0 19044 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_197
timestamp 1667941163
transform 1 0 19228 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_202
timestamp 1667941163
transform 1 0 19688 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_214
timestamp 1667941163
transform 1 0 20792 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_226
timestamp 1667941163
transform 1 0 21896 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_238
timestamp 1667941163
transform 1 0 23000 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_250
timestamp 1667941163
transform 1 0 24104 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_253
timestamp 1667941163
transform 1 0 24380 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_272
timestamp 1667941163
transform 1 0 26128 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_297
timestamp 1667941163
transform 1 0 28428 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_3
timestamp 1667941163
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_15
timestamp 1667941163
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_27
timestamp 1667941163
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_39
timestamp 1667941163
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_51
timestamp 1667941163
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1667941163
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_57
timestamp 1667941163
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_69
timestamp 1667941163
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_81
timestamp 1667941163
transform 1 0 8556 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_93
timestamp 1667941163
transform 1 0 9660 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_105
timestamp 1667941163
transform 1 0 10764 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp 1667941163
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_113
timestamp 1667941163
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_125
timestamp 1667941163
transform 1 0 12604 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_137
timestamp 1667941163
transform 1 0 13708 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_149
timestamp 1667941163
transform 1 0 14812 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_161
timestamp 1667941163
transform 1 0 15916 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_167
timestamp 1667941163
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_169
timestamp 1667941163
transform 1 0 16652 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_187
timestamp 1667941163
transform 1 0 18308 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_195
timestamp 1667941163
transform 1 0 19044 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_213
timestamp 1667941163
transform 1 0 20700 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_221
timestamp 1667941163
transform 1 0 21436 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_225
timestamp 1667941163
transform 1 0 21804 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_236
timestamp 1667941163
transform 1 0 22816 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_256
timestamp 1667941163
transform 1 0 24656 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_276
timestamp 1667941163
transform 1 0 26496 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_281
timestamp 1667941163
transform 1 0 26956 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_23_292
timestamp 1667941163
transform 1 0 27968 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_298
timestamp 1667941163
transform 1 0 28520 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_3
timestamp 1667941163
transform 1 0 1380 0 1 15232
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_24_14
timestamp 1667941163
transform 1 0 2392 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_24_26
timestamp 1667941163
transform 1 0 3496 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_29
timestamp 1667941163
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_41
timestamp 1667941163
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_53
timestamp 1667941163
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_65
timestamp 1667941163
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_77
timestamp 1667941163
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1667941163
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_85
timestamp 1667941163
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_97
timestamp 1667941163
transform 1 0 10028 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_103
timestamp 1667941163
transform 1 0 10580 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_107
timestamp 1667941163
transform 1 0 10948 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_132
timestamp 1667941163
transform 1 0 13248 0 1 15232
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_24_141
timestamp 1667941163
transform 1 0 14076 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_153
timestamp 1667941163
transform 1 0 15180 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_165
timestamp 1667941163
transform 1 0 16284 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_173
timestamp 1667941163
transform 1 0 17020 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_191
timestamp 1667941163
transform 1 0 18676 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_195
timestamp 1667941163
transform 1 0 19044 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_197
timestamp 1667941163
transform 1 0 19228 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_215
timestamp 1667941163
transform 1 0 20884 0 1 15232
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_24_239
timestamp 1667941163
transform 1 0 23092 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_251
timestamp 1667941163
transform 1 0 24196 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_253
timestamp 1667941163
transform 1 0 24380 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_268
timestamp 1667941163
transform 1 0 25760 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_288
timestamp 1667941163
transform 1 0 27600 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_295
timestamp 1667941163
transform 1 0 28244 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_25_3
timestamp 1667941163
transform 1 0 1380 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_25_27
timestamp 1667941163
transform 1 0 3588 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_39
timestamp 1667941163
transform 1 0 4692 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_51
timestamp 1667941163
transform 1 0 5796 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_55
timestamp 1667941163
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_57
timestamp 1667941163
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_69
timestamp 1667941163
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_81
timestamp 1667941163
transform 1 0 8556 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_93
timestamp 1667941163
transform 1 0 9660 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_105
timestamp 1667941163
transform 1 0 10764 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp 1667941163
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_113
timestamp 1667941163
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_125
timestamp 1667941163
transform 1 0 12604 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_137
timestamp 1667941163
transform 1 0 13708 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_149
timestamp 1667941163
transform 1 0 14812 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_161
timestamp 1667941163
transform 1 0 15916 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_167
timestamp 1667941163
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_169
timestamp 1667941163
transform 1 0 16652 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_187
timestamp 1667941163
transform 1 0 18308 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_199
timestamp 1667941163
transform 1 0 19412 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_207
timestamp 1667941163
transform 1 0 20148 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_213
timestamp 1667941163
transform 1 0 20700 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_222
timestamp 1667941163
transform 1 0 21528 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_225
timestamp 1667941163
transform 1 0 21804 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_237
timestamp 1667941163
transform 1 0 22908 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_249
timestamp 1667941163
transform 1 0 24012 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_261
timestamp 1667941163
transform 1 0 25116 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_269
timestamp 1667941163
transform 1 0 25852 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_276
timestamp 1667941163
transform 1 0 26496 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_281
timestamp 1667941163
transform 1 0 26956 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_286
timestamp 1667941163
transform 1 0 27416 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_297
timestamp 1667941163
transform 1 0 28428 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_3
timestamp 1667941163
transform 1 0 1380 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_26_10
timestamp 1667941163
transform 1 0 2024 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_22
timestamp 1667941163
transform 1 0 3128 0 1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_26_29
timestamp 1667941163
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_41
timestamp 1667941163
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_53
timestamp 1667941163
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_65
timestamp 1667941163
transform 1 0 7084 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_77
timestamp 1667941163
transform 1 0 8188 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 1667941163
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_85
timestamp 1667941163
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_97
timestamp 1667941163
transform 1 0 10028 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_109
timestamp 1667941163
transform 1 0 11132 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_121
timestamp 1667941163
transform 1 0 12236 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_133
timestamp 1667941163
transform 1 0 13340 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_139
timestamp 1667941163
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_141
timestamp 1667941163
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_153
timestamp 1667941163
transform 1 0 15180 0 1 16320
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_26_166
timestamp 1667941163
transform 1 0 16376 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_178
timestamp 1667941163
transform 1 0 17480 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_190
timestamp 1667941163
transform 1 0 18584 0 1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_26_197
timestamp 1667941163
transform 1 0 19228 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_26_209
timestamp 1667941163
transform 1 0 20332 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_26_228
timestamp 1667941163
transform 1 0 22080 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_236
timestamp 1667941163
transform 1 0 22816 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_26_246
timestamp 1667941163
transform 1 0 23736 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_26_253
timestamp 1667941163
transform 1 0 24380 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_262
timestamp 1667941163
transform 1 0 25208 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_272
timestamp 1667941163
transform 1 0 26128 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_297
timestamp 1667941163
transform 1 0 28428 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_3
timestamp 1667941163
transform 1 0 1380 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_9
timestamp 1667941163
transform 1 0 1932 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_27_16
timestamp 1667941163
transform 1 0 2576 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_28
timestamp 1667941163
transform 1 0 3680 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_40
timestamp 1667941163
transform 1 0 4784 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_52
timestamp 1667941163
transform 1 0 5888 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_27_57
timestamp 1667941163
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_69
timestamp 1667941163
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_81
timestamp 1667941163
transform 1 0 8556 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_93
timestamp 1667941163
transform 1 0 9660 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_105
timestamp 1667941163
transform 1 0 10764 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_111
timestamp 1667941163
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_113
timestamp 1667941163
transform 1 0 11500 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_125
timestamp 1667941163
transform 1 0 12604 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_137
timestamp 1667941163
transform 1 0 13708 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_27_148
timestamp 1667941163
transform 1 0 14720 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_156
timestamp 1667941163
transform 1 0 15456 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_164
timestamp 1667941163
transform 1 0 16192 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_27_169
timestamp 1667941163
transform 1 0 16652 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_181
timestamp 1667941163
transform 1 0 17756 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_200
timestamp 1667941163
transform 1 0 19504 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_213
timestamp 1667941163
transform 1 0 20700 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_221
timestamp 1667941163
transform 1 0 21436 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_225
timestamp 1667941163
transform 1 0 21804 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_236
timestamp 1667941163
transform 1 0 22816 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_248
timestamp 1667941163
transform 1 0 23920 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_266
timestamp 1667941163
transform 1 0 25576 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_270
timestamp 1667941163
transform 1 0 25944 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_27_274
timestamp 1667941163
transform 1 0 26312 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_27_281
timestamp 1667941163
transform 1 0 26956 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_287
timestamp 1667941163
transform 1 0 27508 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_294
timestamp 1667941163
transform 1 0 28152 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_298
timestamp 1667941163
transform 1 0 28520 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_3
timestamp 1667941163
transform 1 0 1380 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_26
timestamp 1667941163
transform 1 0 3496 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_29
timestamp 1667941163
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_41
timestamp 1667941163
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_53
timestamp 1667941163
transform 1 0 5980 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_65
timestamp 1667941163
transform 1 0 7084 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_77
timestamp 1667941163
transform 1 0 8188 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_83
timestamp 1667941163
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_85
timestamp 1667941163
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_97
timestamp 1667941163
transform 1 0 10028 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_109
timestamp 1667941163
transform 1 0 11132 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_121
timestamp 1667941163
transform 1 0 12236 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_28_133
timestamp 1667941163
transform 1 0 13340 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_138
timestamp 1667941163
transform 1 0 13800 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_141
timestamp 1667941163
transform 1 0 14076 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_28_150
timestamp 1667941163
transform 1 0 14904 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_28_158
timestamp 1667941163
transform 1 0 15640 0 1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_28_166
timestamp 1667941163
transform 1 0 16376 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_178
timestamp 1667941163
transform 1 0 17480 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_28_186
timestamp 1667941163
transform 1 0 18216 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_194
timestamp 1667941163
transform 1 0 18952 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_197
timestamp 1667941163
transform 1 0 19228 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_209
timestamp 1667941163
transform 1 0 20332 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_213
timestamp 1667941163
transform 1 0 20700 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_234
timestamp 1667941163
transform 1 0 22632 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_245
timestamp 1667941163
transform 1 0 23644 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_251
timestamp 1667941163
transform 1 0 24196 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_253
timestamp 1667941163
transform 1 0 24380 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_260
timestamp 1667941163
transform 1 0 25024 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_272
timestamp 1667941163
transform 1 0 26128 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_297
timestamp 1667941163
transform 1 0 28428 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_3
timestamp 1667941163
transform 1 0 1380 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_8
timestamp 1667941163
transform 1 0 1840 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_20
timestamp 1667941163
transform 1 0 2944 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_32
timestamp 1667941163
transform 1 0 4048 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_44
timestamp 1667941163
transform 1 0 5152 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_57
timestamp 1667941163
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_69
timestamp 1667941163
transform 1 0 7452 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_81
timestamp 1667941163
transform 1 0 8556 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_93
timestamp 1667941163
transform 1 0 9660 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_105
timestamp 1667941163
transform 1 0 10764 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_111
timestamp 1667941163
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_113
timestamp 1667941163
transform 1 0 11500 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_29_130
timestamp 1667941163
transform 1 0 13064 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_142
timestamp 1667941163
transform 1 0 14168 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_150
timestamp 1667941163
transform 1 0 14904 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_158
timestamp 1667941163
transform 1 0 15640 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_166
timestamp 1667941163
transform 1 0 16376 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_169
timestamp 1667941163
transform 1 0 16652 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_29_176
timestamp 1667941163
transform 1 0 17296 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_184
timestamp 1667941163
transform 1 0 18032 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_29_206
timestamp 1667941163
transform 1 0 20056 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_214
timestamp 1667941163
transform 1 0 20792 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_220
timestamp 1667941163
transform 1 0 21344 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_225
timestamp 1667941163
transform 1 0 21804 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_236
timestamp 1667941163
transform 1 0 22816 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_246
timestamp 1667941163
transform 1 0 23736 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_29_254
timestamp 1667941163
transform 1 0 24472 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_260
timestamp 1667941163
transform 1 0 25024 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_29_277
timestamp 1667941163
transform 1 0 26588 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_281
timestamp 1667941163
transform 1 0 26956 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_287
timestamp 1667941163
transform 1 0 27508 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_294
timestamp 1667941163
transform 1 0 28152 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_298
timestamp 1667941163
transform 1 0 28520 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_3
timestamp 1667941163
transform 1 0 1380 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_10
timestamp 1667941163
transform 1 0 2024 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_17
timestamp 1667941163
transform 1 0 2668 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_30_25
timestamp 1667941163
transform 1 0 3404 0 1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_30_29
timestamp 1667941163
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_41
timestamp 1667941163
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_53
timestamp 1667941163
transform 1 0 5980 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_65
timestamp 1667941163
transform 1 0 7084 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_77
timestamp 1667941163
transform 1 0 8188 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_83
timestamp 1667941163
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_85
timestamp 1667941163
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_97
timestamp 1667941163
transform 1 0 10028 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_109
timestamp 1667941163
transform 1 0 11132 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_121
timestamp 1667941163
transform 1 0 12236 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_125
timestamp 1667941163
transform 1 0 12604 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_129
timestamp 1667941163
transform 1 0 12972 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_136
timestamp 1667941163
transform 1 0 13616 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_141
timestamp 1667941163
transform 1 0 14076 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_30_148
timestamp 1667941163
transform 1 0 14720 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_156
timestamp 1667941163
transform 1 0 15456 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_165
timestamp 1667941163
transform 1 0 16284 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_185
timestamp 1667941163
transform 1 0 18124 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_192
timestamp 1667941163
transform 1 0 18768 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_197
timestamp 1667941163
transform 1 0 19228 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_30_208
timestamp 1667941163
transform 1 0 20240 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_30_230
timestamp 1667941163
transform 1 0 22264 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_236
timestamp 1667941163
transform 1 0 22816 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_241
timestamp 1667941163
transform 1 0 23276 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_30_249
timestamp 1667941163
transform 1 0 24012 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_253
timestamp 1667941163
transform 1 0 24380 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_30_262
timestamp 1667941163
transform 1 0 25208 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_268
timestamp 1667941163
transform 1 0 25760 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_272
timestamp 1667941163
transform 1 0 26128 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_297
timestamp 1667941163
transform 1 0 28428 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_3
timestamp 1667941163
transform 1 0 1380 0 -1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_31_27
timestamp 1667941163
transform 1 0 3588 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_39
timestamp 1667941163
transform 1 0 4692 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_51
timestamp 1667941163
transform 1 0 5796 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_55
timestamp 1667941163
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_57
timestamp 1667941163
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_69
timestamp 1667941163
transform 1 0 7452 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_81
timestamp 1667941163
transform 1 0 8556 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_93
timestamp 1667941163
transform 1 0 9660 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_105
timestamp 1667941163
transform 1 0 10764 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_111
timestamp 1667941163
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_113
timestamp 1667941163
transform 1 0 11500 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_121
timestamp 1667941163
transform 1 0 12236 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_31_129
timestamp 1667941163
transform 1 0 12972 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_31_140
timestamp 1667941163
transform 1 0 13984 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_147
timestamp 1667941163
transform 1 0 14628 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_159
timestamp 1667941163
transform 1 0 15732 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_166
timestamp 1667941163
transform 1 0 16376 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_169
timestamp 1667941163
transform 1 0 16652 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_31_188
timestamp 1667941163
transform 1 0 18400 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_196
timestamp 1667941163
transform 1 0 19136 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_206
timestamp 1667941163
transform 1 0 20056 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_214
timestamp 1667941163
transform 1 0 20792 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_219
timestamp 1667941163
transform 1 0 21252 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_223
timestamp 1667941163
transform 1 0 21620 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_225
timestamp 1667941163
transform 1 0 21804 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_237
timestamp 1667941163
transform 1 0 22908 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_249
timestamp 1667941163
transform 1 0 24012 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_261
timestamp 1667941163
transform 1 0 25116 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_273
timestamp 1667941163
transform 1 0 26220 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_279
timestamp 1667941163
transform 1 0 26772 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_281
timestamp 1667941163
transform 1 0 26956 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_31_292
timestamp 1667941163
transform 1 0 27968 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_298
timestamp 1667941163
transform 1 0 28520 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_3
timestamp 1667941163
transform 1 0 1380 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_26
timestamp 1667941163
transform 1 0 3496 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_29
timestamp 1667941163
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_41
timestamp 1667941163
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_53
timestamp 1667941163
transform 1 0 5980 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_65
timestamp 1667941163
transform 1 0 7084 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_77
timestamp 1667941163
transform 1 0 8188 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_83
timestamp 1667941163
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_85
timestamp 1667941163
transform 1 0 8924 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_97
timestamp 1667941163
transform 1 0 10028 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_109
timestamp 1667941163
transform 1 0 11132 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_121
timestamp 1667941163
transform 1 0 12236 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_32_129
timestamp 1667941163
transform 1 0 12972 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_136
timestamp 1667941163
transform 1 0 13616 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_141
timestamp 1667941163
transform 1 0 14076 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_32_153
timestamp 1667941163
transform 1 0 15180 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_161
timestamp 1667941163
transform 1 0 15916 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_169
timestamp 1667941163
transform 1 0 16652 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_173
timestamp 1667941163
transform 1 0 17020 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_185
timestamp 1667941163
transform 1 0 18124 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_32_193
timestamp 1667941163
transform 1 0 18860 0 1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_32_197
timestamp 1667941163
transform 1 0 19228 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_209
timestamp 1667941163
transform 1 0 20332 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_221
timestamp 1667941163
transform 1 0 21436 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_233
timestamp 1667941163
transform 1 0 22540 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_245
timestamp 1667941163
transform 1 0 23644 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_251
timestamp 1667941163
transform 1 0 24196 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_253
timestamp 1667941163
transform 1 0 24380 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_32_262
timestamp 1667941163
transform 1 0 25208 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_32_285
timestamp 1667941163
transform 1 0 27324 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_32_294
timestamp 1667941163
transform 1 0 28152 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_298
timestamp 1667941163
transform 1 0 28520 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_33_3
timestamp 1667941163
transform 1 0 1380 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_33_9
timestamp 1667941163
transform 1 0 1932 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_16
timestamp 1667941163
transform 1 0 2576 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_28
timestamp 1667941163
transform 1 0 3680 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_40
timestamp 1667941163
transform 1 0 4784 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_52
timestamp 1667941163
transform 1 0 5888 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_57
timestamp 1667941163
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_69
timestamp 1667941163
transform 1 0 7452 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_81
timestamp 1667941163
transform 1 0 8556 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_93
timestamp 1667941163
transform 1 0 9660 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_105
timestamp 1667941163
transform 1 0 10764 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_111
timestamp 1667941163
transform 1 0 11316 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_113
timestamp 1667941163
transform 1 0 11500 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_131
timestamp 1667941163
transform 1 0 13156 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_143
timestamp 1667941163
transform 1 0 14260 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_153
timestamp 1667941163
transform 1 0 15180 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_33_165
timestamp 1667941163
transform 1 0 16284 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_33_169
timestamp 1667941163
transform 1 0 16652 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_181
timestamp 1667941163
transform 1 0 17756 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_189
timestamp 1667941163
transform 1 0 18492 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_33_194
timestamp 1667941163
transform 1 0 18952 0 -1 20672
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_33_209
timestamp 1667941163
transform 1 0 20332 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_33_221
timestamp 1667941163
transform 1 0 21436 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_33_225
timestamp 1667941163
transform 1 0 21804 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_229
timestamp 1667941163
transform 1 0 22172 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_236
timestamp 1667941163
transform 1 0 22816 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_33_251
timestamp 1667941163
transform 1 0 24196 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_259
timestamp 1667941163
transform 1 0 24932 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_268
timestamp 1667941163
transform 1 0 25760 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_281
timestamp 1667941163
transform 1 0 26956 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_285
timestamp 1667941163
transform 1 0 27324 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_289
timestamp 1667941163
transform 1 0 27692 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_33_296
timestamp 1667941163
transform 1 0 28336 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_34_3
timestamp 1667941163
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_15
timestamp 1667941163
transform 1 0 2484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 1667941163
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_29
timestamp 1667941163
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_41
timestamp 1667941163
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_53
timestamp 1667941163
transform 1 0 5980 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_65
timestamp 1667941163
transform 1 0 7084 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_77
timestamp 1667941163
transform 1 0 8188 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_83
timestamp 1667941163
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_85
timestamp 1667941163
transform 1 0 8924 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_97
timestamp 1667941163
transform 1 0 10028 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_109
timestamp 1667941163
transform 1 0 11132 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_121
timestamp 1667941163
transform 1 0 12236 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_133
timestamp 1667941163
transform 1 0 13340 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_139
timestamp 1667941163
transform 1 0 13892 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_34_141
timestamp 1667941163
transform 1 0 14076 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_149
timestamp 1667941163
transform 1 0 14812 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_156
timestamp 1667941163
transform 1 0 15456 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_160
timestamp 1667941163
transform 1 0 15824 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_166
timestamp 1667941163
transform 1 0 16376 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_178
timestamp 1667941163
transform 1 0 17480 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_34_186
timestamp 1667941163
transform 1 0 18216 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_34_194
timestamp 1667941163
transform 1 0 18952 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_197
timestamp 1667941163
transform 1 0 19228 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_201
timestamp 1667941163
transform 1 0 19596 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_34_218
timestamp 1667941163
transform 1 0 21160 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_224
timestamp 1667941163
transform 1 0 21712 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_34_241
timestamp 1667941163
transform 1 0 23276 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_34_249
timestamp 1667941163
transform 1 0 24012 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_34_253
timestamp 1667941163
transform 1 0 24380 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_34_261
timestamp 1667941163
transform 1 0 25116 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_34_272
timestamp 1667941163
transform 1 0 26128 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_297
timestamp 1667941163
transform 1 0 28428 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_3
timestamp 1667941163
transform 1 0 1380 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_15
timestamp 1667941163
transform 1 0 2484 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_27
timestamp 1667941163
transform 1 0 3588 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_39
timestamp 1667941163
transform 1 0 4692 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_51
timestamp 1667941163
transform 1 0 5796 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_55
timestamp 1667941163
transform 1 0 6164 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_57
timestamp 1667941163
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_69
timestamp 1667941163
transform 1 0 7452 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_81
timestamp 1667941163
transform 1 0 8556 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_93
timestamp 1667941163
transform 1 0 9660 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_105
timestamp 1667941163
transform 1 0 10764 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_111
timestamp 1667941163
transform 1 0 11316 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_113
timestamp 1667941163
transform 1 0 11500 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_125
timestamp 1667941163
transform 1 0 12604 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_137
timestamp 1667941163
transform 1 0 13708 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_149
timestamp 1667941163
transform 1 0 14812 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_166
timestamp 1667941163
transform 1 0 16376 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_169
timestamp 1667941163
transform 1 0 16652 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_187
timestamp 1667941163
transform 1 0 18308 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_207
timestamp 1667941163
transform 1 0 20148 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_213
timestamp 1667941163
transform 1 0 20700 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_220
timestamp 1667941163
transform 1 0 21344 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_225
timestamp 1667941163
transform 1 0 21804 0 -1 21760
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_35_237
timestamp 1667941163
transform 1 0 22908 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_249
timestamp 1667941163
transform 1 0 24012 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_264
timestamp 1667941163
transform 1 0 25392 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_276
timestamp 1667941163
transform 1 0 26496 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_281
timestamp 1667941163
transform 1 0 26956 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_285
timestamp 1667941163
transform 1 0 27324 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_289
timestamp 1667941163
transform 1 0 27692 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_35_296
timestamp 1667941163
transform 1 0 28336 0 -1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_36_3
timestamp 1667941163
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_15
timestamp 1667941163
transform 1 0 2484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 1667941163
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_29
timestamp 1667941163
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_41
timestamp 1667941163
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_53
timestamp 1667941163
transform 1 0 5980 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_65
timestamp 1667941163
transform 1 0 7084 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_77
timestamp 1667941163
transform 1 0 8188 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_83
timestamp 1667941163
transform 1 0 8740 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_85
timestamp 1667941163
transform 1 0 8924 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_97
timestamp 1667941163
transform 1 0 10028 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_109
timestamp 1667941163
transform 1 0 11132 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_121
timestamp 1667941163
transform 1 0 12236 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_133
timestamp 1667941163
transform 1 0 13340 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_139
timestamp 1667941163
transform 1 0 13892 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_141
timestamp 1667941163
transform 1 0 14076 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_153
timestamp 1667941163
transform 1 0 15180 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_36_164
timestamp 1667941163
transform 1 0 16192 0 1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_36_171
timestamp 1667941163
transform 1 0 16836 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_183
timestamp 1667941163
transform 1 0 17940 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_195
timestamp 1667941163
transform 1 0 19044 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_197
timestamp 1667941163
transform 1 0 19228 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_209
timestamp 1667941163
transform 1 0 20332 0 1 21760
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_36_221
timestamp 1667941163
transform 1 0 21436 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_36_233
timestamp 1667941163
transform 1 0 22540 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_240
timestamp 1667941163
transform 1 0 23184 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_244
timestamp 1667941163
transform 1 0 23552 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_36_249
timestamp 1667941163
transform 1 0 24012 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_36_253
timestamp 1667941163
transform 1 0 24380 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_36_263
timestamp 1667941163
transform 1 0 25300 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_275
timestamp 1667941163
transform 1 0 26404 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_297
timestamp 1667941163
transform 1 0 28428 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_3
timestamp 1667941163
transform 1 0 1380 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_15
timestamp 1667941163
transform 1 0 2484 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_27
timestamp 1667941163
transform 1 0 3588 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_39
timestamp 1667941163
transform 1 0 4692 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_51
timestamp 1667941163
transform 1 0 5796 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_55
timestamp 1667941163
transform 1 0 6164 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_57
timestamp 1667941163
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_69
timestamp 1667941163
transform 1 0 7452 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_81
timestamp 1667941163
transform 1 0 8556 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_93
timestamp 1667941163
transform 1 0 9660 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_105
timestamp 1667941163
transform 1 0 10764 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_111
timestamp 1667941163
transform 1 0 11316 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_113
timestamp 1667941163
transform 1 0 11500 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_125
timestamp 1667941163
transform 1 0 12604 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_137
timestamp 1667941163
transform 1 0 13708 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_149
timestamp 1667941163
transform 1 0 14812 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_37_164
timestamp 1667941163
transform 1 0 16192 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_169
timestamp 1667941163
transform 1 0 16652 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_187
timestamp 1667941163
transform 1 0 18308 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_199
timestamp 1667941163
transform 1 0 19412 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_211
timestamp 1667941163
transform 1 0 20516 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_37_223
timestamp 1667941163
transform 1 0 21620 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_225
timestamp 1667941163
transform 1 0 21804 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_232
timestamp 1667941163
transform 1 0 22448 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_244
timestamp 1667941163
transform 1 0 23552 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_250
timestamp 1667941163
transform 1 0 24104 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_37_256
timestamp 1667941163
transform 1 0 24656 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_37_278
timestamp 1667941163
transform 1 0 26680 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_37_281
timestamp 1667941163
transform 1 0 26956 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_37_287
timestamp 1667941163
transform 1 0 27508 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_294
timestamp 1667941163
transform 1 0 28152 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_298
timestamp 1667941163
transform 1 0 28520 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_3
timestamp 1667941163
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_15
timestamp 1667941163
transform 1 0 2484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 1667941163
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_29
timestamp 1667941163
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_41
timestamp 1667941163
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_53
timestamp 1667941163
transform 1 0 5980 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_65
timestamp 1667941163
transform 1 0 7084 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_77
timestamp 1667941163
transform 1 0 8188 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_83
timestamp 1667941163
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_85
timestamp 1667941163
transform 1 0 8924 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_97
timestamp 1667941163
transform 1 0 10028 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_109
timestamp 1667941163
transform 1 0 11132 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_121
timestamp 1667941163
transform 1 0 12236 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_133
timestamp 1667941163
transform 1 0 13340 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_139
timestamp 1667941163
transform 1 0 13892 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_141
timestamp 1667941163
transform 1 0 14076 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_153
timestamp 1667941163
transform 1 0 15180 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_165
timestamp 1667941163
transform 1 0 16284 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_169
timestamp 1667941163
transform 1 0 16652 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_181
timestamp 1667941163
transform 1 0 17756 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_187
timestamp 1667941163
transform 1 0 18308 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_38_193
timestamp 1667941163
transform 1 0 18860 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_38_197
timestamp 1667941163
transform 1 0 19228 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_38_208
timestamp 1667941163
transform 1 0 20240 0 1 22848
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_38_222
timestamp 1667941163
transform 1 0 21528 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_234
timestamp 1667941163
transform 1 0 22632 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_246
timestamp 1667941163
transform 1 0 23736 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_38_253
timestamp 1667941163
transform 1 0 24380 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_261
timestamp 1667941163
transform 1 0 25116 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_38_270
timestamp 1667941163
transform 1 0 25944 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_38_297
timestamp 1667941163
transform 1 0 28428 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_39_3
timestamp 1667941163
transform 1 0 1380 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_15
timestamp 1667941163
transform 1 0 2484 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_27
timestamp 1667941163
transform 1 0 3588 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_39
timestamp 1667941163
transform 1 0 4692 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_51
timestamp 1667941163
transform 1 0 5796 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_55
timestamp 1667941163
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_57
timestamp 1667941163
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_69
timestamp 1667941163
transform 1 0 7452 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_81
timestamp 1667941163
transform 1 0 8556 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_93
timestamp 1667941163
transform 1 0 9660 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_105
timestamp 1667941163
transform 1 0 10764 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_111
timestamp 1667941163
transform 1 0 11316 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_113
timestamp 1667941163
transform 1 0 11500 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_125
timestamp 1667941163
transform 1 0 12604 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_137
timestamp 1667941163
transform 1 0 13708 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_149
timestamp 1667941163
transform 1 0 14812 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_161
timestamp 1667941163
transform 1 0 15916 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_167
timestamp 1667941163
transform 1 0 16468 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_169
timestamp 1667941163
transform 1 0 16652 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_39_176
timestamp 1667941163
transform 1 0 17296 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_184
timestamp 1667941163
transform 1 0 18032 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_202
timestamp 1667941163
transform 1 0 19688 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_222
timestamp 1667941163
transform 1 0 21528 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_225
timestamp 1667941163
transform 1 0 21804 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_232
timestamp 1667941163
transform 1 0 22448 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_244
timestamp 1667941163
transform 1 0 23552 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_39_252
timestamp 1667941163
transform 1 0 24288 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_39_260
timestamp 1667941163
transform 1 0 25024 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_269
timestamp 1667941163
transform 1 0 25852 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_278
timestamp 1667941163
transform 1 0 26680 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_39_281
timestamp 1667941163
transform 1 0 26956 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_39_287
timestamp 1667941163
transform 1 0 27508 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_294
timestamp 1667941163
transform 1 0 28152 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_298
timestamp 1667941163
transform 1 0 28520 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_3
timestamp 1667941163
transform 1 0 1380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_15
timestamp 1667941163
transform 1 0 2484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_27
timestamp 1667941163
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_29
timestamp 1667941163
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_41
timestamp 1667941163
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_53
timestamp 1667941163
transform 1 0 5980 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_65
timestamp 1667941163
transform 1 0 7084 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_77
timestamp 1667941163
transform 1 0 8188 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_83
timestamp 1667941163
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_85
timestamp 1667941163
transform 1 0 8924 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_97
timestamp 1667941163
transform 1 0 10028 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_109
timestamp 1667941163
transform 1 0 11132 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_121
timestamp 1667941163
transform 1 0 12236 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_133
timestamp 1667941163
transform 1 0 13340 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_139
timestamp 1667941163
transform 1 0 13892 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_141
timestamp 1667941163
transform 1 0 14076 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_153
timestamp 1667941163
transform 1 0 15180 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_166
timestamp 1667941163
transform 1 0 16376 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_186
timestamp 1667941163
transform 1 0 18216 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_40_193
timestamp 1667941163
transform 1 0 18860 0 1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_40_197
timestamp 1667941163
transform 1 0 19228 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_209
timestamp 1667941163
transform 1 0 20332 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_217
timestamp 1667941163
transform 1 0 21068 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_40_224
timestamp 1667941163
transform 1 0 21712 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_232
timestamp 1667941163
transform 1 0 22448 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_40_249
timestamp 1667941163
transform 1 0 24012 0 1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_40_253
timestamp 1667941163
transform 1 0 24380 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_265
timestamp 1667941163
transform 1 0 25484 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_40_273
timestamp 1667941163
transform 1 0 26220 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_40_297
timestamp 1667941163
transform 1 0 28428 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_41_3
timestamp 1667941163
transform 1 0 1380 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_15
timestamp 1667941163
transform 1 0 2484 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_27
timestamp 1667941163
transform 1 0 3588 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_39
timestamp 1667941163
transform 1 0 4692 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_51
timestamp 1667941163
transform 1 0 5796 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_55
timestamp 1667941163
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_57
timestamp 1667941163
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_69
timestamp 1667941163
transform 1 0 7452 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_81
timestamp 1667941163
transform 1 0 8556 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_93
timestamp 1667941163
transform 1 0 9660 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_105
timestamp 1667941163
transform 1 0 10764 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_111
timestamp 1667941163
transform 1 0 11316 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_113
timestamp 1667941163
transform 1 0 11500 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_125
timestamp 1667941163
transform 1 0 12604 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_137
timestamp 1667941163
transform 1 0 13708 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_149
timestamp 1667941163
transform 1 0 14812 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_161
timestamp 1667941163
transform 1 0 15916 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_167
timestamp 1667941163
transform 1 0 16468 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_41_169
timestamp 1667941163
transform 1 0 16652 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_41_174
timestamp 1667941163
transform 1 0 17112 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_186
timestamp 1667941163
transform 1 0 18216 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_198
timestamp 1667941163
transform 1 0 19320 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_210
timestamp 1667941163
transform 1 0 20424 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_41_222
timestamp 1667941163
transform 1 0 21528 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_41_225
timestamp 1667941163
transform 1 0 21804 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_41_236
timestamp 1667941163
transform 1 0 22816 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_247
timestamp 1667941163
transform 1 0 23828 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_41_256
timestamp 1667941163
transform 1 0 24656 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_41_270
timestamp 1667941163
transform 1 0 25944 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_278
timestamp 1667941163
transform 1 0 26680 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_281
timestamp 1667941163
transform 1 0 26956 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_289
timestamp 1667941163
transform 1 0 27692 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_41_296
timestamp 1667941163
transform 1 0 28336 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_42_3
timestamp 1667941163
transform 1 0 1380 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_8
timestamp 1667941163
transform 1 0 1840 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_12
timestamp 1667941163
transform 1 0 2208 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_16
timestamp 1667941163
transform 1 0 2576 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_29
timestamp 1667941163
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_41
timestamp 1667941163
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_53
timestamp 1667941163
transform 1 0 5980 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_65
timestamp 1667941163
transform 1 0 7084 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_77
timestamp 1667941163
transform 1 0 8188 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_83
timestamp 1667941163
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_85
timestamp 1667941163
transform 1 0 8924 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_97
timestamp 1667941163
transform 1 0 10028 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_109
timestamp 1667941163
transform 1 0 11132 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_121
timestamp 1667941163
transform 1 0 12236 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_133
timestamp 1667941163
transform 1 0 13340 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_139
timestamp 1667941163
transform 1 0 13892 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_141
timestamp 1667941163
transform 1 0 14076 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_153
timestamp 1667941163
transform 1 0 15180 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_161
timestamp 1667941163
transform 1 0 15916 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_168
timestamp 1667941163
transform 1 0 16560 0 1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_42_175
timestamp 1667941163
transform 1 0 17204 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_187
timestamp 1667941163
transform 1 0 18308 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_42_194
timestamp 1667941163
transform 1 0 18952 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_197
timestamp 1667941163
transform 1 0 19228 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_42_204
timestamp 1667941163
transform 1 0 19872 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_212
timestamp 1667941163
transform 1 0 20608 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_220
timestamp 1667941163
transform 1 0 21344 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_232
timestamp 1667941163
transform 1 0 22448 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_240
timestamp 1667941163
transform 1 0 23184 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_247
timestamp 1667941163
transform 1 0 23828 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_251
timestamp 1667941163
transform 1 0 24196 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_42_253
timestamp 1667941163
transform 1 0 24380 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_42_261
timestamp 1667941163
transform 1 0 25116 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_268
timestamp 1667941163
transform 1 0 25760 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_297
timestamp 1667941163
transform 1 0 28428 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_43_3
timestamp 1667941163
transform 1 0 1380 0 -1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_43_27
timestamp 1667941163
transform 1 0 3588 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_39
timestamp 1667941163
transform 1 0 4692 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_51
timestamp 1667941163
transform 1 0 5796 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_55
timestamp 1667941163
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_57
timestamp 1667941163
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_69
timestamp 1667941163
transform 1 0 7452 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_81
timestamp 1667941163
transform 1 0 8556 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_93
timestamp 1667941163
transform 1 0 9660 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_105
timestamp 1667941163
transform 1 0 10764 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_111
timestamp 1667941163
transform 1 0 11316 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_113
timestamp 1667941163
transform 1 0 11500 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_125
timestamp 1667941163
transform 1 0 12604 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_137
timestamp 1667941163
transform 1 0 13708 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_149
timestamp 1667941163
transform 1 0 14812 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_166
timestamp 1667941163
transform 1 0 16376 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_169
timestamp 1667941163
transform 1 0 16652 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_187
timestamp 1667941163
transform 1 0 18308 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_191
timestamp 1667941163
transform 1 0 18676 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_208
timestamp 1667941163
transform 1 0 20240 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_43_221
timestamp 1667941163
transform 1 0 21436 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_43_225
timestamp 1667941163
transform 1 0 21804 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_249
timestamp 1667941163
transform 1 0 24012 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_262
timestamp 1667941163
transform 1 0 25208 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_270
timestamp 1667941163
transform 1 0 25944 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_43_278
timestamp 1667941163
transform 1 0 26680 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_281
timestamp 1667941163
transform 1 0 26956 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_286
timestamp 1667941163
transform 1 0 27416 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_43_293
timestamp 1667941163
transform 1 0 28060 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_44_3
timestamp 1667941163
transform 1 0 1380 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_44_10
timestamp 1667941163
transform 1 0 2024 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_22
timestamp 1667941163
transform 1 0 3128 0 1 26112
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_44_29
timestamp 1667941163
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_41
timestamp 1667941163
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_53
timestamp 1667941163
transform 1 0 5980 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_65
timestamp 1667941163
transform 1 0 7084 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_77
timestamp 1667941163
transform 1 0 8188 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_83
timestamp 1667941163
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_85
timestamp 1667941163
transform 1 0 8924 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_97
timestamp 1667941163
transform 1 0 10028 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_109
timestamp 1667941163
transform 1 0 11132 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_121
timestamp 1667941163
transform 1 0 12236 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_133
timestamp 1667941163
transform 1 0 13340 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_139
timestamp 1667941163
transform 1 0 13892 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_141
timestamp 1667941163
transform 1 0 14076 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_153
timestamp 1667941163
transform 1 0 15180 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_165
timestamp 1667941163
transform 1 0 16284 0 1 26112
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_44_175
timestamp 1667941163
transform 1 0 17204 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_187
timestamp 1667941163
transform 1 0 18308 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_195
timestamp 1667941163
transform 1 0 19044 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_197
timestamp 1667941163
transform 1 0 19228 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_202
timestamp 1667941163
transform 1 0 19688 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_44_214
timestamp 1667941163
transform 1 0 20792 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_222
timestamp 1667941163
transform 1 0 21528 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_243
timestamp 1667941163
transform 1 0 23460 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_251
timestamp 1667941163
transform 1 0 24196 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_253
timestamp 1667941163
transform 1 0 24380 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_258
timestamp 1667941163
transform 1 0 24840 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_270
timestamp 1667941163
transform 1 0 25944 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_44_297
timestamp 1667941163
transform 1 0 28428 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_45_3
timestamp 1667941163
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_15
timestamp 1667941163
transform 1 0 2484 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_27
timestamp 1667941163
transform 1 0 3588 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_39
timestamp 1667941163
transform 1 0 4692 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_51
timestamp 1667941163
transform 1 0 5796 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_55
timestamp 1667941163
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_57
timestamp 1667941163
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_69
timestamp 1667941163
transform 1 0 7452 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_81
timestamp 1667941163
transform 1 0 8556 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_93
timestamp 1667941163
transform 1 0 9660 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_105
timestamp 1667941163
transform 1 0 10764 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_111
timestamp 1667941163
transform 1 0 11316 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_113
timestamp 1667941163
transform 1 0 11500 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_125
timestamp 1667941163
transform 1 0 12604 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_137
timestamp 1667941163
transform 1 0 13708 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_149
timestamp 1667941163
transform 1 0 14812 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_45_162
timestamp 1667941163
transform 1 0 16008 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_45_169
timestamp 1667941163
transform 1 0 16652 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_45_174
timestamp 1667941163
transform 1 0 17112 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_45_186
timestamp 1667941163
transform 1 0 18216 0 -1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_45_193
timestamp 1667941163
transform 1 0 18860 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_205
timestamp 1667941163
transform 1 0 19964 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_45_217
timestamp 1667941163
transform 1 0 21068 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_222
timestamp 1667941163
transform 1 0 21528 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_225
timestamp 1667941163
transform 1 0 21804 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_45_232
timestamp 1667941163
transform 1 0 22448 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_244
timestamp 1667941163
transform 1 0 23552 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_256
timestamp 1667941163
transform 1 0 24656 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_45_268
timestamp 1667941163
transform 1 0 25760 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_45_273
timestamp 1667941163
transform 1 0 26220 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_279
timestamp 1667941163
transform 1 0 26772 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_45_281
timestamp 1667941163
transform 1 0 26956 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_286
timestamp 1667941163
transform 1 0 27416 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_45_293
timestamp 1667941163
transform 1 0 28060 0 -1 27200
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_46_3
timestamp 1667941163
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_15
timestamp 1667941163
transform 1 0 2484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_27
timestamp 1667941163
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_29
timestamp 1667941163
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_41
timestamp 1667941163
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_53
timestamp 1667941163
transform 1 0 5980 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_65
timestamp 1667941163
transform 1 0 7084 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_77
timestamp 1667941163
transform 1 0 8188 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_83
timestamp 1667941163
transform 1 0 8740 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_85
timestamp 1667941163
transform 1 0 8924 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_97
timestamp 1667941163
transform 1 0 10028 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_109
timestamp 1667941163
transform 1 0 11132 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_121
timestamp 1667941163
transform 1 0 12236 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_133
timestamp 1667941163
transform 1 0 13340 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_139
timestamp 1667941163
transform 1 0 13892 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_141
timestamp 1667941163
transform 1 0 14076 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_162
timestamp 1667941163
transform 1 0 16008 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_168
timestamp 1667941163
transform 1 0 16560 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_46_185
timestamp 1667941163
transform 1 0 18124 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_46_193
timestamp 1667941163
transform 1 0 18860 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_46_197
timestamp 1667941163
transform 1 0 19228 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_46_221
timestamp 1667941163
transform 1 0 21436 0 1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_46_229
timestamp 1667941163
transform 1 0 22172 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_241
timestamp 1667941163
transform 1 0 23276 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_46_250
timestamp 1667941163
transform 1 0 24104 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_46_253
timestamp 1667941163
transform 1 0 24380 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_46_267
timestamp 1667941163
transform 1 0 25668 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_275
timestamp 1667941163
transform 1 0 26404 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_46_297
timestamp 1667941163
transform 1 0 28428 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_3
timestamp 1667941163
transform 1 0 1380 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_47_8
timestamp 1667941163
transform 1 0 1840 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_20
timestamp 1667941163
transform 1 0 2944 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_32
timestamp 1667941163
transform 1 0 4048 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_44
timestamp 1667941163
transform 1 0 5152 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_57
timestamp 1667941163
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_69
timestamp 1667941163
transform 1 0 7452 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_81
timestamp 1667941163
transform 1 0 8556 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_93
timestamp 1667941163
transform 1 0 9660 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_105
timestamp 1667941163
transform 1 0 10764 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_111
timestamp 1667941163
transform 1 0 11316 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_113
timestamp 1667941163
transform 1 0 11500 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_125
timestamp 1667941163
transform 1 0 12604 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_137
timestamp 1667941163
transform 1 0 13708 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_149
timestamp 1667941163
transform 1 0 14812 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_161
timestamp 1667941163
transform 1 0 15916 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_167
timestamp 1667941163
transform 1 0 16468 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_169
timestamp 1667941163
transform 1 0 16652 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_47_181
timestamp 1667941163
transform 1 0 17756 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_188
timestamp 1667941163
transform 1 0 18400 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_200
timestamp 1667941163
transform 1 0 19504 0 -1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_47_207
timestamp 1667941163
transform 1 0 20148 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_219
timestamp 1667941163
transform 1 0 21252 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_223
timestamp 1667941163
transform 1 0 21620 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_225
timestamp 1667941163
transform 1 0 21804 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_47_237
timestamp 1667941163
transform 1 0 22908 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_47_246
timestamp 1667941163
transform 1 0 23736 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_47_255
timestamp 1667941163
transform 1 0 24564 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_47_263
timestamp 1667941163
transform 1 0 25300 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_47_273
timestamp 1667941163
transform 1 0 26220 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_279
timestamp 1667941163
transform 1 0 26772 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_47_281
timestamp 1667941163
transform 1 0 26956 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_288
timestamp 1667941163
transform 1 0 27600 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_295
timestamp 1667941163
transform 1 0 28244 0 -1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_48_3
timestamp 1667941163
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_15
timestamp 1667941163
transform 1 0 2484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 1667941163
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_29
timestamp 1667941163
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_41
timestamp 1667941163
transform 1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_53
timestamp 1667941163
transform 1 0 5980 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_65
timestamp 1667941163
transform 1 0 7084 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_77
timestamp 1667941163
transform 1 0 8188 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_83
timestamp 1667941163
transform 1 0 8740 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_85
timestamp 1667941163
transform 1 0 8924 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_97
timestamp 1667941163
transform 1 0 10028 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_109
timestamp 1667941163
transform 1 0 11132 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_121
timestamp 1667941163
transform 1 0 12236 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_133
timestamp 1667941163
transform 1 0 13340 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_139
timestamp 1667941163
transform 1 0 13892 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_141
timestamp 1667941163
transform 1 0 14076 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_153
timestamp 1667941163
transform 1 0 15180 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_48_166
timestamp 1667941163
transform 1 0 16376 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_170
timestamp 1667941163
transform 1 0 16744 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_48_187
timestamp 1667941163
transform 1 0 18308 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_195
timestamp 1667941163
transform 1 0 19044 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_48_197
timestamp 1667941163
transform 1 0 19228 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_48_215
timestamp 1667941163
transform 1 0 20884 0 1 28288
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_48_225
timestamp 1667941163
transform 1 0 21804 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_237
timestamp 1667941163
transform 1 0 22908 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_48_249
timestamp 1667941163
transform 1 0 24012 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_48_253
timestamp 1667941163
transform 1 0 24380 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_48_263
timestamp 1667941163
transform 1 0 25300 0 1 28288
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_48_287
timestamp 1667941163
transform 1 0 27508 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_3
timestamp 1667941163
transform 1 0 1380 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_15
timestamp 1667941163
transform 1 0 2484 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_27
timestamp 1667941163
transform 1 0 3588 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_39
timestamp 1667941163
transform 1 0 4692 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_51
timestamp 1667941163
transform 1 0 5796 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_55
timestamp 1667941163
transform 1 0 6164 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_57
timestamp 1667941163
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_69
timestamp 1667941163
transform 1 0 7452 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_81
timestamp 1667941163
transform 1 0 8556 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_93
timestamp 1667941163
transform 1 0 9660 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_105
timestamp 1667941163
transform 1 0 10764 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_111
timestamp 1667941163
transform 1 0 11316 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_113
timestamp 1667941163
transform 1 0 11500 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_125
timestamp 1667941163
transform 1 0 12604 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_137
timestamp 1667941163
transform 1 0 13708 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_149
timestamp 1667941163
transform 1 0 14812 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_49_157
timestamp 1667941163
transform 1 0 15548 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_49_163
timestamp 1667941163
transform 1 0 16100 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_167
timestamp 1667941163
transform 1 0 16468 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_169
timestamp 1667941163
transform 1 0 16652 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_181
timestamp 1667941163
transform 1 0 17756 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_185
timestamp 1667941163
transform 1 0 18124 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_49_206
timestamp 1667941163
transform 1 0 20056 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_49_214
timestamp 1667941163
transform 1 0 20792 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_220
timestamp 1667941163
transform 1 0 21344 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_49_225
timestamp 1667941163
transform 1 0 21804 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_49_244
timestamp 1667941163
transform 1 0 23552 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_256
timestamp 1667941163
transform 1 0 24656 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_265
timestamp 1667941163
transform 1 0 25484 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_49_273
timestamp 1667941163
transform 1 0 26220 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_279
timestamp 1667941163
transform 1 0 26772 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_49_281
timestamp 1667941163
transform 1 0 26956 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_287
timestamp 1667941163
transform 1 0 27508 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_49_291
timestamp 1667941163
transform 1 0 27876 0 -1 29376
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_50_3
timestamp 1667941163
transform 1 0 1380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_15
timestamp 1667941163
transform 1 0 2484 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_27
timestamp 1667941163
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_29
timestamp 1667941163
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_41
timestamp 1667941163
transform 1 0 4876 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_53
timestamp 1667941163
transform 1 0 5980 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_65
timestamp 1667941163
transform 1 0 7084 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_77
timestamp 1667941163
transform 1 0 8188 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_83
timestamp 1667941163
transform 1 0 8740 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_85
timestamp 1667941163
transform 1 0 8924 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_97
timestamp 1667941163
transform 1 0 10028 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_109
timestamp 1667941163
transform 1 0 11132 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_121
timestamp 1667941163
transform 1 0 12236 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_133
timestamp 1667941163
transform 1 0 13340 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_139
timestamp 1667941163
transform 1 0 13892 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_141
timestamp 1667941163
transform 1 0 14076 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_153
timestamp 1667941163
transform 1 0 15180 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_159
timestamp 1667941163
transform 1 0 15732 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_163
timestamp 1667941163
transform 1 0 16100 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_167
timestamp 1667941163
transform 1 0 16468 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_50_171
timestamp 1667941163
transform 1 0 16836 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_50_182
timestamp 1667941163
transform 1 0 17848 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_192
timestamp 1667941163
transform 1 0 18768 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_50_197
timestamp 1667941163
transform 1 0 19228 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_50_202
timestamp 1667941163
transform 1 0 19688 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_210
timestamp 1667941163
transform 1 0 20424 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_230
timestamp 1667941163
transform 1 0 22264 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_238
timestamp 1667941163
transform 1 0 23000 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_50_246
timestamp 1667941163
transform 1 0 23736 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_50_253
timestamp 1667941163
transform 1 0 24380 0 1 29376
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_50_264
timestamp 1667941163
transform 1 0 25392 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_50_297
timestamp 1667941163
transform 1 0 28428 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_3
timestamp 1667941163
transform 1 0 1380 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_51_8
timestamp 1667941163
transform 1 0 1840 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_20
timestamp 1667941163
transform 1 0 2944 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_32
timestamp 1667941163
transform 1 0 4048 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_44
timestamp 1667941163
transform 1 0 5152 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_57
timestamp 1667941163
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_69
timestamp 1667941163
transform 1 0 7452 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_81
timestamp 1667941163
transform 1 0 8556 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_93
timestamp 1667941163
transform 1 0 9660 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_105
timestamp 1667941163
transform 1 0 10764 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_111
timestamp 1667941163
transform 1 0 11316 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_113
timestamp 1667941163
transform 1 0 11500 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_125
timestamp 1667941163
transform 1 0 12604 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_137
timestamp 1667941163
transform 1 0 13708 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_149
timestamp 1667941163
transform 1 0 14812 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_51_161
timestamp 1667941163
transform 1 0 15916 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_166
timestamp 1667941163
transform 1 0 16376 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_169
timestamp 1667941163
transform 1 0 16652 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_51_187
timestamp 1667941163
transform 1 0 18308 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_51_199
timestamp 1667941163
transform 1 0 19412 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_209
timestamp 1667941163
transform 1 0 20332 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_213
timestamp 1667941163
transform 1 0 20700 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_51_217
timestamp 1667941163
transform 1 0 21068 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_223
timestamp 1667941163
transform 1 0 21620 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_225
timestamp 1667941163
transform 1 0 21804 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_237
timestamp 1667941163
transform 1 0 22908 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_249
timestamp 1667941163
transform 1 0 24012 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_261
timestamp 1667941163
transform 1 0 25116 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_51_273
timestamp 1667941163
transform 1 0 26220 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_278
timestamp 1667941163
transform 1 0 26680 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_51_281
timestamp 1667941163
transform 1 0 26956 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_51_292
timestamp 1667941163
transform 1 0 27968 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_298
timestamp 1667941163
transform 1 0 28520 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_3
timestamp 1667941163
transform 1 0 1380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_15
timestamp 1667941163
transform 1 0 2484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_27
timestamp 1667941163
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_29
timestamp 1667941163
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_41
timestamp 1667941163
transform 1 0 4876 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_53
timestamp 1667941163
transform 1 0 5980 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_65
timestamp 1667941163
transform 1 0 7084 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_52_77
timestamp 1667941163
transform 1 0 8188 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_82
timestamp 1667941163
transform 1 0 8648 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_85
timestamp 1667941163
transform 1 0 8924 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_52_108
timestamp 1667941163
transform 1 0 11040 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_120
timestamp 1667941163
transform 1 0 12144 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_132
timestamp 1667941163
transform 1 0 13248 0 1 30464
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_52_141
timestamp 1667941163
transform 1 0 14076 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_153
timestamp 1667941163
transform 1 0 15180 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_159
timestamp 1667941163
transform 1 0 15732 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_165
timestamp 1667941163
transform 1 0 16284 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_177
timestamp 1667941163
transform 1 0 17388 0 1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_52_184
timestamp 1667941163
transform 1 0 18032 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_197
timestamp 1667941163
transform 1 0 19228 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_209
timestamp 1667941163
transform 1 0 20332 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_213
timestamp 1667941163
transform 1 0 20700 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_234
timestamp 1667941163
transform 1 0 22632 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_246
timestamp 1667941163
transform 1 0 23736 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_52_253
timestamp 1667941163
transform 1 0 24380 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_257
timestamp 1667941163
transform 1 0 24748 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_265
timestamp 1667941163
transform 1 0 25484 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_272
timestamp 1667941163
transform 1 0 26128 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_52_297
timestamp 1667941163
transform 1 0 28428 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_53_3
timestamp 1667941163
transform 1 0 1380 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_15
timestamp 1667941163
transform 1 0 2484 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_27
timestamp 1667941163
transform 1 0 3588 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_39
timestamp 1667941163
transform 1 0 4692 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_51
timestamp 1667941163
transform 1 0 5796 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_55
timestamp 1667941163
transform 1 0 6164 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_57
timestamp 1667941163
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_69
timestamp 1667941163
transform 1 0 7452 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_81
timestamp 1667941163
transform 1 0 8556 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_93
timestamp 1667941163
transform 1 0 9660 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_105
timestamp 1667941163
transform 1 0 10764 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_111
timestamp 1667941163
transform 1 0 11316 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_113
timestamp 1667941163
transform 1 0 11500 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_125
timestamp 1667941163
transform 1 0 12604 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_137
timestamp 1667941163
transform 1 0 13708 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_149
timestamp 1667941163
transform 1 0 14812 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_53_157
timestamp 1667941163
transform 1 0 15548 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_53_163
timestamp 1667941163
transform 1 0 16100 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_167
timestamp 1667941163
transform 1 0 16468 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_169
timestamp 1667941163
transform 1 0 16652 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_181
timestamp 1667941163
transform 1 0 17756 0 -1 31552
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_53_190
timestamp 1667941163
transform 1 0 18584 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_202
timestamp 1667941163
transform 1 0 19688 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_214
timestamp 1667941163
transform 1 0 20792 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_222
timestamp 1667941163
transform 1 0 21528 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_53_225
timestamp 1667941163
transform 1 0 21804 0 -1 31552
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_53_236
timestamp 1667941163
transform 1 0 22816 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_53_248
timestamp 1667941163
transform 1 0 23920 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_53_254
timestamp 1667941163
transform 1 0 24472 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_278
timestamp 1667941163
transform 1 0 26680 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_281
timestamp 1667941163
transform 1 0 26956 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_290
timestamp 1667941163
transform 1 0 27784 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_53_297
timestamp 1667941163
transform 1 0 28428 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_54_3
timestamp 1667941163
transform 1 0 1380 0 1 31552
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_54_12
timestamp 1667941163
transform 1 0 2208 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_54_24
timestamp 1667941163
transform 1 0 3312 0 1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_54_29
timestamp 1667941163
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_41
timestamp 1667941163
transform 1 0 4876 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_53
timestamp 1667941163
transform 1 0 5980 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_65
timestamp 1667941163
transform 1 0 7084 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_77
timestamp 1667941163
transform 1 0 8188 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_83
timestamp 1667941163
transform 1 0 8740 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_85
timestamp 1667941163
transform 1 0 8924 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_97
timestamp 1667941163
transform 1 0 10028 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_109
timestamp 1667941163
transform 1 0 11132 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_121
timestamp 1667941163
transform 1 0 12236 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_133
timestamp 1667941163
transform 1 0 13340 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_139
timestamp 1667941163
transform 1 0 13892 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_141
timestamp 1667941163
transform 1 0 14076 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_153
timestamp 1667941163
transform 1 0 15180 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_159
timestamp 1667941163
transform 1 0 15732 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_54_165
timestamp 1667941163
transform 1 0 16284 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_171
timestamp 1667941163
transform 1 0 16836 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_54_188
timestamp 1667941163
transform 1 0 18400 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_54_197
timestamp 1667941163
transform 1 0 19228 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_54_202
timestamp 1667941163
transform 1 0 19688 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_54_210
timestamp 1667941163
transform 1 0 20424 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_218
timestamp 1667941163
transform 1 0 21160 0 1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_54_229
timestamp 1667941163
transform 1 0 22172 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_246
timestamp 1667941163
transform 1 0 23736 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_54_253
timestamp 1667941163
transform 1 0 24380 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_54_261
timestamp 1667941163
transform 1 0 25116 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_54_267
timestamp 1667941163
transform 1 0 25668 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_54_275
timestamp 1667941163
transform 1 0 26404 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_54_297
timestamp 1667941163
transform 1 0 28428 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_55_3
timestamp 1667941163
transform 1 0 1380 0 -1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_55_27
timestamp 1667941163
transform 1 0 3588 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_39
timestamp 1667941163
transform 1 0 4692 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_51
timestamp 1667941163
transform 1 0 5796 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_55
timestamp 1667941163
transform 1 0 6164 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_57
timestamp 1667941163
transform 1 0 6348 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_69
timestamp 1667941163
transform 1 0 7452 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_81
timestamp 1667941163
transform 1 0 8556 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_93
timestamp 1667941163
transform 1 0 9660 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_105
timestamp 1667941163
transform 1 0 10764 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_111
timestamp 1667941163
transform 1 0 11316 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_113
timestamp 1667941163
transform 1 0 11500 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_125
timestamp 1667941163
transform 1 0 12604 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_137
timestamp 1667941163
transform 1 0 13708 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_55_149
timestamp 1667941163
transform 1 0 14812 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_155
timestamp 1667941163
transform 1 0 15364 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_164
timestamp 1667941163
transform 1 0 16192 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_55_169
timestamp 1667941163
transform 1 0 16652 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_55_174
timestamp 1667941163
transform 1 0 17112 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_55_182
timestamp 1667941163
transform 1 0 17848 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_188
timestamp 1667941163
transform 1 0 18400 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_200
timestamp 1667941163
transform 1 0 19504 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_204
timestamp 1667941163
transform 1 0 19872 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_212
timestamp 1667941163
transform 1 0 20608 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_55_225
timestamp 1667941163
transform 1 0 21804 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_244
timestamp 1667941163
transform 1 0 23552 0 -1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_55_257
timestamp 1667941163
transform 1 0 24748 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_269
timestamp 1667941163
transform 1 0 25852 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_55_278
timestamp 1667941163
transform 1 0 26680 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_281
timestamp 1667941163
transform 1 0 26956 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_288
timestamp 1667941163
transform 1 0 27600 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_295
timestamp 1667941163
transform 1 0 28244 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_56_3
timestamp 1667941163
transform 1 0 1380 0 1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_56_9
timestamp 1667941163
transform 1 0 1932 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_21
timestamp 1667941163
transform 1 0 3036 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_27
timestamp 1667941163
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_29
timestamp 1667941163
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_41
timestamp 1667941163
transform 1 0 4876 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_53
timestamp 1667941163
transform 1 0 5980 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_65
timestamp 1667941163
transform 1 0 7084 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_77
timestamp 1667941163
transform 1 0 8188 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_83
timestamp 1667941163
transform 1 0 8740 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_85
timestamp 1667941163
transform 1 0 8924 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_97
timestamp 1667941163
transform 1 0 10028 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_109
timestamp 1667941163
transform 1 0 11132 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_121
timestamp 1667941163
transform 1 0 12236 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_133
timestamp 1667941163
transform 1 0 13340 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_139
timestamp 1667941163
transform 1 0 13892 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_141
timestamp 1667941163
transform 1 0 14076 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_153
timestamp 1667941163
transform 1 0 15180 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_157
timestamp 1667941163
transform 1 0 15548 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_167
timestamp 1667941163
transform 1 0 16468 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_178
timestamp 1667941163
transform 1 0 17480 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_56_189
timestamp 1667941163
transform 1 0 18492 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_195
timestamp 1667941163
transform 1 0 19044 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_56_197
timestamp 1667941163
transform 1 0 19228 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_56_208
timestamp 1667941163
transform 1 0 20240 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_219
timestamp 1667941163
transform 1 0 21252 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_229
timestamp 1667941163
transform 1 0 22172 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_233
timestamp 1667941163
transform 1 0 22540 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_56_250
timestamp 1667941163
transform 1 0 24104 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_253
timestamp 1667941163
transform 1 0 24380 0 1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_56_263
timestamp 1667941163
transform 1 0 25300 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_275
timestamp 1667941163
transform 1 0 26404 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_56_297
timestamp 1667941163
transform 1 0 28428 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_3
timestamp 1667941163
transform 1 0 1380 0 -1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_57_10
timestamp 1667941163
transform 1 0 2024 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_22
timestamp 1667941163
transform 1 0 3128 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_34
timestamp 1667941163
transform 1 0 4232 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_46
timestamp 1667941163
transform 1 0 5336 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_57_54
timestamp 1667941163
transform 1 0 6072 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_57_57
timestamp 1667941163
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_69
timestamp 1667941163
transform 1 0 7452 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_81
timestamp 1667941163
transform 1 0 8556 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_93
timestamp 1667941163
transform 1 0 9660 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_105
timestamp 1667941163
transform 1 0 10764 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_111
timestamp 1667941163
transform 1 0 11316 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_113
timestamp 1667941163
transform 1 0 11500 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_125
timestamp 1667941163
transform 1 0 12604 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_137
timestamp 1667941163
transform 1 0 13708 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_149
timestamp 1667941163
transform 1 0 14812 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_161
timestamp 1667941163
transform 1 0 15916 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_167
timestamp 1667941163
transform 1 0 16468 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_169
timestamp 1667941163
transform 1 0 16652 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_57_181
timestamp 1667941163
transform 1 0 17756 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_190
timestamp 1667941163
transform 1 0 18584 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_57_199
timestamp 1667941163
transform 1 0 19412 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_57_214
timestamp 1667941163
transform 1 0 20792 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_57_222
timestamp 1667941163
transform 1 0 21528 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_225
timestamp 1667941163
transform 1 0 21804 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_57_230
timestamp 1667941163
transform 1 0 22264 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_57_238
timestamp 1667941163
transform 1 0 23000 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_243
timestamp 1667941163
transform 1 0 23460 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_57_250
timestamp 1667941163
transform 1 0 24104 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_57_272
timestamp 1667941163
transform 1 0 26128 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_57_281
timestamp 1667941163
transform 1 0 26956 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_286
timestamp 1667941163
transform 1 0 27416 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_290
timestamp 1667941163
transform 1 0 27784 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_294
timestamp 1667941163
transform 1 0 28152 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_298
timestamp 1667941163
transform 1 0 28520 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_58_3
timestamp 1667941163
transform 1 0 1380 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_9
timestamp 1667941163
transform 1 0 1932 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_13
timestamp 1667941163
transform 1 0 2300 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_58_25
timestamp 1667941163
transform 1 0 3404 0 1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_58_29
timestamp 1667941163
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_41
timestamp 1667941163
transform 1 0 4876 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_53
timestamp 1667941163
transform 1 0 5980 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_65
timestamp 1667941163
transform 1 0 7084 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_77
timestamp 1667941163
transform 1 0 8188 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_83
timestamp 1667941163
transform 1 0 8740 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_85
timestamp 1667941163
transform 1 0 8924 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_97
timestamp 1667941163
transform 1 0 10028 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_109
timestamp 1667941163
transform 1 0 11132 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_121
timestamp 1667941163
transform 1 0 12236 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_133
timestamp 1667941163
transform 1 0 13340 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_139
timestamp 1667941163
transform 1 0 13892 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_141
timestamp 1667941163
transform 1 0 14076 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_153
timestamp 1667941163
transform 1 0 15180 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_165
timestamp 1667941163
transform 1 0 16284 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_177
timestamp 1667941163
transform 1 0 17388 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_189
timestamp 1667941163
transform 1 0 18492 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_195
timestamp 1667941163
transform 1 0 19044 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_197
timestamp 1667941163
transform 1 0 19228 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_209
timestamp 1667941163
transform 1 0 20332 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_58_233
timestamp 1667941163
transform 1 0 22540 0 1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_58_240
timestamp 1667941163
transform 1 0 23184 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_58_253
timestamp 1667941163
transform 1 0 24380 0 1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_58_259
timestamp 1667941163
transform 1 0 24932 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_58_271
timestamp 1667941163
transform 1 0 26036 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_294
timestamp 1667941163
transform 1 0 28152 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_298
timestamp 1667941163
transform 1 0 28520 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_59_3
timestamp 1667941163
transform 1 0 1380 0 -1 34816
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_59_27
timestamp 1667941163
transform 1 0 3588 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_39
timestamp 1667941163
transform 1 0 4692 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_51
timestamp 1667941163
transform 1 0 5796 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_55
timestamp 1667941163
transform 1 0 6164 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_57
timestamp 1667941163
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_69
timestamp 1667941163
transform 1 0 7452 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_81
timestamp 1667941163
transform 1 0 8556 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_93
timestamp 1667941163
transform 1 0 9660 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_105
timestamp 1667941163
transform 1 0 10764 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_111
timestamp 1667941163
transform 1 0 11316 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_113
timestamp 1667941163
transform 1 0 11500 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_125
timestamp 1667941163
transform 1 0 12604 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_137
timestamp 1667941163
transform 1 0 13708 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_149
timestamp 1667941163
transform 1 0 14812 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_161
timestamp 1667941163
transform 1 0 15916 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_167
timestamp 1667941163
transform 1 0 16468 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_169
timestamp 1667941163
transform 1 0 16652 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_181
timestamp 1667941163
transform 1 0 17756 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_193
timestamp 1667941163
transform 1 0 18860 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_197
timestamp 1667941163
transform 1 0 19228 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_201
timestamp 1667941163
transform 1 0 19596 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_213
timestamp 1667941163
transform 1 0 20700 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_59_221
timestamp 1667941163
transform 1 0 21436 0 -1 34816
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_59_225
timestamp 1667941163
transform 1 0 21804 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_237
timestamp 1667941163
transform 1 0 22908 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_249
timestamp 1667941163
transform 1 0 24012 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_59_261
timestamp 1667941163
transform 1 0 25116 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_59_278
timestamp 1667941163
transform 1 0 26680 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_281
timestamp 1667941163
transform 1 0 26956 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_59_291
timestamp 1667941163
transform 1 0 27876 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_60_3
timestamp 1667941163
transform 1 0 1380 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_60_16
timestamp 1667941163
transform 1 0 2576 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_23
timestamp 1667941163
transform 1 0 3220 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_27
timestamp 1667941163
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_29
timestamp 1667941163
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_41
timestamp 1667941163
transform 1 0 4876 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_53
timestamp 1667941163
transform 1 0 5980 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_65
timestamp 1667941163
transform 1 0 7084 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_77
timestamp 1667941163
transform 1 0 8188 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_83
timestamp 1667941163
transform 1 0 8740 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_85
timestamp 1667941163
transform 1 0 8924 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_97
timestamp 1667941163
transform 1 0 10028 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_109
timestamp 1667941163
transform 1 0 11132 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_121
timestamp 1667941163
transform 1 0 12236 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_133
timestamp 1667941163
transform 1 0 13340 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_139
timestamp 1667941163
transform 1 0 13892 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_141
timestamp 1667941163
transform 1 0 14076 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_153
timestamp 1667941163
transform 1 0 15180 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_165
timestamp 1667941163
transform 1 0 16284 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_60_187
timestamp 1667941163
transform 1 0 18308 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_60_195
timestamp 1667941163
transform 1 0 19044 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_60_197
timestamp 1667941163
transform 1 0 19228 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_60_215
timestamp 1667941163
transform 1 0 20884 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_235
timestamp 1667941163
transform 1 0 22724 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_60_244
timestamp 1667941163
transform 1 0 23552 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_60_253
timestamp 1667941163
transform 1 0 24380 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_60_258
timestamp 1667941163
transform 1 0 24840 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_265
timestamp 1667941163
transform 1 0 25484 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_272
timestamp 1667941163
transform 1 0 26128 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_60_297
timestamp 1667941163
transform 1 0 28428 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_61_3
timestamp 1667941163
transform 1 0 1380 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_61_27
timestamp 1667941163
transform 1 0 3588 0 -1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_61_43
timestamp 1667941163
transform 1 0 5060 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_61_55
timestamp 1667941163
transform 1 0 6164 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_57
timestamp 1667941163
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_69
timestamp 1667941163
transform 1 0 7452 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_81
timestamp 1667941163
transform 1 0 8556 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_93
timestamp 1667941163
transform 1 0 9660 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_105
timestamp 1667941163
transform 1 0 10764 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_111
timestamp 1667941163
transform 1 0 11316 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_113
timestamp 1667941163
transform 1 0 11500 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_125
timestamp 1667941163
transform 1 0 12604 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_137
timestamp 1667941163
transform 1 0 13708 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_149
timestamp 1667941163
transform 1 0 14812 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_61_166
timestamp 1667941163
transform 1 0 16376 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_169
timestamp 1667941163
transform 1 0 16652 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_61_187
timestamp 1667941163
transform 1 0 18308 0 -1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_61_207
timestamp 1667941163
transform 1 0 20148 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_219
timestamp 1667941163
transform 1 0 21252 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_223
timestamp 1667941163
transform 1 0 21620 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_61_225
timestamp 1667941163
transform 1 0 21804 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_61_247
timestamp 1667941163
transform 1 0 23828 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_268
timestamp 1667941163
transform 1 0 25760 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_275
timestamp 1667941163
transform 1 0 26404 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_279
timestamp 1667941163
transform 1 0 26772 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_61_281
timestamp 1667941163
transform 1 0 26956 0 -1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_61_286
timestamp 1667941163
transform 1 0 27416 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_61_298
timestamp 1667941163
transform 1 0 28520 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_3
timestamp 1667941163
transform 1 0 1380 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_10
timestamp 1667941163
transform 1 0 2024 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_62_26
timestamp 1667941163
transform 1 0 3496 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_62_29
timestamp 1667941163
transform 1 0 3772 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_43
timestamp 1667941163
transform 1 0 5060 0 1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_62_56
timestamp 1667941163
transform 1 0 6256 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_68
timestamp 1667941163
transform 1 0 7360 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_62_80
timestamp 1667941163
transform 1 0 8464 0 1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_62_85
timestamp 1667941163
transform 1 0 8924 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_97
timestamp 1667941163
transform 1 0 10028 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_109
timestamp 1667941163
transform 1 0 11132 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_121
timestamp 1667941163
transform 1 0 12236 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_133
timestamp 1667941163
transform 1 0 13340 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_139
timestamp 1667941163
transform 1 0 13892 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_141
timestamp 1667941163
transform 1 0 14076 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_153
timestamp 1667941163
transform 1 0 15180 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_62_168
timestamp 1667941163
transform 1 0 16560 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_175
timestamp 1667941163
transform 1 0 17204 0 1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_62_182
timestamp 1667941163
transform 1 0 17848 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_62_194
timestamp 1667941163
transform 1 0 18952 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_62_197
timestamp 1667941163
transform 1 0 19228 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_62_205
timestamp 1667941163
transform 1 0 19964 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_62_222
timestamp 1667941163
transform 1 0 21528 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_62_230
timestamp 1667941163
transform 1 0 22264 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_235
timestamp 1667941163
transform 1 0 22724 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_248
timestamp 1667941163
transform 1 0 23920 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_62_253
timestamp 1667941163
transform 1 0 24380 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_62_264
timestamp 1667941163
transform 1 0 25392 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_289
timestamp 1667941163
transform 1 0 27692 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_62_296
timestamp 1667941163
transform 1 0 28336 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_63_3
timestamp 1667941163
transform 1 0 1380 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_19
timestamp 1667941163
transform 1 0 2852 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_35
timestamp 1667941163
transform 1 0 4324 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_51
timestamp 1667941163
transform 1 0 5796 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_55
timestamp 1667941163
transform 1 0 6164 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_57
timestamp 1667941163
transform 1 0 6348 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_69
timestamp 1667941163
transform 1 0 7452 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_81
timestamp 1667941163
transform 1 0 8556 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_93
timestamp 1667941163
transform 1 0 9660 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_105
timestamp 1667941163
transform 1 0 10764 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_111
timestamp 1667941163
transform 1 0 11316 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_113
timestamp 1667941163
transform 1 0 11500 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_125
timestamp 1667941163
transform 1 0 12604 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_137
timestamp 1667941163
transform 1 0 13708 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_149
timestamp 1667941163
transform 1 0 14812 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_161
timestamp 1667941163
transform 1 0 15916 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_167
timestamp 1667941163
transform 1 0 16468 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_63_169
timestamp 1667941163
transform 1 0 16652 0 -1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_63_176
timestamp 1667941163
transform 1 0 17296 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_191
timestamp 1667941163
transform 1 0 18676 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_203
timestamp 1667941163
transform 1 0 19780 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_215
timestamp 1667941163
transform 1 0 20884 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_63_222
timestamp 1667941163
transform 1 0 21528 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_63_225
timestamp 1667941163
transform 1 0 21804 0 -1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_63_234
timestamp 1667941163
transform 1 0 22632 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_246
timestamp 1667941163
transform 1 0 23736 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_258
timestamp 1667941163
transform 1 0 24840 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_63_278
timestamp 1667941163
transform 1 0 26680 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_281
timestamp 1667941163
transform 1 0 26956 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_63_286
timestamp 1667941163
transform 1 0 27416 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_63_293
timestamp 1667941163
transform 1 0 28060 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_64_3
timestamp 1667941163
transform 1 0 1380 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_10
timestamp 1667941163
transform 1 0 2024 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_64_26
timestamp 1667941163
transform 1 0 3496 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_29
timestamp 1667941163
transform 1 0 3772 0 1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_64_43
timestamp 1667941163
transform 1 0 5060 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_55
timestamp 1667941163
transform 1 0 6164 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_67
timestamp 1667941163
transform 1 0 7268 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_79
timestamp 1667941163
transform 1 0 8372 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_83
timestamp 1667941163
transform 1 0 8740 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_85
timestamp 1667941163
transform 1 0 8924 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_97
timestamp 1667941163
transform 1 0 10028 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_109
timestamp 1667941163
transform 1 0 11132 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_121
timestamp 1667941163
transform 1 0 12236 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_133
timestamp 1667941163
transform 1 0 13340 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_139
timestamp 1667941163
transform 1 0 13892 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_141
timestamp 1667941163
transform 1 0 14076 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_153
timestamp 1667941163
transform 1 0 15180 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_165
timestamp 1667941163
transform 1 0 16284 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_178
timestamp 1667941163
transform 1 0 17480 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_64_189
timestamp 1667941163
transform 1 0 18492 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_195
timestamp 1667941163
transform 1 0 19044 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_197
timestamp 1667941163
transform 1 0 19228 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_206
timestamp 1667941163
transform 1 0 20056 0 1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_64_216
timestamp 1667941163
transform 1 0 20976 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_228
timestamp 1667941163
transform 1 0 22080 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_240
timestamp 1667941163
transform 1 0 23184 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_253
timestamp 1667941163
transform 1 0 24380 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_265
timestamp 1667941163
transform 1 0 25484 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_64_273
timestamp 1667941163
transform 1 0 26220 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_64_297
timestamp 1667941163
transform 1 0 28428 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_65_3
timestamp 1667941163
transform 1 0 1380 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_65_27
timestamp 1667941163
transform 1 0 3588 0 -1 38080
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_65_34
timestamp 1667941163
transform 1 0 4232 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_65_46
timestamp 1667941163
transform 1 0 5336 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_65_54
timestamp 1667941163
transform 1 0 6072 0 -1 38080
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_65_57
timestamp 1667941163
transform 1 0 6348 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_69
timestamp 1667941163
transform 1 0 7452 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_81
timestamp 1667941163
transform 1 0 8556 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_93
timestamp 1667941163
transform 1 0 9660 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_105
timestamp 1667941163
transform 1 0 10764 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_111
timestamp 1667941163
transform 1 0 11316 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_113
timestamp 1667941163
transform 1 0 11500 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_125
timestamp 1667941163
transform 1 0 12604 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_137
timestamp 1667941163
transform 1 0 13708 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_149
timestamp 1667941163
transform 1 0 14812 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_161
timestamp 1667941163
transform 1 0 15916 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_167
timestamp 1667941163
transform 1 0 16468 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_169
timestamp 1667941163
transform 1 0 16652 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_181
timestamp 1667941163
transform 1 0 17756 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_187
timestamp 1667941163
transform 1 0 18308 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_65_191
timestamp 1667941163
transform 1 0 18676 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_65_198
timestamp 1667941163
transform 1 0 19320 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_65_213
timestamp 1667941163
transform 1 0 20700 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_65_222
timestamp 1667941163
transform 1 0 21528 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_65_225
timestamp 1667941163
transform 1 0 21804 0 -1 38080
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_65_230
timestamp 1667941163
transform 1 0 22264 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_242
timestamp 1667941163
transform 1 0 23368 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_254
timestamp 1667941163
transform 1 0 24472 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_266
timestamp 1667941163
transform 1 0 25576 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_65_278
timestamp 1667941163
transform 1 0 26680 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_65_281
timestamp 1667941163
transform 1 0 26956 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_65_295
timestamp 1667941163
transform 1 0 28244 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_66_3
timestamp 1667941163
transform 1 0 1380 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_66_26
timestamp 1667941163
transform 1 0 3496 0 1 38080
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_66_29
timestamp 1667941163
transform 1 0 3772 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_41
timestamp 1667941163
transform 1 0 4876 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_53
timestamp 1667941163
transform 1 0 5980 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_65
timestamp 1667941163
transform 1 0 7084 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_77
timestamp 1667941163
transform 1 0 8188 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_83
timestamp 1667941163
transform 1 0 8740 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_85
timestamp 1667941163
transform 1 0 8924 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_97
timestamp 1667941163
transform 1 0 10028 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_109
timestamp 1667941163
transform 1 0 11132 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_121
timestamp 1667941163
transform 1 0 12236 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_133
timestamp 1667941163
transform 1 0 13340 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_139
timestamp 1667941163
transform 1 0 13892 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_141
timestamp 1667941163
transform 1 0 14076 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_153
timestamp 1667941163
transform 1 0 15180 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_165
timestamp 1667941163
transform 1 0 16284 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_177
timestamp 1667941163
transform 1 0 17388 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_66_194
timestamp 1667941163
transform 1 0 18952 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_66_197
timestamp 1667941163
transform 1 0 19228 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_66_212
timestamp 1667941163
transform 1 0 20608 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_221
timestamp 1667941163
transform 1 0 21436 0 1 38080
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_66_230
timestamp 1667941163
transform 1 0 22264 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_66_242
timestamp 1667941163
transform 1 0 23368 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_66_250
timestamp 1667941163
transform 1 0 24104 0 1 38080
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_66_253
timestamp 1667941163
transform 1 0 24380 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_66_265
timestamp 1667941163
transform 1 0 25484 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_272
timestamp 1667941163
transform 1 0 26128 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_66_297
timestamp 1667941163
transform 1 0 28428 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_67_3
timestamp 1667941163
transform 1 0 1380 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_67_8
timestamp 1667941163
transform 1 0 1840 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_67_16
timestamp 1667941163
transform 1 0 2576 0 -1 39168
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_67_39
timestamp 1667941163
transform 1 0 4692 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_51
timestamp 1667941163
transform 1 0 5796 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_55
timestamp 1667941163
transform 1 0 6164 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_57
timestamp 1667941163
transform 1 0 6348 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_69
timestamp 1667941163
transform 1 0 7452 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_81
timestamp 1667941163
transform 1 0 8556 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_93
timestamp 1667941163
transform 1 0 9660 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_105
timestamp 1667941163
transform 1 0 10764 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_111
timestamp 1667941163
transform 1 0 11316 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_113
timestamp 1667941163
transform 1 0 11500 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_125
timestamp 1667941163
transform 1 0 12604 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_137
timestamp 1667941163
transform 1 0 13708 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_149
timestamp 1667941163
transform 1 0 14812 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_161
timestamp 1667941163
transform 1 0 15916 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_167
timestamp 1667941163
transform 1 0 16468 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_169
timestamp 1667941163
transform 1 0 16652 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_181
timestamp 1667941163
transform 1 0 17756 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_67_193
timestamp 1667941163
transform 1 0 18860 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_67_197
timestamp 1667941163
transform 1 0 19228 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_207
timestamp 1667941163
transform 1 0 20148 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_214
timestamp 1667941163
transform 1 0 20792 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_67_221
timestamp 1667941163
transform 1 0 21436 0 -1 39168
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_67_225
timestamp 1667941163
transform 1 0 21804 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_237
timestamp 1667941163
transform 1 0 22908 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_249
timestamp 1667941163
transform 1 0 24012 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_261
timestamp 1667941163
transform 1 0 25116 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_67_273
timestamp 1667941163
transform 1 0 26220 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_67_278
timestamp 1667941163
transform 1 0 26680 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_67_281
timestamp 1667941163
transform 1 0 26956 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_67_286
timestamp 1667941163
transform 1 0 27416 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_67_293
timestamp 1667941163
transform 1 0 28060 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_68_3
timestamp 1667941163
transform 1 0 1380 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_10
timestamp 1667941163
transform 1 0 2024 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_17
timestamp 1667941163
transform 1 0 2668 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_24
timestamp 1667941163
transform 1 0 3312 0 1 39168
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_68_29
timestamp 1667941163
transform 1 0 3772 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_41
timestamp 1667941163
transform 1 0 4876 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_53
timestamp 1667941163
transform 1 0 5980 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_65
timestamp 1667941163
transform 1 0 7084 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_77
timestamp 1667941163
transform 1 0 8188 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_83
timestamp 1667941163
transform 1 0 8740 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_85
timestamp 1667941163
transform 1 0 8924 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_97
timestamp 1667941163
transform 1 0 10028 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_109
timestamp 1667941163
transform 1 0 11132 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_121
timestamp 1667941163
transform 1 0 12236 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_133
timestamp 1667941163
transform 1 0 13340 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_139
timestamp 1667941163
transform 1 0 13892 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_141
timestamp 1667941163
transform 1 0 14076 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_153
timestamp 1667941163
transform 1 0 15180 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_165
timestamp 1667941163
transform 1 0 16284 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_177
timestamp 1667941163
transform 1 0 17388 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_189
timestamp 1667941163
transform 1 0 18492 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_195
timestamp 1667941163
transform 1 0 19044 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_197
timestamp 1667941163
transform 1 0 19228 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_209
timestamp 1667941163
transform 1 0 20332 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_221
timestamp 1667941163
transform 1 0 21436 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_233
timestamp 1667941163
transform 1 0 22540 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_245
timestamp 1667941163
transform 1 0 23644 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_251
timestamp 1667941163
transform 1 0 24196 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_253
timestamp 1667941163
transform 1 0 24380 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_68_265
timestamp 1667941163
transform 1 0 25484 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_68_273
timestamp 1667941163
transform 1 0 26220 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_68_297
timestamp 1667941163
transform 1 0 28428 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_69_3
timestamp 1667941163
transform 1 0 1380 0 -1 40256
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_69_10
timestamp 1667941163
transform 1 0 2024 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_22
timestamp 1667941163
transform 1 0 3128 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_34
timestamp 1667941163
transform 1 0 4232 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_69_46
timestamp 1667941163
transform 1 0 5336 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_69_54
timestamp 1667941163
transform 1 0 6072 0 -1 40256
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_69_57
timestamp 1667941163
transform 1 0 6348 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_69
timestamp 1667941163
transform 1 0 7452 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_81
timestamp 1667941163
transform 1 0 8556 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_93
timestamp 1667941163
transform 1 0 9660 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_105
timestamp 1667941163
transform 1 0 10764 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_111
timestamp 1667941163
transform 1 0 11316 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_113
timestamp 1667941163
transform 1 0 11500 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_125
timestamp 1667941163
transform 1 0 12604 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_137
timestamp 1667941163
transform 1 0 13708 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_149
timestamp 1667941163
transform 1 0 14812 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_161
timestamp 1667941163
transform 1 0 15916 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_167
timestamp 1667941163
transform 1 0 16468 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_169
timestamp 1667941163
transform 1 0 16652 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_181
timestamp 1667941163
transform 1 0 17756 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_193
timestamp 1667941163
transform 1 0 18860 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_205
timestamp 1667941163
transform 1 0 19964 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_217
timestamp 1667941163
transform 1 0 21068 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_223
timestamp 1667941163
transform 1 0 21620 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_225
timestamp 1667941163
transform 1 0 21804 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_237
timestamp 1667941163
transform 1 0 22908 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_249
timestamp 1667941163
transform 1 0 24012 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_261
timestamp 1667941163
transform 1 0 25116 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_273
timestamp 1667941163
transform 1 0 26220 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_279
timestamp 1667941163
transform 1 0 26772 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_69_281
timestamp 1667941163
transform 1 0 26956 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_69_287
timestamp 1667941163
transform 1 0 27508 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_294
timestamp 1667941163
transform 1 0 28152 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_298
timestamp 1667941163
transform 1 0 28520 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_70_3
timestamp 1667941163
transform 1 0 1380 0 1 40256
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_70_14
timestamp 1667941163
transform 1 0 2392 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_70_26
timestamp 1667941163
transform 1 0 3496 0 1 40256
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_70_29
timestamp 1667941163
transform 1 0 3772 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_41
timestamp 1667941163
transform 1 0 4876 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_53
timestamp 1667941163
transform 1 0 5980 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_65
timestamp 1667941163
transform 1 0 7084 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_77
timestamp 1667941163
transform 1 0 8188 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_83
timestamp 1667941163
transform 1 0 8740 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_85
timestamp 1667941163
transform 1 0 8924 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_97
timestamp 1667941163
transform 1 0 10028 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_109
timestamp 1667941163
transform 1 0 11132 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_121
timestamp 1667941163
transform 1 0 12236 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_133
timestamp 1667941163
transform 1 0 13340 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_139
timestamp 1667941163
transform 1 0 13892 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_141
timestamp 1667941163
transform 1 0 14076 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_153
timestamp 1667941163
transform 1 0 15180 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_165
timestamp 1667941163
transform 1 0 16284 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_177
timestamp 1667941163
transform 1 0 17388 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_189
timestamp 1667941163
transform 1 0 18492 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_195
timestamp 1667941163
transform 1 0 19044 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_197
timestamp 1667941163
transform 1 0 19228 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_209
timestamp 1667941163
transform 1 0 20332 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_221
timestamp 1667941163
transform 1 0 21436 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_233
timestamp 1667941163
transform 1 0 22540 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_245
timestamp 1667941163
transform 1 0 23644 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_251
timestamp 1667941163
transform 1 0 24196 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_253
timestamp 1667941163
transform 1 0 24380 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_70_265
timestamp 1667941163
transform 1 0 25484 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_70_273
timestamp 1667941163
transform 1 0 26220 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_70_297
timestamp 1667941163
transform 1 0 28428 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_71_3
timestamp 1667941163
transform 1 0 1380 0 -1 41344
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_71_27
timestamp 1667941163
transform 1 0 3588 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_39
timestamp 1667941163
transform 1 0 4692 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_71_51
timestamp 1667941163
transform 1 0 5796 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_55
timestamp 1667941163
transform 1 0 6164 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_57
timestamp 1667941163
transform 1 0 6348 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_69
timestamp 1667941163
transform 1 0 7452 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_81
timestamp 1667941163
transform 1 0 8556 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_93
timestamp 1667941163
transform 1 0 9660 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_105
timestamp 1667941163
transform 1 0 10764 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_111
timestamp 1667941163
transform 1 0 11316 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_113
timestamp 1667941163
transform 1 0 11500 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_125
timestamp 1667941163
transform 1 0 12604 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_137
timestamp 1667941163
transform 1 0 13708 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_149
timestamp 1667941163
transform 1 0 14812 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_161
timestamp 1667941163
transform 1 0 15916 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_167
timestamp 1667941163
transform 1 0 16468 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_169
timestamp 1667941163
transform 1 0 16652 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_181
timestamp 1667941163
transform 1 0 17756 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_193
timestamp 1667941163
transform 1 0 18860 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_205
timestamp 1667941163
transform 1 0 19964 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_217
timestamp 1667941163
transform 1 0 21068 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_223
timestamp 1667941163
transform 1 0 21620 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_225
timestamp 1667941163
transform 1 0 21804 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_237
timestamp 1667941163
transform 1 0 22908 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_249
timestamp 1667941163
transform 1 0 24012 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_261
timestamp 1667941163
transform 1 0 25116 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_273
timestamp 1667941163
transform 1 0 26220 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_279
timestamp 1667941163
transform 1 0 26772 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_71_281
timestamp 1667941163
transform 1 0 26956 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_71_286
timestamp 1667941163
transform 1 0 27416 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_290
timestamp 1667941163
transform 1 0 27784 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_71_294
timestamp 1667941163
transform 1 0 28152 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_298
timestamp 1667941163
transform 1 0 28520 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_72_3
timestamp 1667941163
transform 1 0 1380 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_72_26
timestamp 1667941163
transform 1 0 3496 0 1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_72_29
timestamp 1667941163
transform 1 0 3772 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_41
timestamp 1667941163
transform 1 0 4876 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_53
timestamp 1667941163
transform 1 0 5980 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_65
timestamp 1667941163
transform 1 0 7084 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_77
timestamp 1667941163
transform 1 0 8188 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_83
timestamp 1667941163
transform 1 0 8740 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_85
timestamp 1667941163
transform 1 0 8924 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_97
timestamp 1667941163
transform 1 0 10028 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_109
timestamp 1667941163
transform 1 0 11132 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_121
timestamp 1667941163
transform 1 0 12236 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_133
timestamp 1667941163
transform 1 0 13340 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_139
timestamp 1667941163
transform 1 0 13892 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_141
timestamp 1667941163
transform 1 0 14076 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_153
timestamp 1667941163
transform 1 0 15180 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_165
timestamp 1667941163
transform 1 0 16284 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_177
timestamp 1667941163
transform 1 0 17388 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_189
timestamp 1667941163
transform 1 0 18492 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_195
timestamp 1667941163
transform 1 0 19044 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_197
timestamp 1667941163
transform 1 0 19228 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_209
timestamp 1667941163
transform 1 0 20332 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_221
timestamp 1667941163
transform 1 0 21436 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_233
timestamp 1667941163
transform 1 0 22540 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_245
timestamp 1667941163
transform 1 0 23644 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_251
timestamp 1667941163
transform 1 0 24196 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_253
timestamp 1667941163
transform 1 0 24380 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_72_265
timestamp 1667941163
transform 1 0 25484 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_72_273
timestamp 1667941163
transform 1 0 26220 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_72_297
timestamp 1667941163
transform 1 0 28428 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_73_3
timestamp 1667941163
transform 1 0 1380 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_10
timestamp 1667941163
transform 1 0 2024 0 -1 42432
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_73_17
timestamp 1667941163
transform 1 0 2668 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_29
timestamp 1667941163
transform 1 0 3772 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_41
timestamp 1667941163
transform 1 0 4876 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_73_53
timestamp 1667941163
transform 1 0 5980 0 -1 42432
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_73_57
timestamp 1667941163
transform 1 0 6348 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_69
timestamp 1667941163
transform 1 0 7452 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_81
timestamp 1667941163
transform 1 0 8556 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_93
timestamp 1667941163
transform 1 0 9660 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_105
timestamp 1667941163
transform 1 0 10764 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_111
timestamp 1667941163
transform 1 0 11316 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_113
timestamp 1667941163
transform 1 0 11500 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_125
timestamp 1667941163
transform 1 0 12604 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_137
timestamp 1667941163
transform 1 0 13708 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_149
timestamp 1667941163
transform 1 0 14812 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_161
timestamp 1667941163
transform 1 0 15916 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_167
timestamp 1667941163
transform 1 0 16468 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_169
timestamp 1667941163
transform 1 0 16652 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_181
timestamp 1667941163
transform 1 0 17756 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_193
timestamp 1667941163
transform 1 0 18860 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_205
timestamp 1667941163
transform 1 0 19964 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_217
timestamp 1667941163
transform 1 0 21068 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_223
timestamp 1667941163
transform 1 0 21620 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_225
timestamp 1667941163
transform 1 0 21804 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_237
timestamp 1667941163
transform 1 0 22908 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_73_249
timestamp 1667941163
transform 1 0 24012 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_73_278
timestamp 1667941163
transform 1 0 26680 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_73_281
timestamp 1667941163
transform 1 0 26956 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_73_292
timestamp 1667941163
transform 1 0 27968 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_298
timestamp 1667941163
transform 1 0 28520 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_74_3
timestamp 1667941163
transform 1 0 1380 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_10
timestamp 1667941163
transform 1 0 2024 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_74_17
timestamp 1667941163
transform 1 0 2668 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_74_25
timestamp 1667941163
transform 1 0 3404 0 1 42432
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_74_29
timestamp 1667941163
transform 1 0 3772 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_41
timestamp 1667941163
transform 1 0 4876 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_53
timestamp 1667941163
transform 1 0 5980 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_65
timestamp 1667941163
transform 1 0 7084 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_77
timestamp 1667941163
transform 1 0 8188 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_83
timestamp 1667941163
transform 1 0 8740 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_85
timestamp 1667941163
transform 1 0 8924 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_97
timestamp 1667941163
transform 1 0 10028 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_109
timestamp 1667941163
transform 1 0 11132 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_121
timestamp 1667941163
transform 1 0 12236 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_133
timestamp 1667941163
transform 1 0 13340 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_139
timestamp 1667941163
transform 1 0 13892 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_141
timestamp 1667941163
transform 1 0 14076 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_153
timestamp 1667941163
transform 1 0 15180 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_165
timestamp 1667941163
transform 1 0 16284 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_177
timestamp 1667941163
transform 1 0 17388 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_189
timestamp 1667941163
transform 1 0 18492 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_195
timestamp 1667941163
transform 1 0 19044 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_197
timestamp 1667941163
transform 1 0 19228 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_209
timestamp 1667941163
transform 1 0 20332 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_221
timestamp 1667941163
transform 1 0 21436 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_233
timestamp 1667941163
transform 1 0 22540 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_245
timestamp 1667941163
transform 1 0 23644 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_251
timestamp 1667941163
transform 1 0 24196 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_253
timestamp 1667941163
transform 1 0 24380 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_74_265
timestamp 1667941163
transform 1 0 25484 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_74_273
timestamp 1667941163
transform 1 0 26220 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_74_297
timestamp 1667941163
transform 1 0 28428 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_75_3
timestamp 1667941163
transform 1 0 1380 0 -1 43520
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_75_30
timestamp 1667941163
transform 1 0 3864 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_42
timestamp 1667941163
transform 1 0 4968 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_75_54
timestamp 1667941163
transform 1 0 6072 0 -1 43520
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_75_57
timestamp 1667941163
transform 1 0 6348 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_69
timestamp 1667941163
transform 1 0 7452 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_81
timestamp 1667941163
transform 1 0 8556 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_93
timestamp 1667941163
transform 1 0 9660 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_105
timestamp 1667941163
transform 1 0 10764 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_111
timestamp 1667941163
transform 1 0 11316 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_113
timestamp 1667941163
transform 1 0 11500 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_125
timestamp 1667941163
transform 1 0 12604 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_137
timestamp 1667941163
transform 1 0 13708 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_149
timestamp 1667941163
transform 1 0 14812 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_161
timestamp 1667941163
transform 1 0 15916 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_167
timestamp 1667941163
transform 1 0 16468 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_169
timestamp 1667941163
transform 1 0 16652 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_181
timestamp 1667941163
transform 1 0 17756 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_193
timestamp 1667941163
transform 1 0 18860 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_205
timestamp 1667941163
transform 1 0 19964 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_217
timestamp 1667941163
transform 1 0 21068 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_223
timestamp 1667941163
transform 1 0 21620 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_225
timestamp 1667941163
transform 1 0 21804 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_237
timestamp 1667941163
transform 1 0 22908 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_249
timestamp 1667941163
transform 1 0 24012 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_75_261
timestamp 1667941163
transform 1 0 25116 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_75_272
timestamp 1667941163
transform 1 0 26128 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_75_281
timestamp 1667941163
transform 1 0 26956 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_75_287
timestamp 1667941163
transform 1 0 27508 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_294
timestamp 1667941163
transform 1 0 28152 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_298
timestamp 1667941163
transform 1 0 28520 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_76_3
timestamp 1667941163
transform 1 0 1380 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_76_26
timestamp 1667941163
transform 1 0 3496 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_76_29
timestamp 1667941163
transform 1 0 3772 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_76_34
timestamp 1667941163
transform 1 0 4232 0 1 43520
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_76_41
timestamp 1667941163
transform 1 0 4876 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_53
timestamp 1667941163
transform 1 0 5980 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_65
timestamp 1667941163
transform 1 0 7084 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_77
timestamp 1667941163
transform 1 0 8188 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_83
timestamp 1667941163
transform 1 0 8740 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_85
timestamp 1667941163
transform 1 0 8924 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_97
timestamp 1667941163
transform 1 0 10028 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_109
timestamp 1667941163
transform 1 0 11132 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_121
timestamp 1667941163
transform 1 0 12236 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_133
timestamp 1667941163
transform 1 0 13340 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_139
timestamp 1667941163
transform 1 0 13892 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_141
timestamp 1667941163
transform 1 0 14076 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_153
timestamp 1667941163
transform 1 0 15180 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_165
timestamp 1667941163
transform 1 0 16284 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_177
timestamp 1667941163
transform 1 0 17388 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_189
timestamp 1667941163
transform 1 0 18492 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_195
timestamp 1667941163
transform 1 0 19044 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_197
timestamp 1667941163
transform 1 0 19228 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_209
timestamp 1667941163
transform 1 0 20332 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_221
timestamp 1667941163
transform 1 0 21436 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_233
timestamp 1667941163
transform 1 0 22540 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_245
timestamp 1667941163
transform 1 0 23644 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_251
timestamp 1667941163
transform 1 0 24196 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_253
timestamp 1667941163
transform 1 0 24380 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_76_265
timestamp 1667941163
transform 1 0 25484 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_290
timestamp 1667941163
transform 1 0 27784 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_76_297
timestamp 1667941163
transform 1 0 28428 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_77_3
timestamp 1667941163
transform 1 0 1380 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_77_14
timestamp 1667941163
transform 1 0 2392 0 -1 44608
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_77_43
timestamp 1667941163
transform 1 0 5060 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_77_55
timestamp 1667941163
transform 1 0 6164 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_57
timestamp 1667941163
transform 1 0 6348 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_69
timestamp 1667941163
transform 1 0 7452 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_81
timestamp 1667941163
transform 1 0 8556 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_93
timestamp 1667941163
transform 1 0 9660 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_105
timestamp 1667941163
transform 1 0 10764 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_111
timestamp 1667941163
transform 1 0 11316 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_113
timestamp 1667941163
transform 1 0 11500 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_125
timestamp 1667941163
transform 1 0 12604 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_137
timestamp 1667941163
transform 1 0 13708 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_149
timestamp 1667941163
transform 1 0 14812 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_161
timestamp 1667941163
transform 1 0 15916 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_167
timestamp 1667941163
transform 1 0 16468 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_169
timestamp 1667941163
transform 1 0 16652 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_181
timestamp 1667941163
transform 1 0 17756 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_193
timestamp 1667941163
transform 1 0 18860 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_205
timestamp 1667941163
transform 1 0 19964 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_217
timestamp 1667941163
transform 1 0 21068 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_223
timestamp 1667941163
transform 1 0 21620 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_225
timestamp 1667941163
transform 1 0 21804 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_237
timestamp 1667941163
transform 1 0 22908 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_77_249
timestamp 1667941163
transform 1 0 24012 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_77_278
timestamp 1667941163
transform 1 0 26680 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_77_281
timestamp 1667941163
transform 1 0 26956 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_77_286
timestamp 1667941163
transform 1 0 27416 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_77_293
timestamp 1667941163
transform 1 0 28060 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_78_3
timestamp 1667941163
transform 1 0 1380 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_9
timestamp 1667941163
transform 1 0 1932 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_78_13
timestamp 1667941163
transform 1 0 2300 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_78_21
timestamp 1667941163
transform 1 0 3036 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_78_26
timestamp 1667941163
transform 1 0 3496 0 1 44608
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_78_29
timestamp 1667941163
transform 1 0 3772 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_41
timestamp 1667941163
transform 1 0 4876 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_53
timestamp 1667941163
transform 1 0 5980 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_65
timestamp 1667941163
transform 1 0 7084 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_77
timestamp 1667941163
transform 1 0 8188 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_83
timestamp 1667941163
transform 1 0 8740 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_85
timestamp 1667941163
transform 1 0 8924 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_97
timestamp 1667941163
transform 1 0 10028 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_109
timestamp 1667941163
transform 1 0 11132 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_121
timestamp 1667941163
transform 1 0 12236 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_133
timestamp 1667941163
transform 1 0 13340 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_139
timestamp 1667941163
transform 1 0 13892 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_141
timestamp 1667941163
transform 1 0 14076 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_153
timestamp 1667941163
transform 1 0 15180 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_165
timestamp 1667941163
transform 1 0 16284 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_177
timestamp 1667941163
transform 1 0 17388 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_189
timestamp 1667941163
transform 1 0 18492 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_195
timestamp 1667941163
transform 1 0 19044 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_197
timestamp 1667941163
transform 1 0 19228 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_209
timestamp 1667941163
transform 1 0 20332 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_78_221
timestamp 1667941163
transform 1 0 21436 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_78_229
timestamp 1667941163
transform 1 0 22172 0 1 44608
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_78_235
timestamp 1667941163
transform 1 0 22724 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_78_247
timestamp 1667941163
transform 1 0 23828 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_78_251
timestamp 1667941163
transform 1 0 24196 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_78_253
timestamp 1667941163
transform 1 0 24380 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_78_258
timestamp 1667941163
transform 1 0 24840 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_265
timestamp 1667941163
transform 1 0 25484 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_272
timestamp 1667941163
transform 1 0 26128 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_78_297
timestamp 1667941163
transform 1 0 28428 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_79_3
timestamp 1667941163
transform 1 0 1380 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_7
timestamp 1667941163
transform 1 0 1748 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_79_11
timestamp 1667941163
transform 1 0 2116 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_18
timestamp 1667941163
transform 1 0 2760 0 -1 45696
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_79_25
timestamp 1667941163
transform 1 0 3404 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_37
timestamp 1667941163
transform 1 0 4508 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_49
timestamp 1667941163
transform 1 0 5612 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_55
timestamp 1667941163
transform 1 0 6164 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_57
timestamp 1667941163
transform 1 0 6348 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_69
timestamp 1667941163
transform 1 0 7452 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_81
timestamp 1667941163
transform 1 0 8556 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_79_96
timestamp 1667941163
transform 1 0 9936 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_79_103
timestamp 1667941163
transform 1 0 10580 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_79_111
timestamp 1667941163
transform 1 0 11316 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_79_113
timestamp 1667941163
transform 1 0 11500 0 -1 45696
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_79_118
timestamp 1667941163
transform 1 0 11960 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_130
timestamp 1667941163
transform 1 0 13064 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_142
timestamp 1667941163
transform 1 0 14168 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_154
timestamp 1667941163
transform 1 0 15272 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_79_166
timestamp 1667941163
transform 1 0 16376 0 -1 45696
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_79_169
timestamp 1667941163
transform 1 0 16652 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_181
timestamp 1667941163
transform 1 0 17756 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_79_193
timestamp 1667941163
transform 1 0 18860 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_197
timestamp 1667941163
transform 1 0 19228 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_79_201
timestamp 1667941163
transform 1 0 19596 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_208
timestamp 1667941163
transform 1 0 20240 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_79_215
timestamp 1667941163
transform 1 0 20884 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_79_223
timestamp 1667941163
transform 1 0 21620 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_79_225
timestamp 1667941163
transform 1 0 21804 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_229
timestamp 1667941163
transform 1 0 22172 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_79_233
timestamp 1667941163
transform 1 0 22540 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_79_240
timestamp 1667941163
transform 1 0 23184 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_79_248
timestamp 1667941163
transform 1 0 23920 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_79_253
timestamp 1667941163
transform 1 0 24380 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_79_278
timestamp 1667941163
transform 1 0 26680 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_79_281
timestamp 1667941163
transform 1 0 26956 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_79_286
timestamp 1667941163
transform 1 0 27416 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_290
timestamp 1667941163
transform 1 0 27784 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_79_294
timestamp 1667941163
transform 1 0 28152 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_298
timestamp 1667941163
transform 1 0 28520 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_80_3
timestamp 1667941163
transform 1 0 1380 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_80_26
timestamp 1667941163
transform 1 0 3496 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_80_29
timestamp 1667941163
transform 1 0 3772 0 1 45696
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_80_34
timestamp 1667941163
transform 1 0 4232 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_46
timestamp 1667941163
transform 1 0 5336 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_58
timestamp 1667941163
transform 1 0 6440 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_80_70
timestamp 1667941163
transform 1 0 7544 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_80_75
timestamp 1667941163
transform 1 0 8004 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_80_83
timestamp 1667941163
transform 1 0 8740 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_80_85
timestamp 1667941163
transform 1 0 8924 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_80_93
timestamp 1667941163
transform 1 0 9660 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_80_97
timestamp 1667941163
transform 1 0 10028 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_104
timestamp 1667941163
transform 1 0 10672 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_80_108
timestamp 1667941163
transform 1 0 11040 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_80_130
timestamp 1667941163
transform 1 0 13064 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_80_137
timestamp 1667941163
transform 1 0 13708 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_80_141
timestamp 1667941163
transform 1 0 14076 0 1 45696
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_80_148
timestamp 1667941163
transform 1 0 14720 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_80_160
timestamp 1667941163
transform 1 0 15824 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_80_164
timestamp 1667941163
transform 1 0 16192 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_168
timestamp 1667941163
transform 1 0 16560 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_80_180
timestamp 1667941163
transform 1 0 17664 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_80_191
timestamp 1667941163
transform 1 0 18676 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_80_195
timestamp 1667941163
transform 1 0 19044 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_80_197
timestamp 1667941163
transform 1 0 19228 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_80_220
timestamp 1667941163
transform 1 0 21344 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_80_249
timestamp 1667941163
transform 1 0 24012 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_80_253
timestamp 1667941163
transform 1 0 24380 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_80_258
timestamp 1667941163
transform 1 0 24840 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_80_287
timestamp 1667941163
transform 1 0 27508 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_294
timestamp 1667941163
transform 1 0 28152 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_80_298
timestamp 1667941163
transform 1 0 28520 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_81_3
timestamp 1667941163
transform 1 0 1380 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_81_9
timestamp 1667941163
transform 1 0 1932 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_16
timestamp 1667941163
transform 1 0 2576 0 -1 46784
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_81_41
timestamp 1667941163
transform 1 0 4876 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_81_53
timestamp 1667941163
transform 1 0 5980 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_81_57
timestamp 1667941163
transform 1 0 6348 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_63
timestamp 1667941163
transform 1 0 6900 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_81_85
timestamp 1667941163
transform 1 0 8924 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_81_110
timestamp 1667941163
transform 1 0 11224 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_81_113
timestamp 1667941163
transform 1 0 11500 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_81_140
timestamp 1667941163
transform 1 0 13984 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_81_165
timestamp 1667941163
transform 1 0 16284 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_81_169
timestamp 1667941163
transform 1 0 16652 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_81_192
timestamp 1667941163
transform 1 0 18768 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_81_217
timestamp 1667941163
transform 1 0 21068 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_223
timestamp 1667941163
transform 1 0 21620 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_81_225
timestamp 1667941163
transform 1 0 21804 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_81_248
timestamp 1667941163
transform 1 0 23920 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_81_256
timestamp 1667941163
transform 1 0 24656 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_81_278
timestamp 1667941163
transform 1 0 26680 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_81_281
timestamp 1667941163
transform 1 0 26956 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_81_286
timestamp 1667941163
transform 1 0 27416 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_81_293
timestamp 1667941163
transform 1 0 28060 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_82_3
timestamp 1667941163
transform 1 0 1380 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_82_26
timestamp 1667941163
transform 1 0 3496 0 1 46784
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_82_29
timestamp 1667941163
transform 1 0 3772 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_82_41
timestamp 1667941163
transform 1 0 4876 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_82_49
timestamp 1667941163
transform 1 0 5612 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_82_54
timestamp 1667941163
transform 1 0 6072 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_82_57
timestamp 1667941163
transform 1 0 6348 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_82_62
timestamp 1667941163
transform 1 0 6808 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_82_70
timestamp 1667941163
transform 1 0 7544 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_82_75
timestamp 1667941163
transform 1 0 8004 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_82_83
timestamp 1667941163
transform 1 0 8740 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_85
timestamp 1667941163
transform 1 0 8924 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_82_110
timestamp 1667941163
transform 1 0 11224 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_82_113
timestamp 1667941163
transform 1 0 11500 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_82_118
timestamp 1667941163
transform 1 0 11960 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_82_126
timestamp 1667941163
transform 1 0 12696 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_82_132
timestamp 1667941163
transform 1 0 13248 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_82_141
timestamp 1667941163
transform 1 0 14076 0 1 46784
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_82_148
timestamp 1667941163
transform 1 0 14720 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_82_160
timestamp 1667941163
transform 1 0 15824 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_82_169
timestamp 1667941163
transform 1 0 16652 0 1 46784
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_82_174
timestamp 1667941163
transform 1 0 17112 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_82_186
timestamp 1667941163
transform 1 0 18216 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_82_190
timestamp 1667941163
transform 1 0 18584 0 1 46784
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_82_197
timestamp 1667941163
transform 1 0 19228 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_82_209
timestamp 1667941163
transform 1 0 20332 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_82_215
timestamp 1667941163
transform 1 0 20884 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_82_222
timestamp 1667941163
transform 1 0 21528 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_82_225
timestamp 1667941163
transform 1 0 21804 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_82_250
timestamp 1667941163
transform 1 0 24104 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_82_253
timestamp 1667941163
transform 1 0 24380 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_82_278
timestamp 1667941163
transform 1 0 26680 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_82_281
timestamp 1667941163
transform 1 0 26956 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_82_286
timestamp 1667941163
transform 1 0 27416 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_82_293
timestamp 1667941163
transform 1 0 28060 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1667941163
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1667941163
transform -1 0 28888 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1667941163
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1667941163
transform -1 0 28888 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1667941163
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1667941163
transform -1 0 28888 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1667941163
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1667941163
transform -1 0 28888 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1667941163
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1667941163
transform -1 0 28888 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1667941163
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1667941163
transform -1 0 28888 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1667941163
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1667941163
transform -1 0 28888 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1667941163
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1667941163
transform -1 0 28888 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1667941163
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1667941163
transform -1 0 28888 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1667941163
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1667941163
transform -1 0 28888 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1667941163
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1667941163
transform -1 0 28888 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1667941163
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1667941163
transform -1 0 28888 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1667941163
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1667941163
transform -1 0 28888 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1667941163
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1667941163
transform -1 0 28888 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1667941163
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1667941163
transform -1 0 28888 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1667941163
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1667941163
transform -1 0 28888 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1667941163
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1667941163
transform -1 0 28888 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1667941163
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1667941163
transform -1 0 28888 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1667941163
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1667941163
transform -1 0 28888 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1667941163
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1667941163
transform -1 0 28888 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1667941163
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1667941163
transform -1 0 28888 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1667941163
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1667941163
transform -1 0 28888 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1667941163
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1667941163
transform -1 0 28888 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1667941163
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1667941163
transform -1 0 28888 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1667941163
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1667941163
transform -1 0 28888 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1667941163
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1667941163
transform -1 0 28888 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1667941163
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1667941163
transform -1 0 28888 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1667941163
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1667941163
transform -1 0 28888 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1667941163
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1667941163
transform -1 0 28888 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1667941163
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1667941163
transform -1 0 28888 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1667941163
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1667941163
transform -1 0 28888 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1667941163
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1667941163
transform -1 0 28888 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1667941163
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1667941163
transform -1 0 28888 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1667941163
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1667941163
transform -1 0 28888 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1667941163
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1667941163
transform -1 0 28888 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1667941163
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1667941163
transform -1 0 28888 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1667941163
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1667941163
transform -1 0 28888 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1667941163
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1667941163
transform -1 0 28888 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1667941163
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1667941163
transform -1 0 28888 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1667941163
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1667941163
transform -1 0 28888 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1667941163
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1667941163
transform -1 0 28888 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1667941163
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1667941163
transform -1 0 28888 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1667941163
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1667941163
transform -1 0 28888 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1667941163
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1667941163
transform -1 0 28888 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1667941163
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1667941163
transform -1 0 28888 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1667941163
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1667941163
transform -1 0 28888 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1667941163
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1667941163
transform -1 0 28888 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1667941163
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1667941163
transform -1 0 28888 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1667941163
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1667941163
transform -1 0 28888 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1667941163
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1667941163
transform -1 0 28888 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1667941163
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1667941163
transform -1 0 28888 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1667941163
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1667941163
transform -1 0 28888 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1667941163
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1667941163
transform -1 0 28888 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1667941163
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1667941163
transform -1 0 28888 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1667941163
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1667941163
transform -1 0 28888 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1667941163
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1667941163
transform -1 0 28888 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1667941163
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1667941163
transform -1 0 28888 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1667941163
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1667941163
transform -1 0 28888 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1667941163
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1667941163
transform -1 0 28888 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1667941163
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1667941163
transform -1 0 28888 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1667941163
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1667941163
transform -1 0 28888 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1667941163
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1667941163
transform -1 0 28888 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1667941163
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1667941163
transform -1 0 28888 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1667941163
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1667941163
transform -1 0 28888 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1667941163
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1667941163
transform -1 0 28888 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 1667941163
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 1667941163
transform -1 0 28888 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 1667941163
transform 1 0 1104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 1667941163
transform -1 0 28888 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_134
timestamp 1667941163
transform 1 0 1104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_135
timestamp 1667941163
transform -1 0 28888 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_136
timestamp 1667941163
transform 1 0 1104 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_137
timestamp 1667941163
transform -1 0 28888 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_138
timestamp 1667941163
transform 1 0 1104 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_139
timestamp 1667941163
transform -1 0 28888 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_140
timestamp 1667941163
transform 1 0 1104 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_141
timestamp 1667941163
transform -1 0 28888 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_142
timestamp 1667941163
transform 1 0 1104 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_143
timestamp 1667941163
transform -1 0 28888 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_144
timestamp 1667941163
transform 1 0 1104 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_145
timestamp 1667941163
transform -1 0 28888 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_146
timestamp 1667941163
transform 1 0 1104 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_147
timestamp 1667941163
transform -1 0 28888 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_148
timestamp 1667941163
transform 1 0 1104 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_149
timestamp 1667941163
transform -1 0 28888 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_150
timestamp 1667941163
transform 1 0 1104 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_151
timestamp 1667941163
transform -1 0 28888 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_152
timestamp 1667941163
transform 1 0 1104 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_153
timestamp 1667941163
transform -1 0 28888 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_154
timestamp 1667941163
transform 1 0 1104 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_155
timestamp 1667941163
transform -1 0 28888 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_156
timestamp 1667941163
transform 1 0 1104 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_157
timestamp 1667941163
transform -1 0 28888 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_158
timestamp 1667941163
transform 1 0 1104 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_159
timestamp 1667941163
transform -1 0 28888 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_160
timestamp 1667941163
transform 1 0 1104 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_161
timestamp 1667941163
transform -1 0 28888 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_162
timestamp 1667941163
transform 1 0 1104 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_163
timestamp 1667941163
transform -1 0 28888 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_164
timestamp 1667941163
transform 1 0 1104 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_165
timestamp 1667941163
transform -1 0 28888 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1667941163
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1667941163
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1667941163
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1667941163
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1667941163
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1667941163
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1667941163
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1667941163
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1667941163
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1667941163
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1667941163
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1667941163
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1667941163
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1667941163
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1667941163
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1667941163
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1667941163
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1667941163
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1667941163
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1667941163
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1667941163
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1667941163
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1667941163
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1667941163
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1667941163
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1667941163
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1667941163
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1667941163
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1667941163
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1667941163
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1667941163
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1667941163
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1667941163
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1667941163
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1667941163
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1667941163
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1667941163
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1667941163
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1667941163
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1667941163
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1667941163
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1667941163
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1667941163
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1667941163
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1667941163
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1667941163
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1667941163
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1667941163
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1667941163
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1667941163
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1667941163
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1667941163
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1667941163
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1667941163
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1667941163
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1667941163
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1667941163
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1667941163
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1667941163
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1667941163
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1667941163
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1667941163
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1667941163
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1667941163
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1667941163
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1667941163
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1667941163
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1667941163
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1667941163
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1667941163
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1667941163
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1667941163
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1667941163
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1667941163
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1667941163
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1667941163
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1667941163
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1667941163
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1667941163
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1667941163
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1667941163
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1667941163
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1667941163
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1667941163
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1667941163
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1667941163
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1667941163
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1667941163
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1667941163
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1667941163
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1667941163
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1667941163
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1667941163
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1667941163
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1667941163
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1667941163
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1667941163
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1667941163
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1667941163
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1667941163
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1667941163
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1667941163
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1667941163
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1667941163
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1667941163
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1667941163
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1667941163
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1667941163
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1667941163
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1667941163
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1667941163
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1667941163
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1667941163
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1667941163
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1667941163
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1667941163
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1667941163
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1667941163
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1667941163
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1667941163
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1667941163
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1667941163
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1667941163
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1667941163
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1667941163
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1667941163
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1667941163
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1667941163
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1667941163
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1667941163
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1667941163
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1667941163
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1667941163
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1667941163
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1667941163
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1667941163
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1667941163
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1667941163
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1667941163
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1667941163
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1667941163
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1667941163
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1667941163
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1667941163
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1667941163
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1667941163
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1667941163
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1667941163
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1667941163
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1667941163
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1667941163
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1667941163
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1667941163
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1667941163
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1667941163
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1667941163
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1667941163
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1667941163
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1667941163
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1667941163
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1667941163
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1667941163
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1667941163
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1667941163
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1667941163
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1667941163
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1667941163
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1667941163
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1667941163
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1667941163
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1667941163
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1667941163
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1667941163
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1667941163
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1667941163
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1667941163
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1667941163
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1667941163
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1667941163
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1667941163
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1667941163
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1667941163
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1667941163
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1667941163
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1667941163
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1667941163
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1667941163
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1667941163
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1667941163
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1667941163
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1667941163
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1667941163
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1667941163
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1667941163
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1667941163
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1667941163
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1667941163
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1667941163
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1667941163
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1667941163
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1667941163
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1667941163
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1667941163
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1667941163
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1667941163
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1667941163
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1667941163
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1667941163
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1667941163
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1667941163
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1667941163
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1667941163
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1667941163
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1667941163
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1667941163
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1667941163
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1667941163
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1667941163
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1667941163
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1667941163
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1667941163
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1667941163
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1667941163
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1667941163
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1667941163
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1667941163
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1667941163
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1667941163
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1667941163
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1667941163
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1667941163
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1667941163
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1667941163
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1667941163
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1667941163
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1667941163
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1667941163
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1667941163
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1667941163
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1667941163
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1667941163
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1667941163
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1667941163
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1667941163
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1667941163
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1667941163
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1667941163
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1667941163
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1667941163
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1667941163
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1667941163
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1667941163
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1667941163
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1667941163
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1667941163
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1667941163
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1667941163
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1667941163
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1667941163
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1667941163
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1667941163
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1667941163
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1667941163
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1667941163
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1667941163
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1667941163
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1667941163
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1667941163
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1667941163
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1667941163
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1667941163
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1667941163
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1667941163
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1667941163
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1667941163
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1667941163
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1667941163
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1667941163
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1667941163
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1667941163
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1667941163
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1667941163
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1667941163
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1667941163
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1667941163
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1667941163
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1667941163
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1667941163
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1667941163
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1667941163
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1667941163
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1667941163
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1667941163
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1667941163
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1667941163
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1667941163
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1667941163
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1667941163
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1667941163
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1667941163
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1667941163
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1667941163
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1667941163
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1667941163
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1667941163
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1667941163
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1667941163
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1667941163
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1667941163
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1667941163
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1667941163
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1667941163
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1667941163
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1667941163
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1667941163
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1667941163
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1667941163
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1667941163
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1667941163
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1667941163
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1667941163
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1667941163
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1667941163
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1667941163
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1667941163
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1667941163
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1667941163
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1667941163
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1667941163
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1667941163
transform 1 0 6256 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1667941163
transform 1 0 11408 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1667941163
transform 1 0 16560 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1667941163
transform 1 0 21712 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1667941163
transform 1 0 26864 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1667941163
transform 1 0 3680 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1667941163
transform 1 0 8832 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1667941163
transform 1 0 13984 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1667941163
transform 1 0 19136 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1667941163
transform 1 0 24288 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1667941163
transform 1 0 6256 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1667941163
transform 1 0 11408 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1667941163
transform 1 0 16560 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1667941163
transform 1 0 21712 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1667941163
transform 1 0 26864 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1667941163
transform 1 0 3680 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1667941163
transform 1 0 8832 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1667941163
transform 1 0 13984 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1667941163
transform 1 0 19136 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1667941163
transform 1 0 24288 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1667941163
transform 1 0 6256 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1667941163
transform 1 0 11408 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1667941163
transform 1 0 16560 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1667941163
transform 1 0 21712 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1667941163
transform 1 0 26864 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1667941163
transform 1 0 3680 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1667941163
transform 1 0 8832 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1667941163
transform 1 0 13984 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1667941163
transform 1 0 19136 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1667941163
transform 1 0 24288 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1667941163
transform 1 0 6256 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1667941163
transform 1 0 11408 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1667941163
transform 1 0 16560 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1667941163
transform 1 0 21712 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1667941163
transform 1 0 26864 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1667941163
transform 1 0 3680 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1667941163
transform 1 0 8832 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1667941163
transform 1 0 13984 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1667941163
transform 1 0 19136 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1667941163
transform 1 0 24288 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1667941163
transform 1 0 6256 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1667941163
transform 1 0 11408 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1667941163
transform 1 0 16560 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1667941163
transform 1 0 21712 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1667941163
transform 1 0 26864 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1667941163
transform 1 0 3680 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1667941163
transform 1 0 8832 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1667941163
transform 1 0 13984 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1667941163
transform 1 0 19136 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1667941163
transform 1 0 24288 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1667941163
transform 1 0 6256 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1667941163
transform 1 0 11408 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1667941163
transform 1 0 16560 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1667941163
transform 1 0 21712 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1667941163
transform 1 0 26864 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1667941163
transform 1 0 3680 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1667941163
transform 1 0 8832 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1667941163
transform 1 0 13984 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1667941163
transform 1 0 19136 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1667941163
transform 1 0 24288 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1667941163
transform 1 0 6256 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1667941163
transform 1 0 11408 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1667941163
transform 1 0 16560 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1667941163
transform 1 0 21712 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1667941163
transform 1 0 26864 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1667941163
transform 1 0 3680 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1667941163
transform 1 0 8832 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1667941163
transform 1 0 13984 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1667941163
transform 1 0 19136 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1667941163
transform 1 0 24288 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1667941163
transform 1 0 6256 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1667941163
transform 1 0 11408 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1667941163
transform 1 0 16560 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1667941163
transform 1 0 21712 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1667941163
transform 1 0 26864 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1667941163
transform 1 0 3680 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1667941163
transform 1 0 8832 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1667941163
transform 1 0 13984 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1667941163
transform 1 0 19136 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1667941163
transform 1 0 24288 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1667941163
transform 1 0 6256 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1667941163
transform 1 0 11408 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1667941163
transform 1 0 16560 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1667941163
transform 1 0 21712 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1667941163
transform 1 0 26864 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1667941163
transform 1 0 3680 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1667941163
transform 1 0 6256 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1667941163
transform 1 0 8832 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1667941163
transform 1 0 11408 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1667941163
transform 1 0 13984 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1667941163
transform 1 0 16560 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1667941163
transform 1 0 19136 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1667941163
transform 1 0 21712 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1667941163
transform 1 0 24288 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1667941163
transform 1 0 26864 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_8  _0475_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 1564 0 1 34816
box -38 -48 1050 592
use sky130_fd_sc_hd__buf_8  _0476_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 2392 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  _0477_
timestamp 1667941163
transform 1 0 3956 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0478_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 2024 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0479_
timestamp 1667941163
transform -1 0 2576 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0480_
timestamp 1667941163
transform -1 0 2116 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0481_
timestamp 1667941163
transform -1 0 27416 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0482_
timestamp 1667941163
transform -1 0 2576 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0483_
timestamp 1667941163
transform -1 0 28060 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0484_
timestamp 1667941163
transform 1 0 2392 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0485_
timestamp 1667941163
transform 1 0 27784 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0486_
timestamp 1667941163
transform 1 0 27968 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0487_
timestamp 1667941163
transform -1 0 13708 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _0488_
timestamp 1667941163
transform 1 0 27140 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0489_
timestamp 1667941163
transform 1 0 27692 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0490_
timestamp 1667941163
transform 1 0 25852 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0491_
timestamp 1667941163
transform -1 0 10672 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0492_
timestamp 1667941163
transform -1 0 10028 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0493_
timestamp 1667941163
transform -1 0 4232 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0494_
timestamp 1667941163
transform -1 0 2392 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0495_
timestamp 1667941163
transform 1 0 27784 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0496_
timestamp 1667941163
transform 1 0 2484 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0497_
timestamp 1667941163
transform 1 0 18400 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0498_
timestamp 1667941163
transform 1 0 10580 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _0499_
timestamp 1667941163
transform -1 0 2852 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0500_
timestamp 1667941163
transform -1 0 27508 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0501_
timestamp 1667941163
transform -1 0 2392 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0502_
timestamp 1667941163
transform -1 0 6072 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0503_
timestamp 1667941163
transform 1 0 28060 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0504_
timestamp 1667941163
transform 1 0 27876 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0505_
timestamp 1667941163
transform 1 0 28152 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0506_
timestamp 1667941163
transform -1 0 2116 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0507_
timestamp 1667941163
transform -1 0 8188 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0508_
timestamp 1667941163
transform -1 0 4876 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0509_
timestamp 1667941163
transform 1 0 2392 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _0510_
timestamp 1667941163
transform 1 0 3956 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0511_
timestamp 1667941163
transform -1 0 27508 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0512_
timestamp 1667941163
transform -1 0 2576 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0513_
timestamp 1667941163
transform 1 0 27692 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0514_
timestamp 1667941163
transform -1 0 20332 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0515_
timestamp 1667941163
transform -1 0 23184 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0516_
timestamp 1667941163
transform -1 0 27416 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0517_
timestamp 1667941163
transform 1 0 27876 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0518_
timestamp 1667941163
transform -1 0 4232 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0519_
timestamp 1667941163
transform -1 0 27508 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0520_
timestamp 1667941163
transform -1 0 27508 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _0521_
timestamp 1667941163
transform -1 0 3496 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0522_
timestamp 1667941163
transform -1 0 2116 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0523_
timestamp 1667941163
transform 1 0 20608 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0524_
timestamp 1667941163
transform 1 0 12788 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0525_
timestamp 1667941163
transform 1 0 27140 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0526_
timestamp 1667941163
transform -1 0 2116 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0527_
timestamp 1667941163
transform 1 0 1748 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0528_
timestamp 1667941163
transform 1 0 1748 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0529_
timestamp 1667941163
transform 1 0 27140 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0530_
timestamp 1667941163
transform 1 0 27232 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0531_
timestamp 1667941163
transform -1 0 2576 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _0532_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 5428 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0533_
timestamp 1667941163
transform 1 0 5336 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0534_
timestamp 1667941163
transform 1 0 25760 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0535_
timestamp 1667941163
transform -1 0 26404 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0536_
timestamp 1667941163
transform 1 0 5980 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0537_
timestamp 1667941163
transform 1 0 2944 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0538_
timestamp 1667941163
transform 1 0 16744 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0539_
timestamp 1667941163
transform 1 0 3956 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0540_
timestamp 1667941163
transform 1 0 25852 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0541_
timestamp 1667941163
transform -1 0 2484 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0542_
timestamp 1667941163
transform 1 0 27140 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _0543_
timestamp 1667941163
transform 1 0 4692 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0544_
timestamp 1667941163
transform -1 0 2024 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0545_
timestamp 1667941163
transform 1 0 25852 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0546_
timestamp 1667941163
transform 1 0 8372 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0547_
timestamp 1667941163
transform -1 0 27416 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0548_
timestamp 1667941163
transform 1 0 14444 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0549_
timestamp 1667941163
transform -1 0 27416 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0550_
timestamp 1667941163
transform -1 0 10028 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0551_
timestamp 1667941163
transform 1 0 28060 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0552_
timestamp 1667941163
transform -1 0 27416 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0553_
timestamp 1667941163
transform -1 0 2668 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _0554_
timestamp 1667941163
transform -1 0 5060 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0555_
timestamp 1667941163
transform 1 0 27968 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0556_
timestamp 1667941163
transform -1 0 27416 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0557_
timestamp 1667941163
transform -1 0 2024 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0558_
timestamp 1667941163
transform -1 0 28060 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0559_
timestamp 1667941163
transform -1 0 2668 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0560_
timestamp 1667941163
transform -1 0 4416 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0561_
timestamp 1667941163
transform 1 0 28060 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0562_
timestamp 1667941163
transform -1 0 22540 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0563_
timestamp 1667941163
transform -1 0 2208 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0564_
timestamp 1667941163
transform 1 0 19320 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _0565_
timestamp 1667941163
transform 1 0 3956 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0566_
timestamp 1667941163
transform -1 0 25484 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0567_
timestamp 1667941163
transform 1 0 16284 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0568_
timestamp 1667941163
transform 1 0 5152 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0569_
timestamp 1667941163
transform -1 0 2300 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0570_
timestamp 1667941163
transform 1 0 23828 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0571_
timestamp 1667941163
transform 1 0 25852 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0572_
timestamp 1667941163
transform 1 0 27600 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0573_
timestamp 1667941163
transform -1 0 8004 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0574_
timestamp 1667941163
transform 1 0 27784 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0575_
timestamp 1667941163
transform -1 0 2392 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _0576_
timestamp 1667941163
transform 1 0 3220 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0577_
timestamp 1667941163
transform 1 0 14260 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0578_
timestamp 1667941163
transform 1 0 10672 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0579_
timestamp 1667941163
transform 1 0 27324 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0580_
timestamp 1667941163
transform 1 0 11960 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0581_
timestamp 1667941163
transform 1 0 21988 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0582_
timestamp 1667941163
transform 1 0 25852 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0583_
timestamp 1667941163
transform 1 0 17112 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0584_
timestamp 1667941163
transform 1 0 25852 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0585_
timestamp 1667941163
transform -1 0 4232 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0586_
timestamp 1667941163
transform -1 0 11960 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0587_
timestamp 1667941163
transform -1 0 3128 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0588_
timestamp 1667941163
transform -1 0 3312 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0589_
timestamp 1667941163
transform 1 0 27968 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0590_
timestamp 1667941163
transform -1 0 27416 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0591_
timestamp 1667941163
transform -1 0 27508 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0592_
timestamp 1667941163
transform 1 0 20424 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0593_
timestamp 1667941163
transform 1 0 26404 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _0594_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 26128 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _0595_
timestamp 1667941163
transform 1 0 20608 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _0596_
timestamp 1667941163
transform 1 0 22080 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0597_
timestamp 1667941163
transform -1 0 18032 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0598_
timestamp 1667941163
transform 1 0 18308 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__a22oi_1  _0599_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 15916 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0600_
timestamp 1667941163
transform 1 0 19872 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0601_
timestamp 1667941163
transform 1 0 19412 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _0602_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 20608 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0603_
timestamp 1667941163
transform -1 0 23184 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _0604_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 21252 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0605_
timestamp 1667941163
transform -1 0 24104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _0606_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 20148 0 -1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0607_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 22172 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0608_
timestamp 1667941163
transform -1 0 17848 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _0609_
timestamp 1667941163
transform -1 0 17480 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0610_
timestamp 1667941163
transform -1 0 19596 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _0611_
timestamp 1667941163
transform -1 0 18584 0 -1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0612_
timestamp 1667941163
transform 1 0 19412 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _0613_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 18216 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _0614_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 20240 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _0615_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 18952 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0616_
timestamp 1667941163
transform -1 0 18492 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _0617_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 18032 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__a32o_1  _0618_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 19504 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0619_
timestamp 1667941163
transform 1 0 17848 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0620_
timestamp 1667941163
transform 1 0 19136 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0621_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 19872 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0622_
timestamp 1667941163
transform 1 0 17664 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _0623_
timestamp 1667941163
transform -1 0 18768 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__a21bo_1  _0624_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 18308 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__a211oi_1  _0625_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 17756 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0626_
timestamp 1667941163
transform 1 0 18492 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _0627_
timestamp 1667941163
transform -1 0 18584 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _0628_
timestamp 1667941163
transform 1 0 19688 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0629_
timestamp 1667941163
transform 1 0 18492 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _0630_
timestamp 1667941163
transform 1 0 18676 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a21boi_2  _0631_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 18216 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _0632_
timestamp 1667941163
transform 1 0 17848 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _0633_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 27140 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _0634_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 27692 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _0635_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 27600 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _0636_
timestamp 1667941163
transform 1 0 23184 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _0637_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 22172 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0638_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 21528 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0639_
timestamp 1667941163
transform -1 0 21528 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_2  _0640_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 19504 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _0641_
timestamp 1667941163
transform 1 0 21436 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__or3b_1  _0642_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 21528 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _0643_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 22264 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _0644_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 19412 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0645_
timestamp 1667941163
transform 1 0 14352 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0646_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 19228 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_2  _0647_
timestamp 1667941163
transform 1 0 21988 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _0648_
timestamp 1667941163
transform 1 0 13340 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _0649_
timestamp 1667941163
transform 1 0 19504 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _0650_
timestamp 1667941163
transform -1 0 13984 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0651_
timestamp 1667941163
transform -1 0 12972 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0652_
timestamp 1667941163
transform 1 0 12512 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _0653_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 14168 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_1  _0654_
timestamp 1667941163
transform -1 0 15732 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0655_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 14260 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__or2b_1  _0656_
timestamp 1667941163
transform -1 0 15180 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0657_
timestamp 1667941163
transform -1 0 15180 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__o21bai_2  _0658_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 12236 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _0659_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 13524 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0660_
timestamp 1667941163
transform 1 0 14536 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_2  _0661_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 14260 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _0662_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 14260 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0663_
timestamp 1667941163
transform -1 0 15916 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0664_
timestamp 1667941163
transform -1 0 15456 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0665_
timestamp 1667941163
transform -1 0 25484 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _0666_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 13248 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _0667_
timestamp 1667941163
transform 1 0 12604 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__clkinv_2  _0668_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 25944 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _0669_
timestamp 1667941163
transform 1 0 24104 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0670_
timestamp 1667941163
transform -1 0 22816 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0671_
timestamp 1667941163
transform -1 0 3036 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0672_
timestamp 1667941163
transform 1 0 24564 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0673_
timestamp 1667941163
transform -1 0 24472 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0674_
timestamp 1667941163
transform -1 0 24932 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_2  _0675_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 24564 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_4  _0676_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 24380 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__or2_2  _0677_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 24196 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _0678_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 24564 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__o221ai_1  _0679_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 25208 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0680_
timestamp 1667941163
transform -1 0 26312 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _0681_
timestamp 1667941163
transform 1 0 24656 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _0682_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 25760 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _0683_
timestamp 1667941163
transform -1 0 24012 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0684_
timestamp 1667941163
transform 1 0 24196 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _0685_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 23552 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__o32a_1  _0686_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 25300 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0687_
timestamp 1667941163
transform 1 0 25116 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _0688_
timestamp 1667941163
transform -1 0 26128 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _0689_
timestamp 1667941163
transform -1 0 26680 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _0690_
timestamp 1667941163
transform -1 0 26680 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0691_
timestamp 1667941163
transform 1 0 25392 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0692_
timestamp 1667941163
transform 1 0 24564 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0693_
timestamp 1667941163
transform -1 0 25760 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _0694_
timestamp 1667941163
transform 1 0 25208 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _0695_
timestamp 1667941163
transform 1 0 24656 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0696_
timestamp 1667941163
transform -1 0 25944 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0697_
timestamp 1667941163
transform 1 0 24840 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0698_
timestamp 1667941163
transform -1 0 25668 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0699_
timestamp 1667941163
transform 1 0 26312 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _0700_
timestamp 1667941163
transform 1 0 27140 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0701_
timestamp 1667941163
transform -1 0 26128 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0702_
timestamp 1667941163
transform -1 0 26220 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0703_
timestamp 1667941163
transform -1 0 25392 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0704_
timestamp 1667941163
transform -1 0 25484 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _0705_
timestamp 1667941163
transform -1 0 26220 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _0706_
timestamp 1667941163
transform 1 0 25116 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__o211ai_1  _0707_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 25300 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _0708_
timestamp 1667941163
transform -1 0 26220 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _0709_
timestamp 1667941163
transform -1 0 24012 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _0710_
timestamp 1667941163
transform 1 0 23920 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _0711_
timestamp 1667941163
transform 1 0 23828 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0712_
timestamp 1667941163
transform 1 0 23368 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__nor3_1  _0713_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 23000 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _0714_
timestamp 1667941163
transform 1 0 21988 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0715_
timestamp 1667941163
transform -1 0 21528 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0716_
timestamp 1667941163
transform -1 0 20700 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0717_
timestamp 1667941163
transform -1 0 21344 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _0718_
timestamp 1667941163
transform 1 0 19872 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0719_
timestamp 1667941163
transform -1 0 18952 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0720_
timestamp 1667941163
transform 1 0 18492 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0721_
timestamp 1667941163
transform 1 0 21068 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0722_
timestamp 1667941163
transform 1 0 20148 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0723_
timestamp 1667941163
transform 1 0 20240 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0724_
timestamp 1667941163
transform 1 0 19872 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0725_
timestamp 1667941163
transform -1 0 19872 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0726_
timestamp 1667941163
transform -1 0 19688 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0727_
timestamp 1667941163
transform 1 0 21988 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0728_
timestamp 1667941163
transform 1 0 20884 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0729_
timestamp 1667941163
transform 1 0 20976 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0730_
timestamp 1667941163
transform 1 0 20608 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0731_
timestamp 1667941163
transform -1 0 19872 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0732_
timestamp 1667941163
transform -1 0 18952 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0733_
timestamp 1667941163
transform 1 0 19412 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0734_
timestamp 1667941163
transform 1 0 18400 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0735_
timestamp 1667941163
transform 1 0 18584 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0736_
timestamp 1667941163
transform 1 0 19504 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0737_
timestamp 1667941163
transform 1 0 18492 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0738_
timestamp 1667941163
transform -1 0 18952 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0739_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 16836 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _0740_
timestamp 1667941163
transform -1 0 16376 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _0741_
timestamp 1667941163
transform 1 0 16836 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0742_
timestamp 1667941163
transform 1 0 16836 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0743_
timestamp 1667941163
transform -1 0 16376 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _0744_
timestamp 1667941163
transform 1 0 16100 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0745_
timestamp 1667941163
transform -1 0 17204 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0746_
timestamp 1667941163
transform 1 0 23092 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _0747_
timestamp 1667941163
transform 1 0 23092 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0748_
timestamp 1667941163
transform 1 0 22448 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0749_
timestamp 1667941163
transform 1 0 23920 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _0750_
timestamp 1667941163
transform -1 0 23736 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0751_
timestamp 1667941163
transform 1 0 23184 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0752_
timestamp 1667941163
transform -1 0 17480 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0753_
timestamp 1667941163
transform 1 0 16836 0 -1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0754_
timestamp 1667941163
transform 1 0 17572 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0755_
timestamp 1667941163
transform -1 0 16376 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _0756_
timestamp 1667941163
transform -1 0 16376 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0757_
timestamp 1667941163
transform -1 0 16836 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0758_
timestamp 1667941163
transform -1 0 16560 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0759_
timestamp 1667941163
transform 1 0 15916 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0760_
timestamp 1667941163
transform -1 0 17204 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0761_
timestamp 1667941163
transform -1 0 16008 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _0762_
timestamp 1667941163
transform 1 0 15548 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0763_
timestamp 1667941163
transform -1 0 17112 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0764_
timestamp 1667941163
transform 1 0 16836 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0765_
timestamp 1667941163
transform 1 0 16468 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0766_
timestamp 1667941163
transform 1 0 17296 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0767_
timestamp 1667941163
transform 1 0 27140 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0768_
timestamp 1667941163
transform 1 0 26036 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0769_
timestamp 1667941163
transform 1 0 27140 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0770_
timestamp 1667941163
transform -1 0 16192 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _0771_
timestamp 1667941163
transform -1 0 16192 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0772_
timestamp 1667941163
transform -1 0 16652 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0773_
timestamp 1667941163
transform 1 0 25852 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0774_
timestamp 1667941163
transform -1 0 26036 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0775_
timestamp 1667941163
transform -1 0 25852 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0776_
timestamp 1667941163
transform -1 0 21344 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0777_
timestamp 1667941163
transform -1 0 21068 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0778_
timestamp 1667941163
transform -1 0 22448 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__a21boi_1  _0779_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 22816 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _0780_
timestamp 1667941163
transform -1 0 23184 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _0781_
timestamp 1667941163
transform 1 0 22356 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__a21boi_1  _0782_
timestamp 1667941163
transform 1 0 20976 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _0783_
timestamp 1667941163
transform -1 0 22816 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _0784_
timestamp 1667941163
transform 1 0 20792 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__a21boi_1  _0785_
timestamp 1667941163
transform 1 0 21160 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _0786_
timestamp 1667941163
transform -1 0 22448 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _0787_
timestamp 1667941163
transform 1 0 20976 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__a21boi_1  _0788_
timestamp 1667941163
transform 1 0 20884 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _0789_
timestamp 1667941163
transform -1 0 22448 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _0790_
timestamp 1667941163
transform 1 0 20792 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _0791_
timestamp 1667941163
transform -1 0 23276 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _0792_
timestamp 1667941163
transform -1 0 23828 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _0793_
timestamp 1667941163
transform -1 0 25024 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_1  _0794_
timestamp 1667941163
transform 1 0 24104 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _0795_
timestamp 1667941163
transform 1 0 23184 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0796_
timestamp 1667941163
transform 1 0 23000 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__o21ba_1  _0797_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 23736 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _0798_
timestamp 1667941163
transform 1 0 22908 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0799_
timestamp 1667941163
transform 1 0 23368 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _0800_
timestamp 1667941163
transform 1 0 22356 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a41o_1  _0801_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 22264 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__and2b_1  _0802_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 22540 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0803_
timestamp 1667941163
transform 1 0 21804 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nand4_1  _0804_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 23736 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _0805_
timestamp 1667941163
transform -1 0 24012 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0806_
timestamp 1667941163
transform -1 0 25024 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0807_
timestamp 1667941163
transform -1 0 24840 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0808_
timestamp 1667941163
transform 1 0 19504 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _0809_
timestamp 1667941163
transform -1 0 19688 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0810_
timestamp 1667941163
transform -1 0 21528 0 -1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0811_
timestamp 1667941163
transform 1 0 18492 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0812_
timestamp 1667941163
transform 1 0 16836 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _0813_
timestamp 1667941163
transform 1 0 20424 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _0814_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 19964 0 1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _0815_
timestamp 1667941163
transform 1 0 20516 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0816_
timestamp 1667941163
transform 1 0 21804 0 1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0817_
timestamp 1667941163
transform -1 0 21436 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0818_
timestamp 1667941163
transform 1 0 20976 0 1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0819_
timestamp 1667941163
transform -1 0 22264 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _0820_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 20700 0 -1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0821_
timestamp 1667941163
transform -1 0 19320 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0822_
timestamp 1667941163
transform 1 0 19596 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _0823_
timestamp 1667941163
transform 1 0 18492 0 1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0824_
timestamp 1667941163
transform -1 0 19228 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0825_
timestamp 1667941163
transform -1 0 18676 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _0826_
timestamp 1667941163
transform -1 0 20056 0 1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0827_
timestamp 1667941163
transform 1 0 18032 0 1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0828_
timestamp 1667941163
transform -1 0 18676 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0829_
timestamp 1667941163
transform -1 0 15364 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0830_
timestamp 1667941163
transform 1 0 15272 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0831_
timestamp 1667941163
transform 1 0 15732 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0832_
timestamp 1667941163
transform -1 0 17112 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _0833_
timestamp 1667941163
transform -1 0 16284 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0834_
timestamp 1667941163
transform 1 0 15824 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0835_
timestamp 1667941163
transform 1 0 15824 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0836_
timestamp 1667941163
transform -1 0 16376 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0837_
timestamp 1667941163
transform 1 0 15824 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0838_
timestamp 1667941163
transform 1 0 15824 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _0839_
timestamp 1667941163
transform 1 0 15732 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _0840_
timestamp 1667941163
transform -1 0 16836 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0841_
timestamp 1667941163
transform -1 0 16192 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0842_
timestamp 1667941163
transform 1 0 15916 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _0843_
timestamp 1667941163
transform 1 0 15732 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _0844_
timestamp 1667941163
transform -1 0 16376 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0845_
timestamp 1667941163
transform -1 0 16376 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0846_
timestamp 1667941163
transform 1 0 16836 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _0847_
timestamp 1667941163
transform 1 0 15640 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _0848_
timestamp 1667941163
transform -1 0 17020 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0849_
timestamp 1667941163
transform 1 0 16008 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0850_
timestamp 1667941163
transform 1 0 16100 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0851_
timestamp 1667941163
transform 1 0 16836 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0852_
timestamp 1667941163
transform -1 0 17940 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a21boi_1  _0853_
timestamp 1667941163
transform 1 0 16836 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _0854_
timestamp 1667941163
transform -1 0 23828 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _0855_
timestamp 1667941163
transform 1 0 22816 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _0856_
timestamp 1667941163
transform -1 0 24840 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0857_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 22540 0 1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _0858_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 21988 0 -1 32640
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _0859_
timestamp 1667941163
transform 1 0 21896 0 1 26112
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _0860_
timestamp 1667941163
transform 1 0 25116 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _0861_
timestamp 1667941163
transform 1 0 25760 0 1 19584
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _0862_
timestamp 1667941163
transform 1 0 25208 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0863_
timestamp 1667941163
transform -1 0 26680 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0864_
timestamp 1667941163
transform 1 0 26036 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0865_
timestamp 1667941163
transform 1 0 22080 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0866_
timestamp 1667941163
transform 1 0 20608 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0867_
timestamp 1667941163
transform 1 0 18032 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0868_
timestamp 1667941163
transform -1 0 20700 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0869_
timestamp 1667941163
transform 1 0 19412 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0870_
timestamp 1667941163
transform 1 0 20792 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0871_
timestamp 1667941163
transform 1 0 18768 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0872_
timestamp 1667941163
transform 1 0 18216 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0873_
timestamp 1667941163
transform 1 0 18676 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0874_
timestamp 1667941163
transform -1 0 26680 0 -1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0875_
timestamp 1667941163
transform 1 0 25208 0 -1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0876_
timestamp 1667941163
transform -1 0 26128 0 -1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0877_
timestamp 1667941163
transform 1 0 16744 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0878_
timestamp 1667941163
transform 1 0 16836 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0879_
timestamp 1667941163
transform 1 0 22356 0 -1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0880_
timestamp 1667941163
transform 1 0 22632 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0881_
timestamp 1667941163
transform 1 0 16836 0 1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0882_
timestamp 1667941163
transform 1 0 16836 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0883_
timestamp 1667941163
transform 1 0 16836 0 -1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0884_
timestamp 1667941163
transform 1 0 16652 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0885_
timestamp 1667941163
transform 1 0 16836 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0886_
timestamp 1667941163
transform 1 0 26128 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0887_
timestamp 1667941163
transform 1 0 16836 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0888_
timestamp 1667941163
transform -1 0 26128 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_4  _0889_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 20516 0 1 29376
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_1  _0890_
timestamp 1667941163
transform 1 0 21804 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0891_
timestamp 1667941163
transform 1 0 19964 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0892_
timestamp 1667941163
transform -1 0 21528 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0893_
timestamp 1667941163
transform -1 0 21160 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0894_
timestamp 1667941163
transform 1 0 24104 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0895_
timestamp 1667941163
transform -1 0 24656 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0896_
timestamp 1667941163
transform 1 0 21620 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0897_
timestamp 1667941163
transform -1 0 26496 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0898_
timestamp 1667941163
transform 1 0 19412 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0899_
timestamp 1667941163
transform 1 0 20056 0 1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0900_
timestamp 1667941163
transform -1 0 22724 0 1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0901_
timestamp 1667941163
transform 1 0 19412 0 1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0902_
timestamp 1667941163
transform 1 0 18676 0 -1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0903_
timestamp 1667941163
transform 1 0 16928 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0904_
timestamp 1667941163
transform 1 0 16836 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0905_
timestamp 1667941163
transform 1 0 16836 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0906_
timestamp 1667941163
transform 1 0 16652 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0907_
timestamp 1667941163
transform 1 0 16928 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0908_
timestamp 1667941163
transform -1 0 18308 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0909_
timestamp 1667941163
transform 1 0 17204 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0910_
timestamp 1667941163
transform 1 0 22540 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _0911_
timestamp 1667941163
transform 1 0 24196 0 -1 35904
box -38 -48 1602 592
use sky130_fd_sc_hd__conb_1  _1012__17 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 6808 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1012_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 6532 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1013__18
timestamp 1667941163
transform 1 0 1748 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1013_
timestamp 1667941163
transform -1 0 3588 0 -1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1014__19
timestamp 1667941163
transform 1 0 16100 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1014_
timestamp 1667941163
transform 1 0 16836 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1015__20
timestamp 1667941163
transform 1 0 3128 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1015_
timestamp 1667941163
transform -1 0 4968 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1016__21
timestamp 1667941163
transform -1 0 27416 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1016_
timestamp 1667941163
transform 1 0 26496 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1017__22
timestamp 1667941163
transform -1 0 3128 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1017_
timestamp 1667941163
transform 1 0 2852 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1018__23
timestamp 1667941163
transform -1 0 27416 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1018_
timestamp 1667941163
transform 1 0 26496 0 1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1019__24
timestamp 1667941163
transform -1 0 5520 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1019_
timestamp 1667941163
transform -1 0 3588 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1020__25
timestamp 1667941163
transform -1 0 28152 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1020_
timestamp 1667941163
transform 1 0 26496 0 1 39168
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1021__26
timestamp 1667941163
transform -1 0 28060 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1021_
timestamp 1667941163
transform -1 0 26680 0 -1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1022__27
timestamp 1667941163
transform -1 0 28152 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1022_
timestamp 1667941163
transform 1 0 26496 0 1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1023__28
timestamp 1667941163
transform -1 0 17664 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1023_
timestamp 1667941163
transform 1 0 17020 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1024__29
timestamp 1667941163
transform -1 0 26128 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1024_
timestamp 1667941163
transform 1 0 25852 0 1 43520
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1025__30
timestamp 1667941163
transform -1 0 3496 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1025_
timestamp 1667941163
transform 1 0 3128 0 -1 44608
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1026__31
timestamp 1667941163
transform -1 0 11960 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1026_
timestamp 1667941163
transform 1 0 11132 0 1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1027__32
timestamp 1667941163
transform 1 0 3956 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1027_
timestamp 1667941163
transform -1 0 4324 0 -1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1028__33
timestamp 1667941163
transform -1 0 28152 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1028_
timestamp 1667941163
transform 1 0 26496 0 1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1029__34
timestamp 1667941163
transform -1 0 28060 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1029_
timestamp 1667941163
transform 1 0 26496 0 1 38080
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1030__35
timestamp 1667941163
transform 1 0 2392 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1030_
timestamp 1667941163
transform 1 0 2760 0 -1 39168
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1031_
timestamp 1667941163
transform 1 0 26496 0 1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1031__36
timestamp 1667941163
transform 1 0 26404 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1032_
timestamp 1667941163
transform 1 0 1564 0 1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1032__37
timestamp 1667941163
transform -1 0 1932 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1033_
timestamp 1667941163
transform 1 0 26496 0 1 44608
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1033__38
timestamp 1667941163
transform -1 0 28060 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1034__39
timestamp 1667941163
transform -1 0 14720 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1034_
timestamp 1667941163
transform 1 0 14352 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1035__40
timestamp 1667941163
transform -1 0 9384 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1035_
timestamp 1667941163
transform 1 0 8924 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1036__41
timestamp 1667941163
transform 1 0 27784 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1036_
timestamp 1667941163
transform -1 0 28428 0 1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1037__42
timestamp 1667941163
transform 1 0 2944 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1037_
timestamp 1667941163
transform -1 0 3496 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1038_
timestamp 1667941163
transform -1 0 28428 0 1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1038__43
timestamp 1667941163
transform 1 0 27876 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1039__44
timestamp 1667941163
transform -1 0 2024 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1039_
timestamp 1667941163
transform 1 0 1564 0 1 38080
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1040_
timestamp 1667941163
transform -1 0 28428 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1040__45
timestamp 1667941163
transform 1 0 27876 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1041__46
timestamp 1667941163
transform -1 0 4324 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1041_
timestamp 1667941163
transform 1 0 3956 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1042__47
timestamp 1667941163
transform 1 0 27416 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1042_
timestamp 1667941163
transform -1 0 28428 0 1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1043_
timestamp 1667941163
transform 1 0 24748 0 1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1043__48
timestamp 1667941163
transform 1 0 24564 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1044__49
timestamp 1667941163
transform -1 0 27416 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1044_
timestamp 1667941163
transform 1 0 26496 0 1 40256
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1045__50
timestamp 1667941163
transform -1 0 17112 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1045_
timestamp 1667941163
transform 1 0 16836 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1046__51
timestamp 1667941163
transform 1 0 4416 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1046_
timestamp 1667941163
transform 1 0 5060 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1047_
timestamp 1667941163
transform 1 0 1656 0 -1 34816
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1047__52
timestamp 1667941163
transform -1 0 2024 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1048__53
timestamp 1667941163
transform -1 0 27416 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1048_
timestamp 1667941163
transform 1 0 26496 0 1 34816
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1049__54
timestamp 1667941163
transform -1 0 8004 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1049_
timestamp 1667941163
transform 1 0 6992 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1050_
timestamp 1667941163
transform 1 0 24748 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1050__55
timestamp 1667941163
transform 1 0 24104 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1051__56
timestamp 1667941163
transform -1 0 2024 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1051_
timestamp 1667941163
transform 1 0 1656 0 -1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1052__57
timestamp 1667941163
transform -1 0 14628 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1052_
timestamp 1667941163
transform 1 0 14260 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1053_
timestamp 1667941163
transform -1 0 13248 0 1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1054_
timestamp 1667941163
transform 1 0 26496 0 1 31552
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1055_
timestamp 1667941163
transform 1 0 11868 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1056_
timestamp 1667941163
transform -1 0 7912 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1057_
timestamp 1667941163
transform 1 0 25668 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1058_
timestamp 1667941163
transform 1 0 25760 0 1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1059_
timestamp 1667941163
transform -1 0 11040 0 1 30464
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1060_
timestamp 1667941163
transform 1 0 26220 0 1 33728
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1061__58
timestamp 1667941163
transform 1 0 27140 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1061_
timestamp 1667941163
transform -1 0 27508 0 1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1062_
timestamp 1667941163
transform 1 0 26496 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1062__59
timestamp 1667941163
transform -1 0 28060 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1063_
timestamp 1667941163
transform 1 0 1656 0 -1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1063__60
timestamp 1667941163
transform -1 0 2024 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1064__61
timestamp 1667941163
transform 1 0 21252 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1064_
timestamp 1667941163
transform 1 0 22080 0 1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1065__62
timestamp 1667941163
transform -1 0 1932 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1065_
timestamp 1667941163
transform 1 0 1656 0 -1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1066__63
timestamp 1667941163
transform -1 0 24840 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1066_
timestamp 1667941163
transform 1 0 24288 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1067__64
timestamp 1667941163
transform 1 0 27692 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1067_
timestamp 1667941163
transform -1 0 28428 0 1 29376
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1068__65
timestamp 1667941163
transform 1 0 21344 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1068_
timestamp 1667941163
transform 1 0 21988 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1069__66
timestamp 1667941163
transform -1 0 20240 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1069_
timestamp 1667941163
transform 1 0 19412 0 1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1070__67
timestamp 1667941163
transform -1 0 1840 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1070_
timestamp 1667941163
transform 1 0 1564 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1071__68
timestamp 1667941163
transform 1 0 20608 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1071_
timestamp 1667941163
transform 1 0 21988 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1072__69
timestamp 1667941163
transform -1 0 13156 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1072_
timestamp 1667941163
transform 1 0 12788 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1073_
timestamp 1667941163
transform 1 0 26496 0 1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1073__70
timestamp 1667941163
transform -1 0 27416 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1074__71
timestamp 1667941163
transform -1 0 2024 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1074_
timestamp 1667941163
transform 1 0 1656 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1075__72
timestamp 1667941163
transform -1 0 1932 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1075_
timestamp 1667941163
transform 1 0 1656 0 -1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1076__73
timestamp 1667941163
transform -1 0 4232 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1076_
timestamp 1667941163
transform -1 0 3588 0 -1 38080
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1077__74
timestamp 1667941163
transform -1 0 28152 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1077_
timestamp 1667941163
transform 1 0 26496 0 1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1078__75
timestamp 1667941163
transform -1 0 28428 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1078_
timestamp 1667941163
transform -1 0 26680 0 -1 42432
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1079_
timestamp 1667941163
transform 1 0 26496 0 1 41344
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1079__76
timestamp 1667941163
transform -1 0 28152 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1080__77
timestamp 1667941163
transform 1 0 2300 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1080_
timestamp 1667941163
transform 1 0 2944 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1081__78
timestamp 1667941163
transform -1 0 28152 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1081_
timestamp 1667941163
transform -1 0 26680 0 -1 44608
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1082_
timestamp 1667941163
transform 1 0 20424 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1082__79
timestamp 1667941163
transform -1 0 20792 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1083_
timestamp 1667941163
transform 1 0 26496 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1083__80
timestamp 1667941163
transform -1 0 27416 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1084_
timestamp 1667941163
transform 1 0 22172 0 1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1084__81
timestamp 1667941163
transform -1 0 22724 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1085__82
timestamp 1667941163
transform -1 0 19688 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1085_
timestamp 1667941163
transform 1 0 19228 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1086__83
timestamp 1667941163
transform 1 0 27784 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1086_
timestamp 1667941163
transform -1 0 28428 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1087__84
timestamp 1667941163
transform -1 0 2024 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1087_
timestamp 1667941163
transform 1 0 1656 0 -1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1088_
timestamp 1667941163
transform 1 0 26496 0 1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1088__85
timestamp 1667941163
transform -1 0 28152 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1089__86
timestamp 1667941163
transform 1 0 2024 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1089_
timestamp 1667941163
transform -1 0 3496 0 1 43520
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1090__87
timestamp 1667941163
transform -1 0 4232 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1090_
timestamp 1667941163
transform 1 0 3956 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1091_
timestamp 1667941163
transform 1 0 7728 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1091__88
timestamp 1667941163
transform -1 0 8096 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1092__89
timestamp 1667941163
transform -1 0 3680 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1092_
timestamp 1667941163
transform -1 0 3496 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1093__90
timestamp 1667941163
transform 1 0 27876 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1093_
timestamp 1667941163
transform -1 0 28428 0 1 30464
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1094__91
timestamp 1667941163
transform 1 0 27692 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1094_
timestamp 1667941163
transform -1 0 28428 0 1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1095_
timestamp 1667941163
transform -1 0 28428 0 1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1095__92
timestamp 1667941163
transform 1 0 27416 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1096__93
timestamp 1667941163
transform -1 0 5428 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1096_
timestamp 1667941163
transform -1 0 3496 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1097__94
timestamp 1667941163
transform -1 0 4876 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1097_
timestamp 1667941163
transform -1 0 3864 0 -1 43520
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1098__95
timestamp 1667941163
transform -1 0 28152 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1098_
timestamp 1667941163
transform 1 0 26496 0 1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1099__96
timestamp 1667941163
transform 1 0 11224 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1099_
timestamp 1667941163
transform 1 0 11684 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1100__97
timestamp 1667941163
transform 1 0 18308 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1100_
timestamp 1667941163
transform 1 0 19136 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1101_
timestamp 1667941163
transform -1 0 3496 0 1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1101__98
timestamp 1667941163
transform 1 0 3128 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1102__99
timestamp 1667941163
transform 1 0 27968 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1102_
timestamp 1667941163
transform -1 0 28428 0 1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1103__100
timestamp 1667941163
transform -1 0 2024 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1103_
timestamp 1667941163
transform 1 0 1656 0 -1 41344
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1104_
timestamp 1667941163
transform 1 0 3680 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1104__101
timestamp 1667941163
transform 1 0 3036 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1105_
timestamp 1667941163
transform 1 0 9292 0 1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1105__102
timestamp 1667941163
transform -1 0 9936 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1106_
timestamp 1667941163
transform 1 0 9292 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1106__103
timestamp 1667941163
transform -1 0 10580 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1107__104
timestamp 1667941163
transform 1 0 26404 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1107_
timestamp 1667941163
transform -1 0 26680 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1108__105
timestamp 1667941163
transform 1 0 27876 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1108_
timestamp 1667941163
transform -1 0 28428 0 1 42432
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1109__106
timestamp 1667941163
transform 1 0 12972 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1109_
timestamp 1667941163
transform -1 0 13984 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1110__107
timestamp 1667941163
transform -1 0 28152 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1110_
timestamp 1667941163
transform -1 0 26680 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1111_
timestamp 1667941163
transform -1 0 28428 0 1 36992
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1111__108
timestamp 1667941163
transform 1 0 28060 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1112__109
timestamp 1667941163
transform 1 0 1748 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1112_
timestamp 1667941163
transform -1 0 3496 0 1 41344
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1113__110
timestamp 1667941163
transform -1 0 28060 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1113_
timestamp 1667941163
transform -1 0 26680 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1114__111
timestamp 1667941163
transform -1 0 1932 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1114_
timestamp 1667941163
transform 1 0 1564 0 1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1115_
timestamp 1667941163
transform 1 0 26496 0 1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1115__112
timestamp 1667941163
transform -1 0 28060 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1116__113
timestamp 1667941163
transform -1 0 1932 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1116_
timestamp 1667941163
transform 1 0 1564 0 1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1117_
timestamp 1667941163
transform 1 0 1564 0 1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1117__114
timestamp 1667941163
transform -1 0 1932 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1118__115
timestamp 1667941163
transform -1 0 1932 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1118_
timestamp 1667941163
transform 1 0 1656 0 -1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1119_
timestamp 1667941163
transform -1 0 3496 0 1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1119__116
timestamp 1667941163
transform 1 0 2116 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_wb_clk_i $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 24012 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_0__f_wb_clk_i
timestamp 1667941163
transform -1 0 20056 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_1__f_wb_clk_i
timestamp 1667941163
transform -1 0 22632 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_2__f_wb_clk_i
timestamp 1667941163
transform -1 0 20056 0 -1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_3__f_wb_clk_i
timestamp 1667941163
transform -1 0 22632 0 1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 24656 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 1667941163
transform -1 0 27876 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1667941163
transform 1 0 1564 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1667941163
transform 1 0 27140 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1667941163
transform 1 0 28152 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1667941163
transform 1 0 18032 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1667941163
transform -1 0 25760 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1667941163
transform -1 0 1840 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1667941163
transform 1 0 27140 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input8 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 16008 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input9 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 9108 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1667941163
transform -1 0 1840 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1667941163
transform 1 0 24564 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1667941163
transform 1 0 26404 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1667941163
transform -1 0 6072 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1667941163
transform -1 0 1840 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input15
timestamp 1667941163
transform -1 0 6808 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input16
timestamp 1667941163
transform -1 0 1840 0 -1 28288
box -38 -48 314 592
<< labels >>
flabel metal3 s 200 36668 800 36908 0 FreeSans 960 0 0 0 active
port 0 nsew signal input
flabel metal2 s 12226 200 12338 800 0 FreeSans 448 90 0 0 io_in[0]
port 1 nsew signal input
flabel metal2 s 12226 49200 12338 49800 0 FreeSans 448 90 0 0 io_in[10]
port 2 nsew signal input
flabel metal3 s 200 40068 800 40308 0 FreeSans 960 0 0 0 io_in[11]
port 3 nsew signal input
flabel metal3 s 29200 43468 29800 43708 0 FreeSans 960 0 0 0 io_in[12]
port 4 nsew signal input
flabel metal2 s 18666 200 18778 800 0 FreeSans 448 90 0 0 io_in[13]
port 5 nsew signal input
flabel metal2 s 5142 49200 5254 49800 0 FreeSans 448 90 0 0 io_in[14]
port 6 nsew signal input
flabel metal3 s 29200 45508 29800 45748 0 FreeSans 960 0 0 0 io_in[15]
port 7 nsew signal input
flabel metal3 s 29200 13548 29800 13788 0 FreeSans 960 0 0 0 io_in[16]
port 8 nsew signal input
flabel metal3 s 200 48228 800 48468 0 FreeSans 960 0 0 0 io_in[17]
port 9 nsew signal input
flabel metal2 s -10 49200 102 49800 0 FreeSans 448 90 0 0 io_in[18]
port 10 nsew signal input
flabel metal3 s 29200 4028 29800 4268 0 FreeSans 960 0 0 0 io_in[19]
port 11 nsew signal input
flabel metal3 s 200 12868 800 13108 0 FreeSans 960 0 0 0 io_in[1]
port 12 nsew signal input
flabel metal3 s 200 23068 800 23308 0 FreeSans 960 0 0 0 io_in[20]
port 13 nsew signal input
flabel metal3 s 200 14908 800 15148 0 FreeSans 960 0 0 0 io_in[21]
port 14 nsew signal input
flabel metal3 s 29200 23068 29800 23308 0 FreeSans 960 0 0 0 io_in[22]
port 15 nsew signal input
flabel metal3 s 200 47548 800 47788 0 FreeSans 960 0 0 0 io_in[23]
port 16 nsew signal input
flabel metal3 s 200 45508 800 45748 0 FreeSans 960 0 0 0 io_in[24]
port 17 nsew signal input
flabel metal2 s 29614 200 29726 800 0 FreeSans 448 90 0 0 io_in[25]
port 18 nsew signal input
flabel metal2 s 28970 200 29082 800 0 FreeSans 448 90 0 0 io_in[26]
port 19 nsew signal input
flabel metal3 s 29200 18988 29800 19228 0 FreeSans 960 0 0 0 io_in[27]
port 20 nsew signal input
flabel metal2 s 26394 200 26506 800 0 FreeSans 448 90 0 0 io_in[28]
port 21 nsew signal input
flabel metal2 s 29614 49200 29726 49800 0 FreeSans 448 90 0 0 io_in[29]
port 22 nsew signal input
flabel metal2 s 12870 200 12982 800 0 FreeSans 448 90 0 0 io_in[2]
port 23 nsew signal input
flabel metal3 s 29200 25788 29800 26028 0 FreeSans 960 0 0 0 io_in[30]
port 24 nsew signal input
flabel metal3 s 200 35308 800 35548 0 FreeSans 960 0 0 0 io_in[31]
port 25 nsew signal input
flabel metal2 s 24462 200 24574 800 0 FreeSans 448 90 0 0 io_in[32]
port 26 nsew signal input
flabel metal3 s 200 20348 800 20588 0 FreeSans 960 0 0 0 io_in[33]
port 27 nsew signal input
flabel metal2 s 20598 49200 20710 49800 0 FreeSans 448 90 0 0 io_in[34]
port 28 nsew signal input
flabel metal2 s 25106 49200 25218 49800 0 FreeSans 448 90 0 0 io_in[35]
port 29 nsew signal input
flabel metal3 s 29200 35308 29800 35548 0 FreeSans 960 0 0 0 io_in[36]
port 30 nsew signal input
flabel metal2 s 25750 49200 25862 49800 0 FreeSans 448 90 0 0 io_in[37]
port 31 nsew signal input
flabel metal2 s 12870 49200 12982 49800 0 FreeSans 448 90 0 0 io_in[3]
port 32 nsew signal input
flabel metal3 s 29200 34628 29800 34868 0 FreeSans 960 0 0 0 io_in[4]
port 33 nsew signal input
flabel metal3 s 29200 48228 29800 48468 0 FreeSans 960 0 0 0 io_in[5]
port 34 nsew signal input
flabel metal3 s 200 24428 800 24668 0 FreeSans 960 0 0 0 io_in[6]
port 35 nsew signal input
flabel metal3 s 200 16948 800 17188 0 FreeSans 960 0 0 0 io_in[7]
port 36 nsew signal input
flabel metal3 s 29200 36668 29800 36908 0 FreeSans 960 0 0 0 io_in[8]
port 37 nsew signal input
flabel metal3 s 200 46868 800 47108 0 FreeSans 960 0 0 0 io_in[9]
port 38 nsew signal input
flabel metal2 s 21242 200 21354 800 0 FreeSans 448 90 0 0 io_oeb[0]
port 39 nsew signal tristate
flabel metal3 s 200 13548 800 13788 0 FreeSans 960 0 0 0 io_oeb[10]
port 40 nsew signal tristate
flabel metal3 s 29200 32588 29800 32828 0 FreeSans 960 0 0 0 io_oeb[11]
port 41 nsew signal tristate
flabel metal3 s 29200 21708 29800 21948 0 FreeSans 960 0 0 0 io_oeb[12]
port 42 nsew signal tristate
flabel metal3 s 29200 21028 29800 21268 0 FreeSans 960 0 0 0 io_oeb[13]
port 43 nsew signal tristate
flabel metal3 s 200 3348 800 3588 0 FreeSans 960 0 0 0 io_oeb[14]
port 44 nsew signal tristate
flabel metal2 s 1278 49200 1390 49800 0 FreeSans 448 90 0 0 io_oeb[15]
port 45 nsew signal tristate
flabel metal3 s 29200 12188 29800 12428 0 FreeSans 960 0 0 0 io_oeb[16]
port 46 nsew signal tristate
flabel metal2 s 10938 200 11050 800 0 FreeSans 448 90 0 0 io_oeb[17]
port 47 nsew signal tristate
flabel metal2 s 18666 49200 18778 49800 0 FreeSans 448 90 0 0 io_oeb[18]
port 48 nsew signal tristate
flabel metal2 s 1922 49200 2034 49800 0 FreeSans 448 90 0 0 io_oeb[19]
port 49 nsew signal tristate
flabel metal3 s 29200 1308 29800 1548 0 FreeSans 960 0 0 0 io_oeb[1]
port 50 nsew signal tristate
flabel metal3 s 29200 27148 29800 27388 0 FreeSans 960 0 0 0 io_oeb[20]
port 51 nsew signal tristate
flabel metal3 s 200 41428 800 41668 0 FreeSans 960 0 0 0 io_oeb[21]
port 52 nsew signal tristate
flabel metal2 s 3854 200 3966 800 0 FreeSans 448 90 0 0 io_oeb[22]
port 53 nsew signal tristate
flabel metal2 s 10294 49200 10406 49800 0 FreeSans 448 90 0 0 io_oeb[23]
port 54 nsew signal tristate
flabel metal2 s 10938 49200 11050 49800 0 FreeSans 448 90 0 0 io_oeb[24]
port 55 nsew signal tristate
flabel metal3 s 29200 8108 29800 8348 0 FreeSans 960 0 0 0 io_oeb[25]
port 56 nsew signal tristate
flabel metal3 s 29200 41428 29800 41668 0 FreeSans 960 0 0 0 io_oeb[26]
port 57 nsew signal tristate
flabel metal2 s 13514 49200 13626 49800 0 FreeSans 448 90 0 0 io_oeb[27]
port 58 nsew signal tristate
flabel metal3 s 29200 3348 29800 3588 0 FreeSans 960 0 0 0 io_oeb[28]
port 59 nsew signal tristate
flabel metal3 s 29200 35988 29800 36228 0 FreeSans 960 0 0 0 io_oeb[29]
port 60 nsew signal tristate
flabel metal2 s 23174 49200 23286 49800 0 FreeSans 448 90 0 0 io_oeb[2]
port 61 nsew signal tristate
flabel metal3 s 200 42108 800 42348 0 FreeSans 960 0 0 0 io_oeb[30]
port 62 nsew signal tristate
flabel metal3 s 29200 2668 29800 2908 0 FreeSans 960 0 0 0 io_oeb[31]
port 63 nsew signal tristate
flabel metal3 s 200 19668 800 19908 0 FreeSans 960 0 0 0 io_oeb[32]
port 64 nsew signal tristate
flabel metal3 s 29200 8788 29800 9028 0 FreeSans 960 0 0 0 io_oeb[33]
port 65 nsew signal tristate
flabel metal3 s 200 49588 800 49828 0 FreeSans 960 0 0 0 io_oeb[34]
port 66 nsew signal tristate
flabel metal3 s 200 17628 800 17868 0 FreeSans 960 0 0 0 io_oeb[35]
port 67 nsew signal tristate
flabel metal3 s 200 8788 800 9028 0 FreeSans 960 0 0 0 io_oeb[36]
port 68 nsew signal tristate
flabel metal3 s 200 14228 800 14468 0 FreeSans 960 0 0 0 io_oeb[37]
port 69 nsew signal tristate
flabel metal2 s 19954 200 20066 800 0 FreeSans 448 90 0 0 io_oeb[3]
port 70 nsew signal tristate
flabel metal3 s 29200 10148 29800 10388 0 FreeSans 960 0 0 0 io_oeb[4]
port 71 nsew signal tristate
flabel metal3 s 200 25788 800 26028 0 FreeSans 960 0 0 0 io_oeb[5]
port 72 nsew signal tristate
flabel metal3 s 29200 24428 29800 24668 0 FreeSans 960 0 0 0 io_oeb[6]
port 73 nsew signal tristate
flabel metal2 s 634 49200 746 49800 0 FreeSans 448 90 0 0 io_oeb[7]
port 74 nsew signal tristate
flabel metal2 s 3210 200 3322 800 0 FreeSans 448 90 0 0 io_oeb[8]
port 75 nsew signal tristate
flabel metal2 s 8362 200 8474 800 0 FreeSans 448 90 0 0 io_oeb[9]
port 76 nsew signal tristate
flabel metal3 s 29200 47548 29800 47788 0 FreeSans 960 0 0 0 io_out[0]
port 77 nsew signal tristate
flabel metal3 s 29200 31908 29800 32148 0 FreeSans 960 0 0 0 io_out[10]
port 78 nsew signal tristate
flabel metal3 s 200 1988 800 2228 0 FreeSans 960 0 0 0 io_out[11]
port 79 nsew signal tristate
flabel metal3 s 200 6068 800 6308 0 FreeSans 960 0 0 0 io_out[12]
port 80 nsew signal tristate
flabel metal3 s 29200 1988 29800 2228 0 FreeSans 960 0 0 0 io_out[13]
port 81 nsew signal tristate
flabel metal3 s 29200 42108 29800 42348 0 FreeSans 960 0 0 0 io_out[14]
port 82 nsew signal tristate
flabel metal3 s 200 33268 800 33508 0 FreeSans 960 0 0 0 io_out[15]
port 83 nsew signal tristate
flabel metal3 s 29200 31228 29800 31468 0 FreeSans 960 0 0 0 io_out[16]
port 84 nsew signal tristate
flabel metal2 s 27038 49200 27150 49800 0 FreeSans 448 90 0 0 io_out[17]
port 85 nsew signal tristate
flabel metal3 s 29200 7428 29800 7668 0 FreeSans 960 0 0 0 io_out[18]
port 86 nsew signal tristate
flabel metal3 s 200 18988 800 19228 0 FreeSans 960 0 0 0 io_out[19]
port 87 nsew signal tristate
flabel metal2 s 16734 49200 16846 49800 0 FreeSans 448 90 0 0 io_out[1]
port 88 nsew signal tristate
flabel metal2 s 22530 49200 22642 49800 0 FreeSans 448 90 0 0 io_out[20]
port 89 nsew signal tristate
flabel metal3 s 200 31908 800 32148 0 FreeSans 960 0 0 0 io_out[21]
port 90 nsew signal tristate
flabel metal2 s 25106 200 25218 800 0 FreeSans 448 90 0 0 io_out[22]
port 91 nsew signal tristate
flabel metal3 s 29200 28508 29800 28748 0 FreeSans 960 0 0 0 io_out[23]
port 92 nsew signal tristate
flabel metal2 s 21886 200 21998 800 0 FreeSans 448 90 0 0 io_out[24]
port 93 nsew signal tristate
flabel metal2 s 19954 49200 20066 49800 0 FreeSans 448 90 0 0 io_out[25]
port 94 nsew signal tristate
flabel metal3 s 200 4028 800 4268 0 FreeSans 960 0 0 0 io_out[26]
port 95 nsew signal tristate
flabel metal2 s 21242 49200 21354 49800 0 FreeSans 448 90 0 0 io_out[27]
port 96 nsew signal tristate
flabel metal2 s 13514 200 13626 800 0 FreeSans 448 90 0 0 io_out[28]
port 97 nsew signal tristate
flabel metal3 s 29200 10828 29800 11068 0 FreeSans 960 0 0 0 io_out[29]
port 98 nsew signal tristate
flabel metal2 s 5786 200 5898 800 0 FreeSans 448 90 0 0 io_out[2]
port 99 nsew signal tristate
flabel metal3 s 200 4708 800 4948 0 FreeSans 960 0 0 0 io_out[30]
port 100 nsew signal tristate
flabel metal3 s 200 11508 800 11748 0 FreeSans 960 0 0 0 io_out[31]
port 101 nsew signal tristate
flabel metal3 s 200 37348 800 37588 0 FreeSans 960 0 0 0 io_out[32]
port 102 nsew signal tristate
flabel metal3 s 29200 15588 29800 15828 0 FreeSans 960 0 0 0 io_out[33]
port 103 nsew signal tristate
flabel metal3 s 29200 42788 29800 43028 0 FreeSans 960 0 0 0 io_out[34]
port 104 nsew signal tristate
flabel metal3 s 29200 40748 29800 40988 0 FreeSans 960 0 0 0 io_out[35]
port 105 nsew signal tristate
flabel metal2 s 2566 49200 2678 49800 0 FreeSans 448 90 0 0 io_out[36]
port 106 nsew signal tristate
flabel metal3 s 29200 46188 29800 46428 0 FreeSans 960 0 0 0 io_out[37]
port 107 nsew signal tristate
flabel metal3 s 200 34628 800 34868 0 FreeSans 960 0 0 0 io_out[3]
port 108 nsew signal tristate
flabel metal3 s 29200 33948 29800 34188 0 FreeSans 960 0 0 0 io_out[4]
port 109 nsew signal tristate
flabel metal2 s 8362 49200 8474 49800 0 FreeSans 448 90 0 0 io_out[5]
port 110 nsew signal tristate
flabel metal2 s 28326 49200 28438 49800 0 FreeSans 448 90 0 0 io_out[6]
port 111 nsew signal tristate
flabel metal3 s 200 15588 800 15828 0 FreeSans 960 0 0 0 io_out[7]
port 112 nsew signal tristate
flabel metal2 s 14802 200 14914 800 0 FreeSans 448 90 0 0 io_out[8]
port 113 nsew signal tristate
flabel metal3 s 200 12188 800 12428 0 FreeSans 960 0 0 0 io_out[9]
port 114 nsew signal tristate
flabel metal3 s 29200 16268 29800 16508 0 FreeSans 960 0 0 0 la1_data_in[0]
port 115 nsew signal input
flabel metal2 s 17378 200 17490 800 0 FreeSans 448 90 0 0 la1_data_in[10]
port 116 nsew signal input
flabel metal3 s 29200 14908 29800 15148 0 FreeSans 960 0 0 0 la1_data_in[11]
port 117 nsew signal input
flabel metal3 s 200 29868 800 30108 0 FreeSans 960 0 0 0 la1_data_in[12]
port 118 nsew signal input
flabel metal2 s 27038 200 27150 800 0 FreeSans 448 90 0 0 la1_data_in[13]
port 119 nsew signal input
flabel metal3 s 200 10148 800 10388 0 FreeSans 960 0 0 0 la1_data_in[14]
port 120 nsew signal input
flabel metal2 s 3210 49200 3322 49800 0 FreeSans 448 90 0 0 la1_data_in[15]
port 121 nsew signal input
flabel metal2 s 15446 49200 15558 49800 0 FreeSans 448 90 0 0 la1_data_in[16]
port 122 nsew signal input
flabel metal2 s 9650 49200 9762 49800 0 FreeSans 448 90 0 0 la1_data_in[17]
port 123 nsew signal input
flabel metal3 s 29200 4708 29800 4948 0 FreeSans 960 0 0 0 la1_data_in[18]
port 124 nsew signal input
flabel metal2 s 4498 49200 4610 49800 0 FreeSans 448 90 0 0 la1_data_in[19]
port 125 nsew signal input
flabel metal2 s 16090 200 16202 800 0 FreeSans 448 90 0 0 la1_data_in[1]
port 126 nsew signal input
flabel metal3 s 200 29188 800 29428 0 FreeSans 960 0 0 0 la1_data_in[20]
port 127 nsew signal input
flabel metal2 s 28970 49200 29082 49800 0 FreeSans 448 90 0 0 la1_data_in[21]
port 128 nsew signal input
flabel metal3 s 29200 17628 29800 17868 0 FreeSans 960 0 0 0 la1_data_in[22]
port 129 nsew signal input
flabel metal3 s 200 628 800 868 0 FreeSans 960 0 0 0 la1_data_in[23]
port 130 nsew signal input
flabel metal2 s 11582 200 11694 800 0 FreeSans 448 90 0 0 la1_data_in[24]
port 131 nsew signal input
flabel metal3 s 200 30548 800 30788 0 FreeSans 960 0 0 0 la1_data_in[25]
port 132 nsew signal input
flabel metal3 s 29200 12868 29800 13108 0 FreeSans 960 0 0 0 la1_data_in[26]
port 133 nsew signal input
flabel metal2 s 23174 200 23286 800 0 FreeSans 448 90 0 0 la1_data_in[27]
port 134 nsew signal input
flabel metal3 s 200 26468 800 26708 0 FreeSans 960 0 0 0 la1_data_in[28]
port 135 nsew signal input
flabel metal3 s 200 40748 800 40988 0 FreeSans 960 0 0 0 la1_data_in[29]
port 136 nsew signal input
flabel metal2 s 9006 200 9118 800 0 FreeSans 448 90 0 0 la1_data_in[2]
port 137 nsew signal input
flabel metal2 s 1278 200 1390 800 0 FreeSans 448 90 0 0 la1_data_in[30]
port 138 nsew signal input
flabel metal3 s 29200 -52 29800 188 0 FreeSans 960 0 0 0 la1_data_in[31]
port 139 nsew signal input
flabel metal3 s 200 25108 800 25348 0 FreeSans 960 0 0 0 la1_data_in[3]
port 140 nsew signal input
flabel metal2 s 23818 49200 23930 49800 0 FreeSans 448 90 0 0 la1_data_in[4]
port 141 nsew signal input
flabel metal3 s 29200 29868 29800 30108 0 FreeSans 960 0 0 0 la1_data_in[5]
port 142 nsew signal input
flabel metal2 s 5786 49200 5898 49800 0 FreeSans 448 90 0 0 la1_data_in[6]
port 143 nsew signal input
flabel metal3 s 200 18308 800 18548 0 FreeSans 960 0 0 0 la1_data_in[7]
port 144 nsew signal input
flabel metal2 s 6430 49200 6542 49800 0 FreeSans 448 90 0 0 la1_data_in[8]
port 145 nsew signal input
flabel metal3 s 200 27828 800 28068 0 FreeSans 960 0 0 0 la1_data_in[9]
port 146 nsew signal input
flabel metal2 s 6430 200 6542 800 0 FreeSans 448 90 0 0 la1_data_out[0]
port 147 nsew signal tristate
flabel metal3 s 29200 19668 29800 19908 0 FreeSans 960 0 0 0 la1_data_out[10]
port 148 nsew signal tristate
flabel metal2 s 18022 200 18134 800 0 FreeSans 448 90 0 0 la1_data_out[11]
port 149 nsew signal tristate
flabel metal3 s 29200 46868 29800 47108 0 FreeSans 960 0 0 0 la1_data_out[12]
port 150 nsew signal tristate
flabel metal3 s 200 44148 800 44388 0 FreeSans 960 0 0 0 la1_data_out[13]
port 151 nsew signal tristate
flabel metal2 s 11582 49200 11694 49800 0 FreeSans 448 90 0 0 la1_data_out[14]
port 152 nsew signal tristate
flabel metal3 s 200 1308 800 1548 0 FreeSans 960 0 0 0 la1_data_out[15]
port 153 nsew signal tristate
flabel metal3 s 29200 23748 29800 23988 0 FreeSans 960 0 0 0 la1_data_out[16]
port 154 nsew signal tristate
flabel metal3 s 29200 39388 29800 39628 0 FreeSans 960 0 0 0 la1_data_out[17]
port 155 nsew signal tristate
flabel metal3 s 200 44828 800 45068 0 FreeSans 960 0 0 0 la1_data_out[18]
port 156 nsew signal tristate
flabel metal3 s 29200 30548 29800 30788 0 FreeSans 960 0 0 0 la1_data_out[19]
port 157 nsew signal tristate
flabel metal3 s 200 35988 800 36228 0 FreeSans 960 0 0 0 la1_data_out[1]
port 158 nsew signal tristate
flabel metal3 s 200 8108 800 8348 0 FreeSans 960 0 0 0 la1_data_out[20]
port 159 nsew signal tristate
flabel metal3 s 29200 44828 29800 45068 0 FreeSans 960 0 0 0 la1_data_out[21]
port 160 nsew signal tristate
flabel metal2 s 14802 49200 14914 49800 0 FreeSans 448 90 0 0 la1_data_out[22]
port 161 nsew signal tristate
flabel metal2 s 9650 200 9762 800 0 FreeSans 448 90 0 0 la1_data_out[23]
port 162 nsew signal tristate
flabel metal3 s 29200 25108 29800 25348 0 FreeSans 960 0 0 0 la1_data_out[24]
port 163 nsew signal tristate
flabel metal3 s 200 2668 800 2908 0 FreeSans 960 0 0 0 la1_data_out[25]
port 164 nsew signal tristate
flabel metal3 s 29200 14228 29800 14468 0 FreeSans 960 0 0 0 la1_data_out[26]
port 165 nsew signal tristate
flabel metal3 s 200 38708 800 38948 0 FreeSans 960 0 0 0 la1_data_out[27]
port 166 nsew signal tristate
flabel metal3 s 29200 5388 29800 5628 0 FreeSans 960 0 0 0 la1_data_out[28]
port 167 nsew signal tristate
flabel metal2 s 4498 200 4610 800 0 FreeSans 448 90 0 0 la1_data_out[29]
port 168 nsew signal tristate
flabel metal2 s 16734 200 16846 800 0 FreeSans 448 90 0 0 la1_data_out[2]
port 169 nsew signal tristate
flabel metal3 s 29200 20348 29800 20588 0 FreeSans 960 0 0 0 la1_data_out[30]
port 170 nsew signal tristate
flabel metal3 s 29200 48908 29800 49148 0 FreeSans 960 0 0 0 la1_data_out[31]
port 171 nsew signal tristate
flabel metal3 s 200 7428 800 7668 0 FreeSans 960 0 0 0 la1_data_out[3]
port 172 nsew signal tristate
flabel metal3 s 29200 6748 29800 6988 0 FreeSans 960 0 0 0 la1_data_out[4]
port 173 nsew signal tristate
flabel metal2 s 2566 200 2678 800 0 FreeSans 448 90 0 0 la1_data_out[5]
port 174 nsew signal tristate
flabel metal3 s 29200 26468 29800 26708 0 FreeSans 960 0 0 0 la1_data_out[6]
port 175 nsew signal tristate
flabel metal2 s 634 200 746 800 0 FreeSans 448 90 0 0 la1_data_out[7]
port 176 nsew signal tristate
flabel metal3 s 29200 40068 29800 40308 0 FreeSans 960 0 0 0 la1_data_out[8]
port 177 nsew signal tristate
flabel metal2 s 27682 49200 27794 49800 0 FreeSans 448 90 0 0 la1_data_out[9]
port 178 nsew signal tristate
flabel metal3 s 29200 9468 29800 9708 0 FreeSans 960 0 0 0 la1_oenb[0]
port 179 nsew signal input
flabel metal2 s 26394 49200 26506 49800 0 FreeSans 448 90 0 0 la1_oenb[10]
port 180 nsew signal input
flabel metal3 s 200 22388 800 22628 0 FreeSans 960 0 0 0 la1_oenb[11]
port 181 nsew signal input
flabel metal3 s 200 23748 800 23988 0 FreeSans 960 0 0 0 la1_oenb[12]
port 182 nsew signal input
flabel metal2 s 23818 200 23930 800 0 FreeSans 448 90 0 0 la1_oenb[13]
port 183 nsew signal input
flabel metal2 s -10 200 102 800 0 FreeSans 448 90 0 0 la1_oenb[14]
port 184 nsew signal input
flabel metal2 s 28326 200 28438 800 0 FreeSans 448 90 0 0 la1_oenb[15]
port 185 nsew signal input
flabel metal3 s 200 28508 800 28748 0 FreeSans 960 0 0 0 la1_oenb[16]
port 186 nsew signal input
flabel metal3 s 200 42788 800 43028 0 FreeSans 960 0 0 0 la1_oenb[17]
port 187 nsew signal input
flabel metal2 s 7718 49200 7830 49800 0 FreeSans 448 90 0 0 la1_oenb[18]
port 188 nsew signal input
flabel metal3 s 200 21028 800 21268 0 FreeSans 960 0 0 0 la1_oenb[19]
port 189 nsew signal input
flabel metal2 s 7074 200 7186 800 0 FreeSans 448 90 0 0 la1_oenb[1]
port 190 nsew signal input
flabel metal2 s 1922 200 2034 800 0 FreeSans 448 90 0 0 la1_oenb[20]
port 191 nsew signal input
flabel metal2 s 16090 49200 16202 49800 0 FreeSans 448 90 0 0 la1_oenb[21]
port 192 nsew signal input
flabel metal2 s 7074 49200 7186 49800 0 FreeSans 448 90 0 0 la1_oenb[22]
port 193 nsew signal input
flabel metal2 s 19310 200 19422 800 0 FreeSans 448 90 0 0 la1_oenb[23]
port 194 nsew signal input
flabel metal2 s 21886 49200 21998 49800 0 FreeSans 448 90 0 0 la1_oenb[24]
port 195 nsew signal input
flabel metal3 s 29200 18308 29800 18548 0 FreeSans 960 0 0 0 la1_oenb[25]
port 196 nsew signal input
flabel metal3 s 200 31228 800 31468 0 FreeSans 960 0 0 0 la1_oenb[26]
port 197 nsew signal input
flabel metal3 s 29200 38028 29800 38268 0 FreeSans 960 0 0 0 la1_oenb[27]
port 198 nsew signal input
flabel metal2 s 7718 200 7830 800 0 FreeSans 448 90 0 0 la1_oenb[28]
port 199 nsew signal input
flabel metal2 s 14158 200 14270 800 0 FreeSans 448 90 0 0 la1_oenb[29]
port 200 nsew signal input
flabel metal3 s 200 6748 800 6988 0 FreeSans 960 0 0 0 la1_oenb[2]
port 201 nsew signal input
flabel metal3 s 29200 37348 29800 37588 0 FreeSans 960 0 0 0 la1_oenb[30]
port 202 nsew signal input
flabel metal2 s 22530 200 22642 800 0 FreeSans 448 90 0 0 la1_oenb[31]
port 203 nsew signal input
flabel metal2 s 18022 49200 18134 49800 0 FreeSans 448 90 0 0 la1_oenb[3]
port 204 nsew signal input
flabel metal2 s 17378 49200 17490 49800 0 FreeSans 448 90 0 0 la1_oenb[4]
port 205 nsew signal input
flabel metal3 s 200 39388 800 39628 0 FreeSans 960 0 0 0 la1_oenb[5]
port 206 nsew signal input
flabel metal3 s 200 46188 800 46428 0 FreeSans 960 0 0 0 la1_oenb[6]
port 207 nsew signal input
flabel metal2 s 27682 200 27794 800 0 FreeSans 448 90 0 0 la1_oenb[7]
port 208 nsew signal input
flabel metal3 s 200 9468 800 9708 0 FreeSans 960 0 0 0 la1_oenb[8]
port 209 nsew signal input
flabel metal3 s 200 33948 800 34188 0 FreeSans 960 0 0 0 la1_oenb[9]
port 210 nsew signal input
flabel metal4 s 4417 2128 4737 47376 0 FreeSans 1920 90 0 0 vccd1
port 211 nsew power bidirectional
flabel metal4 s 11363 2128 11683 47376 0 FreeSans 1920 90 0 0 vccd1
port 211 nsew power bidirectional
flabel metal4 s 18309 2128 18629 47376 0 FreeSans 1920 90 0 0 vccd1
port 211 nsew power bidirectional
flabel metal4 s 25255 2128 25575 47376 0 FreeSans 1920 90 0 0 vccd1
port 211 nsew power bidirectional
flabel metal4 s 7890 2128 8210 47376 0 FreeSans 1920 90 0 0 vssd1
port 212 nsew ground bidirectional
flabel metal4 s 14836 2128 15156 47376 0 FreeSans 1920 90 0 0 vssd1
port 212 nsew ground bidirectional
flabel metal4 s 21782 2128 22102 47376 0 FreeSans 1920 90 0 0 vssd1
port 212 nsew ground bidirectional
flabel metal4 s 28728 2128 29048 47376 0 FreeSans 1920 90 0 0 vssd1
port 212 nsew ground bidirectional
flabel metal3 s 29200 29188 29800 29428 0 FreeSans 960 0 0 0 wb_clk_i
port 213 nsew signal input
rlabel metal1 14996 47328 14996 47328 0 vccd1
rlabel via1 15076 46784 15076 46784 0 vssd1
rlabel metal1 22489 32402 22489 32402 0 _0000_
rlabel metal2 22218 33762 22218 33762 0 _0001_
rlabel metal2 21758 26554 21758 26554 0 _0002_
rlabel metal1 25571 18326 25571 18326 0 _0003_
rlabel via1 26077 19822 26077 19822 0 _0004_
rlabel metal1 25709 22678 25709 22678 0 _0005_
rlabel metal2 26082 31110 26082 31110 0 _0006_
rlabel metal2 26174 28322 26174 28322 0 _0007_
rlabel metal1 22673 29138 22673 29138 0 _0008_
rlabel metal1 20700 16218 20700 16218 0 _0009_
rlabel via1 18349 17238 18349 17238 0 _0010_
rlabel metal1 20332 14042 20332 14042 0 _0011_
rlabel metal1 19688 14586 19688 14586 0 _0012_
rlabel via1 21109 18734 21109 18734 0 _0013_
rlabel metal2 18906 25670 18906 25670 0 _0014_
rlabel metal1 18579 23766 18579 23766 0 _0015_
rlabel metal1 18952 20570 18952 20570 0 _0016_
rlabel metal1 16964 24174 16964 24174 0 _0017_
rlabel metal2 17158 25670 17158 25670 0 _0018_
rlabel metal1 22586 36006 22586 36006 0 _0019_
rlabel metal1 23087 32878 23087 32878 0 _0020_
rlabel metal1 17383 34986 17383 34986 0 _0021_
rlabel metal1 16882 21862 16882 21862 0 _0022_
rlabel via1 17153 35734 17153 35734 0 _0023_
rlabel metal2 17066 27234 17066 27234 0 _0024_
rlabel via1 17153 16082 17153 16082 0 _0025_
rlabel metal1 26813 15470 26813 15470 0 _0026_
rlabel metal1 16866 22678 16866 22678 0 _0027_
rlabel metal2 25806 14178 25806 14178 0 _0028_
rlabel metal2 20838 29852 20838 29852 0 _0029_
rlabel metal1 22259 20910 22259 20910 0 _0030_
rlabel metal2 20838 26418 20838 26418 0 _0031_
rlabel metal1 21114 23290 21114 23290 0 _0032_
rlabel via1 20842 20910 20842 20910 0 _0033_
rlabel via1 24421 17170 24421 17170 0 _0034_
rlabel metal1 24016 15062 24016 15062 0 _0035_
rlabel metal1 21742 15402 21742 15402 0 _0036_
rlabel metal1 24978 14042 24978 14042 0 _0037_
rlabel metal1 19632 28526 19632 28526 0 _0038_
rlabel via1 20373 36142 20373 36142 0 _0039_
rlabel metal1 22310 37638 22310 37638 0 _0040_
rlabel metal1 19458 38794 19458 38794 0 _0041_
rlabel metal1 18722 36550 18722 36550 0 _0042_
rlabel metal1 17148 31790 17148 31790 0 _0043_
rlabel metal1 17056 30226 17056 30226 0 _0044_
rlabel metal1 16964 28526 16964 28526 0 _0045_
rlabel via1 16969 18734 16969 18734 0 _0046_
rlabel via1 17245 19414 17245 19414 0 _0047_
rlabel metal1 17940 14586 17940 14586 0 _0048_
rlabel metal1 17250 14042 17250 14042 0 _0049_
rlabel metal2 22862 23970 22862 23970 0 _0050_
rlabel metal2 24794 35462 24794 35462 0 _0051_
rlabel metal2 2622 36448 2622 36448 0 _0052_
rlabel metal2 3266 37740 3266 37740 0 _0053_
rlabel metal2 2530 18802 2530 18802 0 _0054_
rlabel metal1 2530 45424 2530 45424 0 _0055_
rlabel metal1 4830 4624 4830 4624 0 _0056_
rlabel metal1 3404 25262 3404 25262 0 _0057_
rlabel metal1 2070 5270 2070 5270 0 _0058_
rlabel metal1 5474 6766 5474 6766 0 _0059_
rlabel metal1 2622 3060 2622 3060 0 _0060_
rlabel metal1 4370 6732 4370 6732 0 _0061_
rlabel metal1 16974 2584 16974 2584 0 _0062_
rlabel metal1 4094 36618 4094 36618 0 _0063_
rlabel metal1 20838 31790 20838 31790 0 _0064_
rlabel metal1 23966 35054 23966 35054 0 _0065_
rlabel metal1 23598 36550 23598 36550 0 _0066_
rlabel metal2 16606 32300 16606 32300 0 _0067_
rlabel metal1 18400 32878 18400 32878 0 _0068_
rlabel metal1 19090 32504 19090 32504 0 _0069_
rlabel metal1 21022 32980 21022 32980 0 _0070_
rlabel metal1 19826 26554 19826 26554 0 _0071_
rlabel metal2 20562 32640 20562 32640 0 _0072_
rlabel metal1 20562 33558 20562 33558 0 _0073_
rlabel metal1 21436 32878 21436 32878 0 _0074_
rlabel metal1 20562 33456 20562 33456 0 _0075_
rlabel metal2 21942 33082 21942 33082 0 _0076_
rlabel metal2 19182 32640 19182 32640 0 _0077_
rlabel metal1 16836 32878 16836 32878 0 _0078_
rlabel metal1 18538 32334 18538 32334 0 _0079_
rlabel metal1 18446 37876 18446 37876 0 _0080_
rlabel metal1 18354 33286 18354 33286 0 _0081_
rlabel metal1 19688 31994 19688 31994 0 _0082_
rlabel metal1 20194 32946 20194 32946 0 _0083_
rlabel metal2 19458 33320 19458 33320 0 _0084_
rlabel metal1 19320 32402 19320 32402 0 _0085_
rlabel metal2 18078 32572 18078 32572 0 _0086_
rlabel metal1 18653 32470 18653 32470 0 _0087_
rlabel metal1 19274 32198 19274 32198 0 _0088_
rlabel metal1 18262 13260 18262 13260 0 _0089_
rlabel metal1 19780 12614 19780 12614 0 _0090_
rlabel metal1 18768 10166 18768 10166 0 _0091_
rlabel metal1 17894 10676 17894 10676 0 _0092_
rlabel metal2 18262 11288 18262 11288 0 _0093_
rlabel metal2 18170 10268 18170 10268 0 _0094_
rlabel metal2 18262 10387 18262 10387 0 _0095_
rlabel metal1 17526 13294 17526 13294 0 _0096_
rlabel metal1 18676 13158 18676 13158 0 _0097_
rlabel metal2 19274 10812 19274 10812 0 _0098_
rlabel metal1 19044 11322 19044 11322 0 _0099_
rlabel metal1 18814 10778 18814 10778 0 _0100_
rlabel metal1 18860 11866 18860 11866 0 _0101_
rlabel metal2 18814 27404 18814 27404 0 _0102_
rlabel metal2 24702 18598 24702 18598 0 _0103_
rlabel metal2 26634 25262 26634 25262 0 _0104_
rlabel metal1 25622 27370 25622 27370 0 _0105_
rlabel metal1 23322 18598 23322 18598 0 _0106_
rlabel metal2 21482 27268 21482 27268 0 _0107_
rlabel metal2 21390 37094 21390 37094 0 _0108_
rlabel metal1 21022 28526 21022 28526 0 _0109_
rlabel metal1 21344 21862 21344 21862 0 _0110_
rlabel metal1 22218 31994 22218 31994 0 _0111_
rlabel metal1 15916 19754 15916 19754 0 _0112_
rlabel metal2 14490 19992 14490 19992 0 _0113_
rlabel metal1 16376 19414 16376 19414 0 _0114_
rlabel metal1 14398 17204 14398 17204 0 _0115_
rlabel via1 13455 18258 13455 18258 0 _0116_
rlabel metal2 14766 18020 14766 18020 0 _0117_
rlabel metal2 12282 18496 12282 18496 0 _0118_
rlabel metal1 12972 18938 12972 18938 0 _0119_
rlabel metal1 14904 20434 14904 20434 0 _0120_
rlabel metal1 14904 19482 14904 19482 0 _0121_
rlabel metal2 14674 18190 14674 18190 0 _0122_
rlabel metal2 14674 20230 14674 20230 0 _0123_
rlabel metal1 14076 17714 14076 17714 0 _0124_
rlabel metal2 14582 17612 14582 17612 0 _0125_
rlabel metal2 15410 20434 15410 20434 0 _0126_
rlabel metal2 24978 34850 24978 34850 0 _0127_
rlabel metal2 13110 20230 13110 20230 0 _0128_
rlabel metal1 23322 18258 23322 18258 0 _0129_
rlabel metal2 24518 29716 24518 29716 0 _0130_
rlabel metal2 24702 26044 24702 26044 0 _0131_
rlabel metal2 25116 31892 25116 31892 0 _0132_
rlabel metal2 24932 32878 24932 32878 0 _0133_
rlabel metal1 24334 28526 24334 28526 0 _0134_
rlabel metal1 25829 31790 25829 31790 0 _0135_
rlabel metal1 25070 21964 25070 21964 0 _0136_
rlabel metal1 24978 18938 24978 18938 0 _0137_
rlabel metal1 25208 20434 25208 20434 0 _0138_
rlabel metal1 21298 12240 21298 12240 0 _0139_
rlabel metal1 21022 21488 21022 21488 0 _0140_
rlabel metal1 24978 22168 24978 22168 0 _0141_
rlabel metal1 25116 23698 25116 23698 0 _0142_
rlabel metal1 24380 20366 24380 20366 0 _0143_
rlabel metal2 25162 21692 25162 21692 0 _0144_
rlabel metal2 25622 21114 25622 21114 0 _0145_
rlabel metal2 25622 24786 25622 24786 0 _0146_
rlabel metal2 26266 24242 26266 24242 0 _0147_
rlabel metal2 25806 24310 25806 24310 0 _0148_
rlabel metal1 25714 25296 25714 25296 0 _0149_
rlabel metal1 25760 25466 25760 25466 0 _0150_
rlabel metal2 25254 24990 25254 24990 0 _0151_
rlabel metal1 25438 23120 25438 23120 0 _0152_
rlabel metal1 25254 31790 25254 31790 0 _0153_
rlabel metal1 25760 31926 25760 31926 0 _0154_
rlabel metal1 26864 25738 26864 25738 0 _0155_
rlabel metal1 26404 30702 26404 30702 0 _0156_
rlabel metal1 25438 28526 25438 28526 0 _0157_
rlabel metal1 24288 29478 24288 29478 0 _0158_
rlabel metal1 24748 29070 24748 29070 0 _0159_
rlabel metal2 25898 27268 25898 27268 0 _0160_
rlabel metal1 25070 27642 25070 27642 0 _0161_
rlabel metal2 25714 28220 25714 28220 0 _0162_
rlabel metal2 24610 28934 24610 28934 0 _0163_
rlabel metal1 23414 29274 23414 29274 0 _0164_
rlabel metal2 23966 25466 23966 25466 0 _0165_
rlabel metal1 23184 29614 23184 29614 0 _0166_
rlabel metal1 21666 15130 21666 15130 0 _0167_
rlabel metal1 20792 16082 20792 16082 0 _0168_
rlabel metal1 16790 36686 16790 36686 0 _0169_
rlabel metal1 19872 17034 19872 17034 0 _0170_
rlabel metal1 18630 17850 18630 17850 0 _0171_
rlabel metal1 20746 12818 20746 12818 0 _0172_
rlabel metal1 20516 12954 20516 12954 0 _0173_
rlabel metal1 19780 13498 19780 13498 0 _0174_
rlabel metal2 19458 14212 19458 14212 0 _0175_
rlabel metal1 21574 18258 21574 18258 0 _0176_
rlabel metal1 21252 18394 21252 18394 0 _0177_
rlabel metal1 19642 25296 19642 25296 0 _0178_
rlabel metal1 19090 25262 19090 25262 0 _0179_
rlabel metal1 19044 23086 19044 23086 0 _0180_
rlabel metal2 18814 23732 18814 23732 0 _0181_
rlabel metal2 19550 20740 19550 20740 0 _0182_
rlabel metal2 18722 20604 18722 20604 0 _0183_
rlabel metal1 24150 36210 24150 36210 0 _0184_
rlabel metal2 16882 23902 16882 23902 0 _0185_
rlabel metal2 17250 24310 17250 24310 0 _0186_
rlabel metal2 16146 25466 16146 25466 0 _0187_
rlabel metal1 16744 25262 16744 25262 0 _0188_
rlabel metal2 23138 35530 23138 35530 0 _0189_
rlabel metal1 23092 36142 23092 36142 0 _0190_
rlabel metal2 23690 31994 23690 31994 0 _0191_
rlabel metal1 23368 31994 23368 31994 0 _0192_
rlabel metal1 17250 36754 17250 36754 0 _0193_
rlabel metal2 17802 36346 17802 36346 0 _0194_
rlabel metal2 16330 21114 16330 21114 0 _0195_
rlabel metal1 16284 21114 16284 21114 0 _0196_
rlabel metal1 16330 35666 16330 35666 0 _0197_
rlabel metal1 16790 36142 16790 36142 0 _0198_
rlabel metal1 15640 27030 15640 27030 0 _0199_
rlabel metal1 16422 26962 16422 26962 0 _0200_
rlabel metal1 16790 11866 16790 11866 0 _0201_
rlabel metal1 17204 12206 17204 12206 0 _0202_
rlabel metal1 26726 15130 26726 15130 0 _0203_
rlabel metal1 26910 16082 26910 16082 0 _0204_
rlabel metal2 16146 22202 16146 22202 0 _0205_
rlabel metal1 16100 22202 16100 22202 0 _0206_
rlabel metal2 25898 13124 25898 13124 0 _0207_
rlabel metal2 25622 13702 25622 13702 0 _0208_
rlabel metal1 21110 29274 21110 29274 0 _0209_
rlabel metal1 21436 21998 21436 21998 0 _0210_
rlabel metal1 22678 20570 22678 20570 0 _0211_
rlabel metal2 22770 21692 22770 21692 0 _0212_
rlabel metal2 21298 25772 21298 25772 0 _0213_
rlabel metal2 22402 25092 22402 25092 0 _0214_
rlabel metal2 21482 23596 21482 23596 0 _0215_
rlabel metal1 21712 23290 21712 23290 0 _0216_
rlabel metal1 21252 21522 21252 21522 0 _0217_
rlabel metal1 21252 21386 21252 21386 0 _0218_
rlabel metal2 24242 18564 24242 18564 0 _0219_
rlabel metal1 23230 17646 23230 17646 0 _0220_
rlabel metal2 24610 17000 24610 17000 0 _0221_
rlabel metal2 23230 17884 23230 17884 0 _0222_
rlabel metal2 23506 17034 23506 17034 0 _0223_
rlabel metal1 23368 12886 23368 12886 0 _0224_
rlabel metal2 23782 13430 23782 13430 0 _0225_
rlabel metal1 22448 12954 22448 12954 0 _0226_
rlabel metal2 22310 13634 22310 13634 0 _0227_
rlabel metal1 21850 13838 21850 13838 0 _0228_
rlabel metal1 24748 13498 24748 13498 0 _0229_
rlabel metal1 24367 13158 24367 13158 0 _0230_
rlabel metal2 24610 13702 24610 13702 0 _0231_
rlabel metal2 19642 29818 19642 29818 0 _0232_
rlabel metal1 20056 38454 20056 38454 0 _0233_
rlabel metal1 16882 18938 16882 18938 0 _0234_
rlabel metal2 18078 37026 18078 37026 0 _0235_
rlabel metal2 20470 37808 20470 37808 0 _0236_
rlabel metal1 20654 38522 20654 38522 0 _0237_
rlabel metal1 21712 38522 21712 38522 0 _0238_
rlabel metal1 21268 38250 21268 38250 0 _0239_
rlabel metal1 21712 37842 21712 37842 0 _0240_
rlabel metal1 19688 37842 19688 37842 0 _0241_
rlabel metal1 18630 37808 18630 37808 0 _0242_
rlabel metal1 19198 38250 19198 38250 0 _0243_
rlabel metal1 18952 38522 18952 38522 0 _0244_
rlabel metal2 18262 37536 18262 37536 0 _0245_
rlabel metal1 18876 37162 18876 37162 0 _0246_
rlabel metal2 18446 36924 18446 36924 0 _0247_
rlabel metal1 15456 32198 15456 32198 0 _0248_
rlabel metal1 15740 32538 15740 32538 0 _0249_
rlabel metal1 16721 32402 16721 32402 0 _0250_
rlabel metal2 16054 31280 16054 31280 0 _0251_
rlabel metal1 16016 30634 16016 30634 0 _0252_
rlabel metal1 16192 30226 16192 30226 0 _0253_
rlabel metal1 15916 17646 15916 17646 0 _0254_
rlabel metal1 16054 28458 16054 28458 0 _0255_
rlabel metal1 16468 28730 16468 28730 0 _0256_
rlabel metal1 16330 18258 16330 18258 0 _0257_
rlabel metal1 16238 17850 16238 17850 0 _0258_
rlabel metal2 16330 18870 16330 18870 0 _0259_
rlabel metal1 15824 16762 15824 16762 0 _0260_
rlabel metal2 17250 18496 17250 18496 0 _0261_
rlabel metal1 16422 18938 16422 18938 0 _0262_
rlabel metal1 16744 14586 16744 14586 0 _0263_
rlabel metal1 16706 14246 16706 14246 0 _0264_
rlabel metal1 17480 14382 17480 14382 0 _0265_
rlabel metal2 23322 24140 23322 24140 0 _0266_
rlabel metal2 6762 3706 6762 3706 0 _0267_
rlabel metal2 3082 35428 3082 35428 0 _0268_
rlabel metal2 17066 3230 17066 3230 0 _0269_
rlabel metal2 4738 7582 4738 7582 0 _0270_
rlabel metal1 26358 6698 26358 6698 0 _0271_
rlabel metal2 3082 5950 3082 5950 0 _0272_
rlabel metal1 27002 26010 27002 26010 0 _0273_
rlabel metal2 1886 3604 1886 3604 0 _0274_
rlabel metal2 26450 38930 26450 38930 0 _0275_
rlabel metal2 26450 45934 26450 45934 0 _0276_
rlabel metal2 26726 18156 26726 18156 0 _0277_
rlabel metal2 17250 3196 17250 3196 0 _0278_
rlabel metal1 26036 43418 26036 43418 0 _0279_
rlabel metal1 3726 43962 3726 43962 0 _0280_
rlabel metal2 11822 45730 11822 45730 0 _0281_
rlabel metal2 4094 9214 4094 9214 0 _0282_
rlabel metal2 26726 23324 26726 23324 0 _0283_
rlabel metal2 26726 38556 26726 38556 0 _0284_
rlabel metal2 2990 39134 2990 39134 0 _0285_
rlabel metal2 28106 32674 28106 32674 0 _0286_
rlabel metal1 2116 8058 2116 8058 0 _0287_
rlabel metal2 27278 44642 27278 44642 0 _0288_
rlabel metal2 14582 46308 14582 46308 0 _0289_
rlabel metal2 9154 3230 9154 3230 0 _0290_
rlabel metal2 28198 25058 28198 25058 0 _0291_
rlabel metal2 2530 3298 2530 3298 0 _0292_
rlabel metal2 28198 14892 28198 14892 0 _0293_
rlabel metal2 1794 38828 1794 38828 0 _0294_
rlabel metal2 28198 5916 28198 5916 0 _0295_
rlabel metal2 4186 6494 4186 6494 0 _0296_
rlabel metal2 28198 20706 28198 20706 0 _0297_
rlabel metal1 25162 45050 25162 45050 0 _0298_
rlabel metal1 26634 39066 26634 39066 0 _0299_
rlabel metal2 16422 46308 16422 46308 0 _0300_
rlabel metal2 5290 3026 5290 3026 0 _0301_
rlabel metal1 2024 34170 2024 34170 0 _0302_
rlabel metal1 26358 34986 26358 34986 0 _0303_
rlabel metal2 7866 46308 7866 46308 0 _0304_
rlabel metal1 25852 46614 25852 46614 0 _0305_
rlabel metal2 2254 15844 2254 15844 0 _0306_
rlabel metal1 14444 2618 14444 2618 0 _0307_
rlabel metal1 11914 15538 11914 15538 0 _0308_
rlabel metal2 26726 32028 26726 32028 0 _0309_
rlabel metal2 12098 3740 12098 3740 0 _0310_
rlabel metal1 6578 6834 6578 6834 0 _0311_
rlabel metal2 25898 4012 25898 4012 0 _0312_
rlabel metal1 26128 36074 26128 36074 0 _0313_
rlabel metal1 9660 30770 9660 30770 0 _0314_
rlabel metal2 27278 33762 27278 33762 0 _0315_
rlabel metal2 27278 45730 27278 45730 0 _0316_
rlabel metal1 27002 6426 27002 6426 0 _0317_
rlabel metal1 2208 18938 2208 18938 0 _0318_
rlabel metal1 22356 45594 22356 45594 0 _0319_
rlabel metal2 2070 32164 2070 32164 0 _0320_
rlabel metal2 24518 3230 24518 3230 0 _0321_
rlabel metal2 27738 29410 27738 29410 0 _0322_
rlabel metal2 22218 3230 22218 3230 0 _0323_
rlabel metal1 19550 45594 19550 45594 0 _0324_
rlabel metal1 1886 5338 1886 5338 0 _0325_
rlabel metal2 22402 45968 22402 45968 0 _0326_
rlabel metal2 13018 4590 13018 4590 0 _0327_
rlabel metal2 26726 11356 26726 11356 0 _0328_
rlabel metal1 1932 4794 1932 4794 0 _0329_
rlabel metal2 1886 11492 1886 11492 0 _0330_
rlabel metal1 2346 37230 2346 37230 0 _0331_
rlabel metal2 26726 16796 26726 16796 0 _0332_
rlabel metal2 26450 42670 26450 42670 0 _0333_
rlabel metal1 27048 41514 27048 41514 0 _0334_
rlabel metal2 4094 46308 4094 46308 0 _0335_
rlabel metal2 26450 44846 26450 44846 0 _0336_
rlabel metal2 20654 7004 20654 7004 0 _0337_
rlabel metal1 27002 4250 27002 4250 0 _0338_
rlabel metal2 23046 46240 23046 46240 0 _0339_
rlabel metal2 19458 3230 19458 3230 0 _0340_
rlabel metal1 28014 9690 28014 9690 0 _0341_
rlabel metal2 2438 25636 2438 25636 0 _0342_
rlabel metal2 27370 23426 27370 23426 0 _0343_
rlabel metal1 2898 42738 2898 42738 0 _0344_
rlabel metal2 4186 4318 4186 4318 0 _0345_
rlabel metal1 7820 3978 7820 3978 0 _0346_
rlabel metal2 1978 13090 1978 13090 0 _0347_
rlabel metal2 28198 30940 28198 30940 0 _0348_
rlabel metal2 28014 18530 28014 18530 0 _0349_
rlabel metal2 28198 21794 28198 21794 0 _0350_
rlabel metal1 4600 2346 4600 2346 0 _0351_
rlabel metal2 3634 43758 3634 43758 0 _0352_
rlabel metal1 27048 12614 27048 12614 0 _0353_
rlabel metal2 11914 3230 11914 3230 0 _0354_
rlabel metal1 18952 46138 18952 46138 0 _0355_
rlabel metal1 2944 45526 2944 45526 0 _0356_
rlabel metal2 27922 27234 27922 27234 0 _0357_
rlabel metal2 2254 40868 2254 40868 0 _0358_
rlabel metal1 4002 2618 4002 2618 0 _0359_
rlabel metal2 9890 46546 9890 46546 0 _0360_
rlabel metal2 10534 46308 10534 46308 0 _0361_
rlabel metal2 26450 7582 26450 7582 0 _0362_
rlabel metal2 27830 42466 27830 42466 0 _0363_
rlabel metal2 13570 46308 13570 46308 0 _0364_
rlabel metal1 27278 3706 27278 3706 0 _0365_
rlabel metal2 27922 37026 27922 37026 0 _0366_
rlabel metal2 3266 41820 3266 41820 0 _0367_
rlabel metal2 26450 2652 26450 2652 0 _0368_
rlabel metal2 1794 20060 1794 20060 0 _0369_
rlabel metal2 27278 8738 27278 8738 0 _0370_
rlabel metal2 1978 45730 1978 45730 0 _0371_
rlabel metal2 2438 17442 2438 17442 0 _0372_
rlabel metal2 1886 9044 1886 9044 0 _0373_
rlabel metal2 2898 14178 2898 14178 0 _0374_
rlabel metal3 1786 36788 1786 36788 0 active
rlabel metal2 22586 17986 22586 17986 0 clknet_0_wb_clk_i
rlabel metal1 16836 21522 16836 21522 0 clknet_2_0__leaf_wb_clk_i
rlabel metal1 21758 20978 21758 20978 0 clknet_2_1__leaf_wb_clk_i
rlabel metal1 19780 35054 19780 35054 0 clknet_2_2__leaf_wb_clk_i
rlabel metal1 22080 32402 22080 32402 0 clknet_2_3__leaf_wb_clk_i
rlabel metal1 20976 37230 20976 37230 0 frequency_counter_0.clk_counter\[0\]
rlabel metal1 16652 13906 16652 13906 0 frequency_counter_0.clk_counter\[10\]
rlabel metal1 18630 13906 18630 13906 0 frequency_counter_0.clk_counter\[11\]
rlabel metal1 20700 37230 20700 37230 0 frequency_counter_0.clk_counter\[1\]
rlabel metal1 21850 38250 21850 38250 0 frequency_counter_0.clk_counter\[2\]
rlabel metal1 20608 37706 20608 37706 0 frequency_counter_0.clk_counter\[3\]
rlabel metal1 19596 34578 19596 34578 0 frequency_counter_0.clk_counter\[4\]
rlabel metal2 18354 31484 18354 31484 0 frequency_counter_0.clk_counter\[5\]
rlabel metal1 18124 30362 18124 30362 0 frequency_counter_0.clk_counter\[6\]
rlabel metal1 18308 29818 18308 29818 0 frequency_counter_0.clk_counter\[7\]
rlabel metal1 16928 16762 16928 16762 0 frequency_counter_0.clk_counter\[8\]
rlabel metal1 17618 16490 17618 16490 0 frequency_counter_0.clk_counter\[9\]
rlabel metal1 24794 35020 24794 35020 0 frequency_counter_0.digit
rlabel metal2 23782 20298 23782 20298 0 frequency_counter_0.edge_counter\[0\]
rlabel metal1 26864 18258 26864 18258 0 frequency_counter_0.edge_counter\[1\]
rlabel metal1 25921 20910 25921 20910 0 frequency_counter_0.edge_counter\[2\]
rlabel metal1 24472 23630 24472 23630 0 frequency_counter_0.edge_counter\[3\]
rlabel metal2 26174 27438 26174 27438 0 frequency_counter_0.edge_counter\[4\]
rlabel metal2 26174 29376 26174 29376 0 frequency_counter_0.edge_counter\[5\]
rlabel metal2 23506 29274 23506 29274 0 frequency_counter_0.edge_counter\[6\]
rlabel metal2 24794 36380 24794 36380 0 frequency_counter_0.edge_detect0.q0
rlabel metal1 24886 34000 24886 34000 0 frequency_counter_0.edge_detect0.q1
rlabel metal1 25024 32878 25024 32878 0 frequency_counter_0.edge_detect0.q2
rlabel metal1 13340 15538 13340 15538 0 frequency_counter_0.segments\[0\]
rlabel metal1 26450 31790 26450 31790 0 frequency_counter_0.segments\[1\]
rlabel metal2 11914 10880 11914 10880 0 frequency_counter_0.segments\[2\]
rlabel metal1 7820 6834 7820 6834 0 frequency_counter_0.segments\[3\]
rlabel metal1 25714 3604 25714 3604 0 frequency_counter_0.segments\[4\]
rlabel metal1 25622 35258 25622 35258 0 frequency_counter_0.segments\[5\]
rlabel metal1 11822 30702 11822 30702 0 frequency_counter_0.segments\[6\]
rlabel metal1 20056 20366 20056 20366 0 frequency_counter_0.seven_segment0.load
rlabel metal1 22962 14042 22962 14042 0 frequency_counter_0.seven_segment0.ten_count\[0\]
rlabel metal2 23046 17476 23046 17476 0 frequency_counter_0.seven_segment0.ten_count\[1\]
rlabel metal1 21827 13294 21827 13294 0 frequency_counter_0.seven_segment0.ten_count\[2\]
rlabel metal1 20378 13396 20378 13396 0 frequency_counter_0.seven_segment0.ten_count\[3\]
rlabel metal2 22586 16830 22586 16830 0 frequency_counter_0.seven_segment0.ten_count_reg\[0\]
rlabel metal1 19872 17306 19872 17306 0 frequency_counter_0.seven_segment0.ten_count_reg\[1\]
rlabel metal1 19320 14858 19320 14858 0 frequency_counter_0.seven_segment0.ten_count_reg\[2\]
rlabel metal2 20838 17136 20838 17136 0 frequency_counter_0.seven_segment0.ten_count_reg\[3\]
rlabel metal1 22632 20366 22632 20366 0 frequency_counter_0.seven_segment0.unit_count\[0\]
rlabel metal1 21206 26418 21206 26418 0 frequency_counter_0.seven_segment0.unit_count\[1\]
rlabel metal2 20102 24004 20102 24004 0 frequency_counter_0.seven_segment0.unit_count\[2\]
rlabel metal2 19734 21556 19734 21556 0 frequency_counter_0.seven_segment0.unit_count\[3\]
rlabel metal1 22310 18394 22310 18394 0 frequency_counter_0.seven_segment0.unit_count_reg\[0\]
rlabel metal1 20148 17714 20148 17714 0 frequency_counter_0.seven_segment0.unit_count_reg\[1\]
rlabel metal1 19734 23086 19734 23086 0 frequency_counter_0.seven_segment0.unit_count_reg\[2\]
rlabel metal1 20010 20570 20010 20570 0 frequency_counter_0.seven_segment0.unit_count_reg\[3\]
rlabel metal1 21850 36754 21850 36754 0 frequency_counter_0.state\[0\]
rlabel metal1 21758 31790 21758 31790 0 frequency_counter_0.state\[1\]
rlabel metal2 24426 30974 24426 30974 0 frequency_counter_0.state\[2\]
rlabel metal1 18814 24378 18814 24378 0 frequency_counter_0.update_period\[0\]
rlabel metal2 18354 13396 18354 13396 0 frequency_counter_0.update_period\[10\]
rlabel metal2 18078 13600 18078 13600 0 frequency_counter_0.update_period\[11\]
rlabel metal1 19090 26010 19090 26010 0 frequency_counter_0.update_period\[1\]
rlabel metal1 23644 36006 23644 36006 0 frequency_counter_0.update_period\[2\]
rlabel metal2 24058 33286 24058 33286 0 frequency_counter_0.update_period\[3\]
rlabel metal1 17618 37162 17618 37162 0 frequency_counter_0.update_period\[4\]
rlabel metal1 18630 32810 18630 32810 0 frequency_counter_0.update_period\[5\]
rlabel metal2 18078 33133 18078 33133 0 frequency_counter_0.update_period\[6\]
rlabel metal2 17940 32980 17940 32980 0 frequency_counter_0.update_period\[7\]
rlabel metal1 17756 15878 17756 15878 0 frequency_counter_0.update_period\[8\]
rlabel metal1 19918 10030 19918 10030 0 frequency_counter_0.update_period\[9\]
rlabel via2 27370 36771 27370 36771 0 io_in[8]
rlabel metal2 21298 2710 21298 2710 0 io_oeb[0]
rlabel metal3 1142 13668 1142 13668 0 io_oeb[10]
rlabel metal3 28405 32300 28405 32300 0 io_oeb[11]
rlabel metal1 26358 18802 26358 18802 0 io_oeb[12]
rlabel metal2 27554 21607 27554 21607 0 io_oeb[13]
rlabel metal3 1740 3468 1740 3468 0 io_oeb[14]
rlabel metal1 1012 43350 1012 43350 0 io_oeb[15]
rlabel metal3 28850 12308 28850 12308 0 io_oeb[16]
rlabel metal1 11592 2958 11592 2958 0 io_oeb[17]
rlabel metal1 19642 46444 19642 46444 0 io_oeb[18]
rlabel metal2 1978 48188 1978 48188 0 io_oeb[19]
rlabel metal3 28436 1428 28436 1428 0 io_oeb[1]
rlabel via2 27554 27523 27554 27523 0 io_oeb[20]
rlabel metal2 2806 41293 2806 41293 0 io_oeb[21]
rlabel metal1 4094 2958 4094 2958 0 io_oeb[22]
rlabel metal2 10350 48188 10350 48188 0 io_oeb[23]
rlabel metal2 10994 47882 10994 47882 0 io_oeb[24]
rlabel metal2 26174 7769 26174 7769 0 io_oeb[25]
rlabel metal1 26358 42602 26358 42602 0 io_oeb[26]
rlabel metal2 13478 47209 13478 47209 0 io_oeb[27]
rlabel metal2 26174 3757 26174 3757 0 io_oeb[28]
rlabel metal2 26174 36635 26174 36635 0 io_oeb[29]
rlabel metal2 23230 48188 23230 48188 0 io_oeb[2]
rlabel metal3 1142 42228 1142 42228 0 io_oeb[30]
rlabel metal2 26174 2635 26174 2635 0 io_oeb[31]
rlabel metal3 1740 19788 1740 19788 0 io_oeb[32]
rlabel metal3 28850 8908 28850 8908 0 io_oeb[33]
rlabel metal2 2990 47855 2990 47855 0 io_oeb[34]
rlabel via2 2806 17731 2806 17731 0 io_oeb[35]
rlabel metal3 1740 8908 1740 8908 0 io_oeb[36]
rlabel metal3 1142 14348 1142 14348 0 io_oeb[37]
rlabel metal2 20010 1860 20010 1860 0 io_oeb[3]
rlabel metal2 27554 10183 27554 10183 0 io_oeb[4]
rlabel metal3 1740 25908 1740 25908 0 io_oeb[5]
rlabel metal3 28850 24548 28850 24548 0 io_oeb[6]
rlabel metal1 874 43826 874 43826 0 io_oeb[7]
rlabel metal1 4140 3978 4140 3978 0 io_oeb[8]
rlabel metal2 8418 2404 8418 2404 0 io_oeb[9]
rlabel metal1 28520 40562 28520 40562 0 io_out[0]
rlabel metal3 28850 32028 28850 32028 0 io_out[10]
rlabel metal2 12466 2924 12466 2924 0 io_out[11]
rlabel metal3 2384 6188 2384 6188 0 io_out[12]
rlabel metal3 29823 2108 29823 2108 0 io_out[13]
rlabel metal3 28390 42228 28390 42228 0 io_out[14]
rlabel metal3 2108 33388 2108 33388 0 io_out[15]
rlabel metal1 26726 34068 26726 34068 0 io_out[16]
rlabel metal1 27048 46002 27048 46002 0 io_out[17]
rlabel metal3 29846 7548 29846 7548 0 io_out[18]
rlabel metal3 1418 19108 1418 19108 0 io_out[19]
rlabel metal1 17342 46444 17342 46444 0 io_out[1]
rlabel metal2 22586 47644 22586 47644 0 io_out[20]
rlabel metal3 1740 32028 1740 32028 0 io_out[21]
rlabel metal2 25162 1860 25162 1860 0 io_out[22]
rlabel metal2 27554 29155 27554 29155 0 io_out[23]
rlabel metal2 21942 1231 21942 1231 0 io_out[24]
rlabel metal2 20010 47644 20010 47644 0 io_out[25]
rlabel metal3 1740 4148 1740 4148 0 io_out[26]
rlabel metal2 21298 47848 21298 47848 0 io_out[27]
rlabel metal2 13570 2404 13570 2404 0 io_out[28]
rlabel metal3 29846 10948 29846 10948 0 io_out[29]
rlabel metal2 5842 2166 5842 2166 0 io_out[2]
rlabel metal3 1924 4828 1924 4828 0 io_out[30]
rlabel metal3 1740 11628 1740 11628 0 io_out[31]
rlabel metal3 1188 37468 1188 37468 0 io_out[32]
rlabel metal3 28988 15708 28988 15708 0 io_out[33]
rlabel metal2 26082 42517 26082 42517 0 io_out[34]
rlabel metal3 28436 40868 28436 40868 0 io_out[35]
rlabel metal1 4186 46444 4186 46444 0 io_out[36]
rlabel metal2 26082 45305 26082 45305 0 io_out[37]
rlabel metal2 2806 34629 2806 34629 0 io_out[3]
rlabel metal3 28436 34068 28436 34068 0 io_out[4]
rlabel metal2 8418 47882 8418 47882 0 io_out[5]
rlabel metal2 28382 47882 28382 47882 0 io_out[6]
rlabel metal3 1740 15708 1740 15708 0 io_out[7]
rlabel metal2 14858 1231 14858 1231 0 io_out[8]
rlabel metal3 2108 12308 2108 12308 0 io_out[9]
rlabel metal1 29164 16082 29164 16082 0 la1_data_in[0]
rlabel metal2 17434 1367 17434 1367 0 la1_data_in[10]
rlabel metal2 25530 15249 25530 15249 0 la1_data_in[11]
rlabel metal3 1142 29988 1142 29988 0 la1_data_in[12]
rlabel metal2 27094 1588 27094 1588 0 la1_data_in[13]
rlabel metal2 16146 1554 16146 1554 0 la1_data_in[1]
rlabel metal2 9062 1588 9062 1588 0 la1_data_in[2]
rlabel metal3 1142 25228 1142 25228 0 la1_data_in[3]
rlabel metal1 24334 45934 24334 45934 0 la1_data_in[4]
rlabel metal2 26634 30107 26634 30107 0 la1_data_in[5]
rlabel metal2 5842 48154 5842 48154 0 la1_data_in[6]
rlabel metal3 1142 18428 1142 18428 0 la1_data_in[7]
rlabel metal1 6532 47022 6532 47022 0 la1_data_in[8]
rlabel metal3 1142 27948 1142 27948 0 la1_data_in[9]
rlabel metal1 6693 2890 6693 2890 0 la1_data_out[0]
rlabel metal3 28988 19788 28988 19788 0 la1_data_out[10]
rlabel metal2 18078 1622 18078 1622 0 la1_data_out[11]
rlabel metal3 27746 46988 27746 46988 0 la1_data_out[12]
rlabel metal3 2154 44268 2154 44268 0 la1_data_out[13]
rlabel metal2 11822 46767 11822 46767 0 la1_data_out[14]
rlabel metal3 2016 1428 2016 1428 0 la1_data_out[15]
rlabel metal3 29846 23868 29846 23868 0 la1_data_out[16]
rlabel metal3 28988 39508 28988 39508 0 la1_data_out[17]
rlabel metal2 4278 41905 4278 41905 0 la1_data_out[18]
rlabel metal3 28436 30668 28436 30668 0 la1_data_out[19]
rlabel metal3 1188 36108 1188 36108 0 la1_data_out[1]
rlabel metal3 1832 8228 1832 8228 0 la1_data_out[20]
rlabel metal3 28850 44948 28850 44948 0 la1_data_out[21]
rlabel metal1 14812 46478 14812 46478 0 la1_data_out[22]
rlabel metal2 9706 1860 9706 1860 0 la1_data_out[23]
rlabel metal2 27554 25279 27554 25279 0 la1_data_out[24]
rlabel metal3 1142 2788 1142 2788 0 la1_data_out[25]
rlabel metal2 27554 14399 27554 14399 0 la1_data_out[26]
rlabel metal2 2806 38607 2806 38607 0 la1_data_out[27]
rlabel metal2 27554 5491 27554 5491 0 la1_data_out[28]
rlabel metal1 4416 6222 4416 6222 0 la1_data_out[29]
rlabel metal1 17066 2958 17066 2958 0 la1_data_out[2]
rlabel metal2 27554 20723 27554 20723 0 la1_data_out[30]
rlabel metal3 27976 49028 27976 49028 0 la1_data_out[31]
rlabel metal3 1878 7548 1878 7548 0 la1_data_out[3]
rlabel metal3 28850 6868 28850 6868 0 la1_data_out[4]
rlabel metal2 2622 1792 2622 1792 0 la1_data_out[5]
rlabel metal3 28850 26588 28850 26588 0 la1_data_out[6]
rlabel metal2 690 2404 690 2404 0 la1_data_out[7]
rlabel metal3 29846 40188 29846 40188 0 la1_data_out[8]
rlabel metal1 26818 45390 26818 45390 0 la1_data_out[9]
rlabel metal2 1610 36890 1610 36890 0 net1
rlabel metal2 1794 25024 1794 25024 0 net10
rlabel metal2 1702 41548 1702 41548 0 net100
rlabel metal1 3496 2958 3496 2958 0 net101
rlabel metal1 9522 45458 9522 45458 0 net102
rlabel metal1 9844 46410 9844 46410 0 net103
rlabel metal2 26634 7820 26634 7820 0 net104
rlabel metal1 28244 42738 28244 42738 0 net105
rlabel metal2 13938 46784 13938 46784 0 net106
rlabel metal1 27278 4046 27278 4046 0 net107
rlabel metal1 28336 36346 28336 36346 0 net108
rlabel metal2 3450 42126 3450 42126 0 net109
rlabel metal1 24104 45798 24104 45798 0 net11
rlabel metal1 27232 2482 27232 2482 0 net110
rlabel metal2 1610 20060 1610 20060 0 net111
rlabel metal1 27830 8500 27830 8500 0 net112
rlabel metal2 1610 46172 1610 46172 0 net113
rlabel metal1 1656 17170 1656 17170 0 net114
rlabel metal2 1702 9792 1702 9792 0 net115
rlabel metal1 2346 13940 2346 13940 0 net116
rlabel metal1 25530 36006 25530 36006 0 net117
rlabel metal1 25990 33456 25990 33456 0 net118
rlabel metal1 25438 32470 25438 32470 0 net12
rlabel metal2 6026 42058 6026 42058 0 net13
rlabel metal2 15226 19822 15226 19822 0 net14
rlabel metal2 6762 41446 6762 41446 0 net15
rlabel metal2 1794 27608 1794 27608 0 net16
rlabel metal2 6578 3468 6578 3468 0 net17
rlabel metal1 2760 36210 2760 36210 0 net18
rlabel metal1 16606 3026 16606 3026 0 net19
rlabel metal1 26460 36754 26460 36754 0 net2
rlabel metal2 4922 7582 4922 7582 0 net20
rlabel metal1 26864 6834 26864 6834 0 net21
rlabel metal2 2898 5984 2898 5984 0 net22
rlabel metal2 26542 26588 26542 26588 0 net23
rlabel metal1 4232 4046 4232 4046 0 net24
rlabel metal1 27232 39474 27232 39474 0 net25
rlabel metal1 26680 45458 26680 45458 0 net26
rlabel metal1 26542 17748 26542 17748 0 net27
rlabel metal1 17066 2516 17066 2516 0 net28
rlabel metal2 25898 44336 25898 44336 0 net29
rlabel metal1 26128 16490 26128 16490 0 net3
rlabel metal2 3174 44608 3174 44608 0 net30
rlabel metal1 11454 46002 11454 46002 0 net31
rlabel metal2 4278 8908 4278 8908 0 net32
rlabel metal1 26542 23188 26542 23188 0 net33
rlabel metal2 26542 38590 26542 38590 0 net34
rlabel metal2 2806 39168 2806 39168 0 net35
rlabel metal1 26588 32402 26588 32402 0 net36
rlabel metal1 1656 8058 1656 8058 0 net37
rlabel metal2 27830 44540 27830 44540 0 net38
rlabel metal2 14398 46784 14398 46784 0 net39
rlabel metal2 18078 7718 18078 7718 0 net4
rlabel metal2 8970 3264 8970 3264 0 net40
rlabel metal2 28382 25500 28382 25500 0 net41
rlabel metal1 3312 3570 3312 3570 0 net42
rlabel metal1 28244 13906 28244 13906 0 net43
rlabel metal1 1610 38420 1610 38420 0 net44
rlabel metal1 28244 5202 28244 5202 0 net45
rlabel metal1 4048 5882 4048 5882 0 net46
rlabel metal1 28014 20366 28014 20366 0 net47
rlabel metal2 24794 46036 24794 46036 0 net48
rlabel metal2 26542 40732 26542 40732 0 net49
rlabel metal1 27508 15130 27508 15130 0 net5
rlabel metal2 16882 46784 16882 46784 0 net50
rlabel metal1 4876 3502 4876 3502 0 net51
rlabel metal1 1748 33490 1748 33490 0 net52
rlabel metal2 26542 35292 26542 35292 0 net53
rlabel metal2 7038 46784 7038 46784 0 net54
rlabel metal2 24334 45968 24334 45968 0 net55
rlabel metal1 1748 16558 1748 16558 0 net56
rlabel metal2 14306 3264 14306 3264 0 net57
rlabel metal2 27462 46512 27462 46512 0 net58
rlabel metal2 27830 7548 27830 7548 0 net59
rlabel metal1 1840 30022 1840 30022 0 net6
rlabel metal1 1748 18938 1748 18938 0 net60
rlabel metal2 22218 46614 22218 46614 0 net61
rlabel metal2 1702 32640 1702 32640 0 net62
rlabel metal2 24334 3264 24334 3264 0 net63
rlabel metal2 28382 29852 28382 29852 0 net64
rlabel metal1 21804 3026 21804 3026 0 net65
rlabel metal1 19734 45458 19734 45458 0 net66
rlabel metal2 1610 6256 1610 6256 0 net67
rlabel metal1 21436 46546 21436 46546 0 net68
rlabel metal2 12834 4352 12834 4352 0 net69
rlabel metal1 27140 2618 27140 2618 0 net7
rlabel metal1 26864 10642 26864 10642 0 net70
rlabel metal1 1748 7174 1748 7174 0 net71
rlabel metal2 1702 11968 1702 11968 0 net72
rlabel metal1 3772 37774 3772 37774 0 net73
rlabel metal1 26542 16660 26542 16660 0 net74
rlabel metal1 26956 42194 26956 42194 0 net75
rlabel metal1 27232 41446 27232 41446 0 net76
rlabel metal1 2760 46478 2760 46478 0 net77
rlabel metal1 27094 44302 27094 44302 0 net78
rlabel metal1 20516 4114 20516 4114 0 net79
rlabel metal1 16560 2618 16560 2618 0 net8
rlabel metal1 26864 3026 26864 3026 0 net80
rlabel metal2 22494 46070 22494 46070 0 net81
rlabel metal2 19274 3264 19274 3264 0 net82
rlabel metal2 28382 10268 28382 10268 0 net83
rlabel metal1 1748 26350 1748 26350 0 net84
rlabel metal2 27922 23426 27922 23426 0 net85
rlabel metal1 3266 43826 3266 43826 0 net86
rlabel metal2 4002 4352 4002 4352 0 net87
rlabel metal1 7820 3706 7820 3706 0 net88
rlabel metal2 3450 13532 3450 13532 0 net89
rlabel metal1 12650 24038 12650 24038 0 net9
rlabel metal1 28198 33286 28198 33286 0 net90
rlabel metal2 28382 18972 28382 18972 0 net91
rlabel metal1 27646 21556 27646 21556 0 net92
rlabel metal2 4048 3060 4048 3060 0 net93
rlabel metal1 4232 43282 4232 43282 0 net94
rlabel metal1 27232 12682 27232 12682 0 net95
rlabel metal2 11730 3264 11730 3264 0 net96
rlabel metal1 18860 46546 18860 46546 0 net97
rlabel metal1 3450 45458 3450 45458 0 net98
rlabel metal1 28290 27506 28290 27506 0 net99
rlabel metal1 24380 25942 24380 25942 0 wb_clk_i
<< properties >>
string FIXED_BBOX 0 0 30000 50000
<< end >>
