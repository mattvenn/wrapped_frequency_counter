magic
tech sky130A
magscale 1 2
timestamp 1647457561
<< viali >>
rect 23213 47073 23247 47107
rect 25973 47073 26007 47107
rect 1777 47005 1811 47039
rect 2973 47005 3007 47039
rect 3801 47005 3835 47039
rect 6377 47005 6411 47039
rect 7113 47005 7147 47039
rect 7849 47005 7883 47039
rect 14105 47005 14139 47039
rect 16681 47005 16715 47039
rect 18153 47005 18187 47039
rect 19441 47005 19475 47039
rect 22017 47005 22051 47039
rect 26433 47005 26467 47039
rect 26985 47005 27019 47039
rect 28089 47005 28123 47039
rect 22201 46937 22235 46971
rect 26249 46937 26283 46971
rect 6561 46869 6595 46903
rect 7297 46869 7331 46903
rect 27077 46665 27111 46699
rect 23213 46597 23247 46631
rect 25605 46597 25639 46631
rect 1685 46529 1719 46563
rect 3985 46529 4019 46563
rect 7849 46529 7883 46563
rect 13829 46529 13863 46563
rect 16681 46529 16715 46563
rect 19441 46529 19475 46563
rect 26985 46529 27019 46563
rect 1869 46461 1903 46495
rect 2237 46461 2271 46495
rect 4169 46461 4203 46495
rect 4445 46461 4479 46495
rect 8033 46461 8067 46495
rect 8401 46461 8435 46495
rect 10977 46461 11011 46495
rect 11529 46461 11563 46495
rect 11713 46461 11747 46495
rect 11989 46461 12023 46495
rect 14013 46461 14047 46495
rect 14289 46461 14323 46495
rect 16865 46461 16899 46495
rect 17141 46461 17175 46495
rect 19625 46461 19659 46495
rect 19993 46461 20027 46495
rect 23765 46461 23799 46495
rect 23949 46461 23983 46495
rect 23029 46393 23063 46427
rect 10149 46325 10183 46359
rect 22109 46325 22143 46359
rect 26341 46325 26375 46359
rect 27905 46325 27939 46359
rect 2145 46121 2179 46155
rect 3157 46121 3191 46155
rect 8033 46121 8067 46155
rect 13461 46121 13495 46155
rect 16681 46121 16715 46155
rect 24409 46121 24443 46155
rect 3801 45985 3835 46019
rect 4261 45985 4295 46019
rect 9597 45985 9631 46019
rect 10149 45985 10183 46019
rect 19717 45985 19751 46019
rect 21281 45985 21315 46019
rect 22017 45985 22051 46019
rect 22569 45985 22603 46019
rect 26341 45985 26375 46019
rect 28181 45985 28215 46019
rect 1593 45917 1627 45951
rect 2237 45917 2271 45951
rect 3249 45917 3283 45951
rect 7941 45917 7975 45951
rect 13553 45917 13587 45951
rect 14289 45917 14323 45951
rect 16589 45917 16623 45951
rect 18245 45917 18279 45951
rect 25881 45917 25915 45951
rect 3985 45849 4019 45883
rect 9781 45849 9815 45883
rect 14473 45849 14507 45883
rect 16129 45849 16163 45883
rect 19901 45849 19935 45883
rect 22201 45849 22235 45883
rect 27997 45849 28031 45883
rect 18337 45781 18371 45815
rect 25789 45781 25823 45815
rect 9873 45577 9907 45611
rect 14473 45577 14507 45611
rect 20545 45577 20579 45611
rect 22109 45577 22143 45611
rect 4537 45509 4571 45543
rect 10701 45509 10735 45543
rect 18337 45509 18371 45543
rect 22753 45509 22787 45543
rect 23397 45509 23431 45543
rect 26249 45509 26283 45543
rect 27537 45509 27571 45543
rect 1593 45441 1627 45475
rect 4629 45441 4663 45475
rect 9965 45441 9999 45475
rect 10609 45441 10643 45475
rect 14381 45441 14415 45475
rect 18153 45441 18187 45475
rect 20453 45441 20487 45475
rect 22017 45441 22051 45475
rect 22845 45441 22879 45475
rect 23305 45441 23339 45475
rect 26433 45441 26467 45475
rect 27445 45441 27479 45475
rect 1777 45373 1811 45407
rect 2053 45373 2087 45407
rect 15025 45373 15059 45407
rect 18705 45373 18739 45407
rect 25973 45373 26007 45407
rect 1961 45033 1995 45067
rect 19533 45033 19567 45067
rect 20177 45033 20211 45067
rect 22661 45033 22695 45067
rect 12541 44897 12575 44931
rect 27537 44897 27571 44931
rect 28181 44897 28215 44931
rect 2053 44829 2087 44863
rect 10701 44829 10735 44863
rect 11161 44829 11195 44863
rect 19441 44829 19475 44863
rect 11345 44761 11379 44795
rect 27997 44761 28031 44795
rect 11621 44489 11655 44523
rect 27629 44489 27663 44523
rect 2329 44353 2363 44387
rect 11713 44353 11747 44387
rect 27537 44353 27571 44387
rect 1501 44149 1535 44183
rect 2237 44149 2271 44183
rect 2789 44149 2823 44183
rect 26433 44149 26467 44183
rect 1409 43809 1443 43843
rect 1593 43809 1627 43843
rect 2881 43809 2915 43843
rect 27997 43809 28031 43843
rect 25881 43741 25915 43775
rect 26341 43741 26375 43775
rect 26525 43673 26559 43707
rect 27077 43401 27111 43435
rect 2513 43265 2547 43299
rect 27169 43265 27203 43299
rect 27813 43265 27847 43299
rect 2697 43197 2731 43231
rect 3065 43197 3099 43231
rect 27721 43061 27755 43095
rect 2973 42721 3007 42755
rect 26341 42721 26375 42755
rect 26525 42721 26559 42755
rect 28181 42721 28215 42755
rect 1777 42653 1811 42687
rect 3065 42653 3099 42687
rect 27721 42177 27755 42211
rect 2789 42109 2823 42143
rect 4445 42109 4479 42143
rect 4629 42109 4663 42143
rect 1593 41973 1627 42007
rect 26433 41973 26467 42007
rect 27077 41973 27111 42007
rect 27813 41973 27847 42007
rect 3893 41769 3927 41803
rect 4629 41769 4663 41803
rect 1409 41633 1443 41667
rect 3249 41633 3283 41667
rect 26341 41633 26375 41667
rect 28181 41633 28215 41667
rect 3985 41565 4019 41599
rect 3065 41497 3099 41531
rect 26525 41497 26559 41531
rect 1593 41089 1627 41123
rect 26433 41089 26467 41123
rect 27169 41089 27203 41123
rect 1777 41021 1811 41055
rect 3249 41021 3283 41055
rect 25973 41021 26007 41055
rect 26249 41021 26283 41055
rect 27077 41021 27111 41055
rect 28089 40885 28123 40919
rect 2053 40681 2087 40715
rect 2697 40681 2731 40715
rect 27537 40545 27571 40579
rect 28181 40545 28215 40579
rect 2145 40477 2179 40511
rect 2789 40477 2823 40511
rect 27997 40409 28031 40443
rect 27813 40137 27847 40171
rect 27721 40001 27755 40035
rect 27077 39797 27111 39831
rect 21465 39525 21499 39559
rect 20729 39457 20763 39491
rect 26341 39457 26375 39491
rect 28181 39457 28215 39491
rect 20453 39389 20487 39423
rect 20545 39389 20579 39423
rect 21189 39389 21223 39423
rect 21465 39389 21499 39423
rect 26525 39321 26559 39355
rect 20729 39253 20763 39287
rect 21281 39253 21315 39287
rect 27629 39049 27663 39083
rect 19441 38913 19475 38947
rect 19625 38913 19659 38947
rect 20913 38913 20947 38947
rect 21833 38913 21867 38947
rect 22201 38913 22235 38947
rect 27721 38913 27755 38947
rect 20821 38845 20855 38879
rect 22109 38845 22143 38879
rect 20545 38777 20579 38811
rect 1685 38709 1719 38743
rect 19441 38709 19475 38743
rect 20821 38709 20855 38743
rect 21925 38709 21959 38743
rect 22293 38709 22327 38743
rect 26433 38709 26467 38743
rect 20637 38437 20671 38471
rect 1409 38369 1443 38403
rect 2789 38369 2823 38403
rect 21097 38369 21131 38403
rect 26341 38369 26375 38403
rect 28181 38369 28215 38403
rect 19257 38301 19291 38335
rect 19524 38301 19558 38335
rect 21373 38301 21407 38335
rect 23765 38301 23799 38335
rect 1593 38233 1627 38267
rect 23498 38233 23532 38267
rect 26525 38233 26559 38267
rect 22385 38165 22419 38199
rect 2145 37961 2179 37995
rect 19901 37961 19935 37995
rect 21081 37961 21115 37995
rect 22845 37961 22879 37995
rect 27721 37961 27755 37995
rect 21281 37893 21315 37927
rect 2237 37825 2271 37859
rect 20177 37825 20211 37859
rect 20269 37825 20303 37859
rect 22201 37825 22235 37859
rect 22385 37825 22419 37859
rect 22477 37825 22511 37859
rect 22569 37825 22603 37859
rect 27813 37825 27847 37859
rect 20085 37757 20119 37791
rect 20361 37757 20395 37791
rect 1593 37621 1627 37655
rect 20913 37621 20947 37655
rect 21097 37621 21131 37655
rect 19901 37417 19935 37451
rect 21373 37417 21407 37451
rect 27445 37281 27479 37315
rect 28089 37281 28123 37315
rect 1409 37213 1443 37247
rect 3249 37213 3283 37247
rect 20177 37213 20211 37247
rect 20913 37213 20947 37247
rect 21189 37213 21223 37247
rect 26801 37213 26835 37247
rect 3065 37145 3099 37179
rect 19901 37145 19935 37179
rect 21925 37145 21959 37179
rect 22109 37145 22143 37179
rect 20085 37077 20119 37111
rect 21005 37077 21039 37111
rect 26617 37077 26651 37111
rect 2789 36873 2823 36907
rect 1869 36737 1903 36771
rect 2697 36737 2731 36771
rect 17969 36737 18003 36771
rect 22661 36737 22695 36771
rect 27813 36737 27847 36771
rect 18245 36669 18279 36703
rect 2145 36533 2179 36567
rect 22569 36533 22603 36567
rect 27905 36533 27939 36567
rect 20085 36329 20119 36363
rect 27537 36193 27571 36227
rect 27997 36193 28031 36227
rect 28181 36193 28215 36227
rect 18061 36125 18095 36159
rect 20361 36125 20395 36159
rect 22017 36125 22051 36159
rect 22201 36125 22235 36159
rect 22661 36125 22695 36159
rect 22845 36125 22879 36159
rect 22937 36125 22971 36159
rect 23029 36125 23063 36159
rect 25237 36125 25271 36159
rect 18429 36057 18463 36091
rect 20085 36057 20119 36091
rect 20269 36057 20303 36091
rect 21005 36057 21039 36091
rect 22109 36057 22143 36091
rect 25421 36057 25455 36091
rect 20913 35989 20947 36023
rect 23305 35989 23339 36023
rect 20177 35785 20211 35819
rect 16957 35717 16991 35751
rect 18245 35717 18279 35751
rect 20821 35717 20855 35751
rect 24418 35717 24452 35751
rect 17141 35649 17175 35683
rect 17693 35649 17727 35683
rect 18797 35649 18831 35683
rect 19064 35649 19098 35683
rect 21065 35649 21099 35683
rect 21189 35649 21223 35683
rect 22477 35649 22511 35683
rect 25605 35649 25639 35683
rect 27629 35649 27663 35683
rect 21287 35581 21321 35615
rect 22385 35581 22419 35615
rect 24685 35581 24719 35615
rect 26157 35581 26191 35615
rect 1501 35445 1535 35479
rect 2329 35445 2363 35479
rect 22845 35445 22879 35479
rect 23305 35445 23339 35479
rect 26985 35445 27019 35479
rect 20637 35241 20671 35275
rect 22477 35241 22511 35275
rect 27261 35241 27295 35275
rect 22753 35173 22787 35207
rect 1409 35105 1443 35139
rect 2789 35105 2823 35139
rect 18337 35105 18371 35139
rect 20269 35105 20303 35139
rect 22845 35105 22879 35139
rect 25881 35105 25915 35139
rect 18061 35037 18095 35071
rect 19625 35037 19659 35071
rect 19809 35037 19843 35071
rect 20453 35037 20487 35071
rect 21465 35037 21499 35071
rect 22661 35037 22695 35071
rect 22937 35037 22971 35071
rect 23121 35037 23155 35071
rect 25329 35037 25363 35071
rect 26148 35037 26182 35071
rect 27721 35037 27755 35071
rect 1593 34969 1627 35003
rect 21281 34969 21315 35003
rect 24961 34969 24995 35003
rect 27997 34969 28031 35003
rect 19717 34901 19751 34935
rect 21097 34901 21131 34935
rect 1777 34629 1811 34663
rect 18613 34629 18647 34663
rect 21005 34629 21039 34663
rect 21123 34629 21157 34663
rect 27445 34629 27479 34663
rect 3617 34561 3651 34595
rect 18061 34561 18095 34595
rect 20821 34561 20855 34595
rect 20913 34561 20947 34595
rect 22017 34561 22051 34595
rect 22201 34561 22235 34595
rect 26177 34561 26211 34595
rect 26433 34561 26467 34595
rect 27077 34561 27111 34595
rect 3433 34493 3467 34527
rect 20637 34493 20671 34527
rect 21281 34493 21315 34527
rect 21833 34425 21867 34459
rect 22201 34357 22235 34391
rect 25053 34357 25087 34391
rect 2605 34153 2639 34187
rect 20177 34153 20211 34187
rect 21373 34153 21407 34187
rect 23489 34153 23523 34187
rect 23673 34153 23707 34187
rect 21281 34017 21315 34051
rect 21465 34017 21499 34051
rect 24409 34017 24443 34051
rect 27537 34017 27571 34051
rect 28181 34017 28215 34051
rect 2697 33949 2731 33983
rect 19257 33949 19291 33983
rect 19441 33949 19475 33983
rect 20361 33949 20395 33983
rect 20453 33949 20487 33983
rect 20729 33949 20763 33983
rect 21557 33949 21591 33983
rect 25789 33949 25823 33983
rect 20545 33881 20579 33915
rect 23857 33881 23891 33915
rect 24593 33881 24627 33915
rect 27997 33881 28031 33915
rect 19349 33813 19383 33847
rect 23657 33813 23691 33847
rect 25145 33813 25179 33847
rect 19349 33609 19383 33643
rect 24593 33609 24627 33643
rect 27169 33609 27203 33643
rect 22661 33541 22695 33575
rect 23480 33541 23514 33575
rect 27997 33541 28031 33575
rect 17969 33473 18003 33507
rect 18236 33473 18270 33507
rect 19809 33473 19843 33507
rect 20085 33473 20119 33507
rect 20177 33473 20211 33507
rect 27077 33473 27111 33507
rect 27721 33473 27755 33507
rect 23213 33405 23247 33439
rect 19901 33337 19935 33371
rect 20361 33269 20395 33303
rect 22569 33269 22603 33303
rect 25789 33269 25823 33303
rect 26433 33269 26467 33303
rect 19717 33065 19751 33099
rect 23029 33065 23063 33099
rect 19993 32997 20027 33031
rect 20085 32997 20119 33031
rect 23489 32997 23523 33031
rect 26341 32929 26375 32963
rect 28089 32929 28123 32963
rect 19901 32861 19935 32895
rect 20177 32861 20211 32895
rect 20361 32861 20395 32895
rect 22385 32861 22419 32895
rect 22569 32861 22603 32895
rect 22661 32861 22695 32895
rect 22753 32861 22787 32895
rect 23765 32861 23799 32895
rect 25881 32861 25915 32895
rect 23489 32793 23523 32827
rect 25789 32793 25823 32827
rect 26525 32793 26559 32827
rect 23673 32725 23707 32759
rect 20821 32521 20855 32555
rect 20361 32453 20395 32487
rect 26249 32453 26283 32487
rect 27813 32453 27847 32487
rect 16681 32385 16715 32419
rect 16937 32385 16971 32419
rect 19993 32385 20027 32419
rect 20177 32385 20211 32419
rect 21005 32385 21039 32419
rect 21189 32385 21223 32419
rect 22017 32385 22051 32419
rect 26985 32385 27019 32419
rect 27721 32385 27755 32419
rect 22109 32317 22143 32351
rect 25973 32317 26007 32351
rect 26433 32317 26467 32351
rect 1501 32181 1535 32215
rect 18061 32181 18095 32215
rect 22293 32181 22327 32215
rect 27077 32181 27111 32215
rect 22293 31977 22327 32011
rect 23489 31977 23523 32011
rect 16681 31909 16715 31943
rect 20269 31909 20303 31943
rect 1409 31841 1443 31875
rect 1869 31841 1903 31875
rect 17601 31841 17635 31875
rect 17785 31841 17819 31875
rect 22385 31841 22419 31875
rect 25605 31841 25639 31875
rect 27261 31841 27295 31875
rect 16497 31773 16531 31807
rect 18705 31773 18739 31807
rect 19257 31773 19291 31807
rect 19441 31773 19475 31807
rect 19625 31773 19659 31807
rect 20085 31773 20119 31807
rect 20269 31773 20303 31807
rect 21925 31773 21959 31807
rect 22109 31773 22143 31807
rect 22259 31773 22293 31807
rect 22477 31773 22511 31807
rect 23581 31773 23615 31807
rect 27445 31773 27479 31807
rect 28089 31773 28123 31807
rect 1593 31705 1627 31739
rect 17141 31637 17175 31671
rect 17509 31637 17543 31671
rect 18521 31637 18555 31671
rect 1869 31433 1903 31467
rect 16865 31433 16899 31467
rect 23949 31433 23983 31467
rect 17233 31365 17267 31399
rect 18512 31365 18546 31399
rect 1961 31297 1995 31331
rect 17049 31297 17083 31331
rect 21833 31297 21867 31331
rect 22017 31297 22051 31331
rect 22825 31297 22859 31331
rect 27813 31297 27847 31331
rect 18245 31229 18279 31263
rect 22569 31229 22603 31263
rect 19625 31093 19659 31127
rect 21833 31093 21867 31127
rect 27905 31093 27939 31127
rect 21281 30889 21315 30923
rect 20177 30821 20211 30855
rect 22017 30821 22051 30855
rect 27537 30753 27571 30787
rect 27997 30753 28031 30787
rect 28181 30753 28215 30787
rect 14841 30685 14875 30719
rect 15025 30685 15059 30719
rect 15669 30685 15703 30719
rect 17141 30685 17175 30719
rect 20453 30685 20487 30719
rect 20913 30685 20947 30719
rect 24961 30685 24995 30719
rect 25145 30685 25179 30719
rect 14657 30617 14691 30651
rect 17325 30617 17359 30651
rect 19257 30617 19291 30651
rect 19441 30617 19475 30651
rect 20177 30617 20211 30651
rect 20361 30617 20395 30651
rect 21097 30617 21131 30651
rect 21833 30617 21867 30651
rect 15485 30549 15519 30583
rect 16957 30549 16991 30583
rect 25053 30549 25087 30583
rect 17325 30345 17359 30379
rect 22477 30345 22511 30379
rect 14924 30277 14958 30311
rect 17693 30277 17727 30311
rect 23029 30277 23063 30311
rect 1409 30209 1443 30243
rect 16681 30209 16715 30243
rect 19257 30209 19291 30243
rect 19717 30209 19751 30243
rect 19809 30209 19843 30243
rect 19993 30209 20027 30243
rect 20683 30209 20717 30243
rect 20818 30209 20852 30243
rect 20913 30209 20947 30243
rect 21097 30209 21131 30243
rect 21833 30209 21867 30243
rect 22017 30209 22051 30243
rect 22109 30209 22143 30243
rect 22201 30209 22235 30243
rect 25136 30209 25170 30243
rect 27169 30209 27203 30243
rect 27997 30209 28031 30243
rect 14657 30141 14691 30175
rect 17785 30141 17819 30175
rect 17877 30141 17911 30175
rect 18981 30141 19015 30175
rect 24869 30141 24903 30175
rect 19165 30073 19199 30107
rect 20453 30073 20487 30107
rect 23213 30073 23247 30107
rect 1593 30005 1627 30039
rect 16037 30005 16071 30039
rect 16865 30005 16899 30039
rect 19257 30005 19291 30039
rect 19993 30005 20027 30039
rect 26249 30005 26283 30039
rect 27077 30005 27111 30039
rect 27905 30005 27939 30039
rect 14749 29801 14783 29835
rect 16129 29801 16163 29835
rect 21649 29801 21683 29835
rect 22109 29801 22143 29835
rect 15209 29665 15243 29699
rect 15301 29665 15335 29699
rect 21833 29665 21867 29699
rect 26525 29665 26559 29699
rect 28181 29665 28215 29699
rect 15945 29597 15979 29631
rect 16865 29597 16899 29631
rect 17132 29597 17166 29631
rect 19257 29597 19291 29631
rect 19513 29597 19547 29631
rect 21557 29597 21591 29631
rect 22569 29597 22603 29631
rect 22753 29597 22787 29631
rect 23213 29597 23247 29631
rect 23397 29597 23431 29631
rect 23489 29597 23523 29631
rect 23581 29597 23615 29631
rect 25789 29597 25823 29631
rect 26341 29597 26375 29631
rect 22661 29529 22695 29563
rect 23857 29529 23891 29563
rect 25522 29529 25556 29563
rect 15117 29461 15151 29495
rect 18245 29461 18279 29495
rect 20637 29461 20671 29495
rect 24409 29461 24443 29495
rect 27169 29257 27203 29291
rect 27353 29121 27387 29155
rect 27997 28917 28031 28951
rect 21833 28713 21867 28747
rect 23581 28713 23615 28747
rect 17693 28645 17727 28679
rect 27537 28577 27571 28611
rect 28181 28577 28215 28611
rect 21741 28509 21775 28543
rect 22477 28509 22511 28543
rect 22661 28509 22695 28543
rect 23121 28509 23155 28543
rect 23397 28509 23431 28543
rect 14197 28441 14231 28475
rect 14381 28441 14415 28475
rect 17325 28441 17359 28475
rect 27997 28441 28031 28475
rect 14565 28373 14599 28407
rect 17785 28373 17819 28407
rect 22569 28373 22603 28407
rect 23213 28373 23247 28407
rect 16129 28169 16163 28203
rect 20729 28169 20763 28203
rect 22109 28169 22143 28203
rect 25513 28169 25547 28203
rect 27353 28169 27387 28203
rect 15761 28101 15795 28135
rect 15961 28101 15995 28135
rect 23673 28101 23707 28135
rect 24378 28101 24412 28135
rect 1409 28033 1443 28067
rect 13636 28033 13670 28067
rect 16865 28033 16899 28067
rect 18337 28033 18371 28067
rect 18521 28033 18555 28067
rect 18613 28033 18647 28067
rect 19441 28033 19475 28067
rect 19717 28033 19751 28067
rect 20177 28033 20211 28067
rect 20545 28033 20579 28067
rect 20637 28033 20671 28067
rect 22385 28033 22419 28067
rect 23029 28033 23063 28067
rect 23213 28033 23247 28067
rect 23305 28033 23339 28067
rect 23397 28033 23431 28067
rect 27261 28033 27295 28067
rect 13369 27965 13403 27999
rect 17417 27965 17451 27999
rect 19625 27965 19659 27999
rect 22109 27965 22143 27999
rect 24133 27965 24167 27999
rect 17693 27897 17727 27931
rect 1593 27829 1627 27863
rect 14749 27829 14783 27863
rect 15945 27829 15979 27863
rect 16681 27829 16715 27863
rect 17877 27829 17911 27863
rect 18337 27829 18371 27863
rect 18797 27829 18831 27863
rect 19257 27829 19291 27863
rect 22293 27829 22327 27863
rect 28089 27829 28123 27863
rect 13553 27625 13587 27659
rect 14197 27625 14231 27659
rect 23029 27625 23063 27659
rect 17049 27557 17083 27591
rect 21649 27557 21683 27591
rect 22385 27557 22419 27591
rect 14657 27489 14691 27523
rect 14749 27489 14783 27523
rect 17509 27489 17543 27523
rect 17785 27489 17819 27523
rect 19717 27489 19751 27523
rect 20269 27489 20303 27523
rect 20821 27489 20855 27523
rect 27537 27489 27571 27523
rect 28181 27489 28215 27523
rect 13369 27421 13403 27455
rect 15669 27421 15703 27455
rect 15936 27421 15970 27455
rect 19809 27421 19843 27455
rect 20453 27421 20487 27455
rect 22201 27421 22235 27455
rect 23213 27421 23247 27455
rect 23489 27421 23523 27455
rect 21281 27353 21315 27387
rect 21465 27353 21499 27387
rect 27997 27353 28031 27387
rect 14565 27285 14599 27319
rect 20729 27285 20763 27319
rect 23397 27285 23431 27319
rect 15761 27081 15795 27115
rect 16773 27081 16807 27115
rect 20269 27081 20303 27115
rect 27721 27081 27755 27115
rect 20821 27013 20855 27047
rect 21005 27013 21039 27047
rect 15945 26945 15979 26979
rect 16129 26945 16163 26979
rect 16681 26945 16715 26979
rect 16865 26945 16899 26979
rect 17325 26945 17359 26979
rect 18245 26945 18279 26979
rect 18429 26945 18463 26979
rect 18889 26945 18923 26979
rect 19156 26945 19190 26979
rect 22109 26945 22143 26979
rect 22753 26945 22787 26979
rect 22937 26945 22971 26979
rect 27629 26945 27663 26979
rect 17785 26877 17819 26911
rect 21833 26877 21867 26911
rect 22017 26877 22051 26911
rect 17601 26809 17635 26843
rect 18245 26741 18279 26775
rect 21925 26741 21959 26775
rect 22937 26741 22971 26775
rect 17969 26537 18003 26571
rect 17785 26469 17819 26503
rect 19257 26469 19291 26503
rect 21833 26469 21867 26503
rect 17509 26401 17543 26435
rect 21557 26401 21591 26435
rect 14749 26333 14783 26367
rect 15577 26333 15611 26367
rect 15853 26333 15887 26367
rect 19257 26333 19291 26367
rect 19441 26333 19475 26367
rect 19533 26333 19567 26367
rect 19993 26333 20027 26367
rect 21373 26333 21407 26367
rect 21465 26333 21499 26367
rect 21649 26333 21683 26367
rect 22293 26333 22327 26367
rect 22477 26333 22511 26367
rect 22753 26333 22787 26367
rect 23213 26333 23247 26367
rect 23305 26333 23339 26367
rect 23489 26333 23523 26367
rect 24409 26333 24443 26367
rect 27261 26333 27295 26367
rect 28089 26333 28123 26367
rect 15761 26265 15795 26299
rect 20085 26265 20119 26299
rect 22661 26265 22695 26299
rect 24654 26265 24688 26299
rect 14565 26197 14599 26231
rect 15393 26197 15427 26231
rect 23673 26197 23707 26231
rect 25789 26197 25823 26231
rect 15393 25993 15427 26027
rect 19165 25993 19199 26027
rect 22661 25993 22695 26027
rect 14280 25925 14314 25959
rect 24501 25925 24535 25959
rect 12541 25857 12575 25891
rect 12725 25857 12759 25891
rect 12909 25857 12943 25891
rect 13553 25857 13587 25891
rect 17785 25857 17819 25891
rect 17877 25857 17911 25891
rect 18153 25857 18187 25891
rect 19073 25857 19107 25891
rect 19257 25857 19291 25891
rect 22477 25857 22511 25891
rect 23121 25857 23155 25891
rect 23305 25857 23339 25891
rect 23397 25857 23431 25891
rect 23535 25857 23569 25891
rect 24225 25857 24259 25891
rect 24317 25857 24351 25891
rect 25145 25857 25179 25891
rect 27537 25857 27571 25891
rect 14013 25789 14047 25823
rect 18061 25789 18095 25823
rect 22293 25789 22327 25823
rect 24501 25721 24535 25755
rect 25053 25721 25087 25755
rect 1501 25653 1535 25687
rect 13369 25653 13403 25687
rect 17601 25653 17635 25687
rect 23765 25653 23799 25687
rect 27629 25653 27663 25687
rect 14933 25449 14967 25483
rect 15117 25449 15151 25483
rect 22201 25449 22235 25483
rect 22661 25449 22695 25483
rect 23765 25449 23799 25483
rect 16497 25381 16531 25415
rect 1409 25313 1443 25347
rect 2789 25313 2823 25347
rect 13553 25313 13587 25347
rect 22845 25313 22879 25347
rect 22937 25313 22971 25347
rect 23121 25313 23155 25347
rect 27537 25313 27571 25347
rect 27997 25313 28031 25347
rect 28181 25313 28215 25347
rect 5549 25245 5583 25279
rect 13286 25245 13320 25279
rect 16313 25245 16347 25279
rect 21925 25245 21959 25279
rect 22017 25245 22051 25279
rect 23029 25245 23063 25279
rect 23673 25245 23707 25279
rect 23857 25245 23891 25279
rect 25789 25245 25823 25279
rect 1593 25177 1627 25211
rect 4997 25177 5031 25211
rect 15301 25177 15335 25211
rect 16129 25177 16163 25211
rect 22201 25177 22235 25211
rect 25522 25177 25556 25211
rect 12173 25109 12207 25143
rect 15101 25109 15135 25143
rect 15945 25109 15979 25143
rect 16221 25109 16255 25143
rect 24409 25109 24443 25143
rect 1777 24905 1811 24939
rect 12725 24905 12759 24939
rect 15301 24905 15335 24939
rect 17785 24905 17819 24939
rect 13093 24837 13127 24871
rect 1869 24769 1903 24803
rect 4353 24769 4387 24803
rect 4997 24769 5031 24803
rect 6377 24769 6411 24803
rect 15301 24769 15335 24803
rect 15485 24769 15519 24803
rect 16681 24769 16715 24803
rect 17601 24769 17635 24803
rect 17693 24769 17727 24803
rect 18889 24769 18923 24803
rect 21281 24769 21315 24803
rect 26433 24769 26467 24803
rect 26985 24769 27019 24803
rect 27721 24769 27755 24803
rect 4077 24701 4111 24735
rect 5181 24701 5215 24735
rect 6561 24701 6595 24735
rect 13185 24701 13219 24735
rect 13369 24701 13403 24735
rect 18061 24701 18095 24735
rect 21833 24701 21867 24735
rect 22109 24701 22143 24735
rect 25973 24701 26007 24735
rect 26249 24701 26283 24735
rect 27813 24701 27847 24735
rect 16773 24565 16807 24599
rect 17141 24565 17175 24599
rect 18981 24565 19015 24599
rect 19993 24565 20027 24599
rect 27169 24565 27203 24599
rect 15945 24361 15979 24395
rect 16681 24361 16715 24395
rect 19441 24361 19475 24395
rect 22293 24361 22327 24395
rect 18613 24225 18647 24259
rect 20821 24225 20855 24259
rect 27537 24225 27571 24259
rect 1409 24157 1443 24191
rect 4997 24157 5031 24191
rect 12173 24157 12207 24191
rect 15301 24157 15335 24191
rect 16589 24157 16623 24191
rect 18337 24157 18371 24191
rect 21281 24157 21315 24191
rect 25881 24157 25915 24191
rect 28181 24157 28215 24191
rect 5457 24089 5491 24123
rect 16129 24089 16163 24123
rect 20554 24089 20588 24123
rect 22385 24089 22419 24123
rect 25053 24089 25087 24123
rect 27997 24089 28031 24123
rect 1593 24021 1627 24055
rect 12357 24021 12391 24055
rect 15117 24021 15151 24055
rect 15761 24021 15795 24055
rect 15929 24021 15963 24055
rect 17049 24021 17083 24055
rect 21465 24021 21499 24055
rect 17601 23817 17635 23851
rect 18521 23817 18555 23851
rect 27721 23817 27755 23851
rect 4905 23749 4939 23783
rect 15016 23749 15050 23783
rect 21833 23749 21867 23783
rect 22033 23749 22067 23783
rect 22845 23749 22879 23783
rect 27445 23749 27479 23783
rect 4721 23681 4755 23715
rect 12633 23681 12667 23715
rect 17141 23681 17175 23715
rect 19645 23681 19679 23715
rect 20821 23681 20855 23715
rect 21189 23681 21223 23715
rect 25605 23681 25639 23715
rect 12725 23613 12759 23647
rect 12909 23613 12943 23647
rect 14749 23613 14783 23647
rect 19901 23613 19935 23647
rect 26157 23613 26191 23647
rect 22661 23545 22695 23579
rect 12265 23477 12299 23511
rect 16129 23477 16163 23511
rect 17233 23477 17267 23511
rect 20637 23477 20671 23511
rect 21097 23477 21131 23511
rect 22017 23477 22051 23511
rect 22201 23477 22235 23511
rect 13553 23273 13587 23307
rect 15393 23273 15427 23307
rect 15577 23273 15611 23307
rect 17509 23273 17543 23307
rect 19901 23273 19935 23307
rect 20821 23273 20855 23307
rect 21649 23273 21683 23307
rect 27997 23273 28031 23307
rect 15945 23205 15979 23239
rect 18429 23205 18463 23239
rect 23121 23205 23155 23239
rect 24869 23205 24903 23239
rect 22293 23137 22327 23171
rect 23673 23137 23707 23171
rect 12173 23069 12207 23103
rect 12440 23069 12474 23103
rect 16589 23069 16623 23103
rect 16865 23069 16899 23103
rect 18153 23069 18187 23103
rect 18245 23069 18279 23103
rect 19257 23069 19291 23103
rect 19441 23069 19475 23103
rect 19533 23069 19567 23103
rect 19625 23069 19659 23103
rect 22477 23069 22511 23103
rect 24593 23069 24627 23103
rect 24685 23069 24719 23103
rect 24869 23069 24903 23103
rect 25605 23069 25639 23103
rect 26065 23069 26099 23103
rect 26893 23069 26927 23103
rect 27905 23069 27939 23103
rect 16773 23001 16807 23035
rect 17325 23001 17359 23035
rect 17525 23001 17559 23035
rect 18429 23001 18463 23035
rect 20637 23001 20671 23035
rect 20853 23001 20887 23035
rect 21465 23001 21499 23035
rect 21681 23001 21715 23035
rect 23581 23001 23615 23035
rect 15577 22933 15611 22967
rect 16405 22933 16439 22967
rect 17693 22933 17727 22967
rect 21005 22933 21039 22967
rect 21833 22933 21867 22967
rect 22661 22933 22695 22967
rect 23489 22933 23523 22967
rect 25421 22933 25455 22967
rect 12909 22729 12943 22763
rect 18981 22729 19015 22763
rect 20269 22729 20303 22763
rect 24225 22729 24259 22763
rect 12541 22661 12575 22695
rect 12725 22661 12759 22695
rect 21833 22661 21867 22695
rect 22033 22661 22067 22695
rect 14482 22593 14516 22627
rect 14749 22593 14783 22627
rect 18889 22593 18923 22627
rect 19073 22593 19107 22627
rect 20085 22593 20119 22627
rect 22845 22593 22879 22627
rect 23101 22593 23135 22627
rect 24961 22593 24995 22627
rect 25217 22593 25251 22627
rect 27169 22593 27203 22627
rect 27721 22593 27755 22627
rect 27813 22457 27847 22491
rect 13369 22389 13403 22423
rect 22017 22389 22051 22423
rect 22201 22389 22235 22423
rect 26341 22389 26375 22423
rect 27077 22389 27111 22423
rect 14289 22185 14323 22219
rect 22937 22185 22971 22219
rect 25053 22185 25087 22219
rect 23857 22117 23891 22151
rect 25421 22049 25455 22083
rect 26525 22049 26559 22083
rect 28181 22049 28215 22083
rect 1593 21981 1627 22015
rect 14105 21981 14139 22015
rect 19993 21981 20027 22015
rect 21005 21981 21039 22015
rect 22753 21981 22787 22015
rect 24593 21981 24627 22015
rect 25237 21981 25271 22015
rect 25513 21981 25547 22015
rect 26341 21981 26375 22015
rect 24501 21913 24535 21947
rect 19809 21845 19843 21879
rect 20821 21845 20855 21879
rect 17233 21641 17267 21675
rect 18061 21641 18095 21675
rect 18245 21641 18279 21675
rect 19717 21641 19751 21675
rect 15485 21573 15519 21607
rect 17877 21573 17911 21607
rect 19073 21573 19107 21607
rect 20637 21573 20671 21607
rect 24777 21573 24811 21607
rect 2145 21505 2179 21539
rect 15301 21505 15335 21539
rect 15577 21505 15611 21539
rect 17325 21505 17359 21539
rect 18153 21505 18187 21539
rect 19901 21505 19935 21539
rect 20361 21505 20395 21539
rect 20453 21505 20487 21539
rect 21097 21505 21131 21539
rect 21281 21505 21315 21539
rect 22017 21505 22051 21539
rect 22201 21505 22235 21539
rect 27721 21505 27755 21539
rect 22293 21437 22327 21471
rect 24133 21437 24167 21471
rect 24593 21437 24627 21471
rect 26157 21437 26191 21471
rect 20637 21369 20671 21403
rect 2053 21301 2087 21335
rect 15117 21301 15151 21335
rect 18429 21301 18463 21335
rect 18981 21301 19015 21335
rect 21097 21301 21131 21335
rect 21833 21301 21867 21335
rect 27629 21301 27663 21335
rect 15025 21097 15059 21131
rect 17049 21097 17083 21131
rect 19257 21097 19291 21131
rect 14841 21029 14875 21063
rect 1409 20961 1443 20995
rect 25237 20961 25271 20995
rect 25329 20961 25363 20995
rect 26341 20961 26375 20995
rect 26525 20961 26559 20995
rect 28181 20961 28215 20995
rect 12449 20893 12483 20927
rect 13093 20893 13127 20927
rect 14289 20893 14323 20927
rect 15669 20893 15703 20927
rect 15853 20893 15887 20927
rect 16957 20893 16991 20927
rect 17933 20893 17967 20927
rect 18061 20893 18095 20927
rect 18153 20893 18187 20927
rect 19441 20893 19475 20927
rect 19533 20893 19567 20927
rect 19717 20893 19751 20927
rect 19809 20893 19843 20927
rect 21005 20893 21039 20927
rect 21465 20893 21499 20927
rect 21732 20893 21766 20927
rect 23305 20893 23339 20927
rect 1593 20825 1627 20859
rect 3249 20825 3283 20859
rect 12081 20825 12115 20859
rect 12265 20825 12299 20859
rect 15209 20825 15243 20859
rect 18337 20825 18371 20859
rect 12909 20757 12943 20791
rect 14105 20757 14139 20791
rect 14999 20757 15033 20791
rect 15669 20757 15703 20791
rect 20821 20757 20855 20791
rect 22845 20757 22879 20791
rect 23489 20757 23523 20791
rect 24777 20757 24811 20791
rect 25145 20757 25179 20791
rect 18337 20553 18371 20587
rect 18705 20553 18739 20587
rect 21097 20553 21131 20587
rect 22569 20553 22603 20587
rect 25881 20553 25915 20587
rect 14096 20485 14130 20519
rect 15669 20485 15703 20519
rect 17233 20485 17267 20519
rect 19984 20485 20018 20519
rect 23756 20485 23790 20519
rect 15899 20451 15933 20485
rect 12256 20417 12290 20451
rect 13829 20417 13863 20451
rect 18521 20417 18555 20451
rect 18797 20417 18831 20451
rect 22661 20417 22695 20451
rect 23489 20417 23523 20451
rect 25789 20417 25823 20451
rect 27353 20417 27387 20451
rect 28089 20417 28123 20451
rect 2329 20349 2363 20383
rect 2513 20349 2547 20383
rect 2973 20349 3007 20383
rect 11989 20349 12023 20383
rect 19717 20349 19751 20383
rect 22477 20349 22511 20383
rect 25973 20349 26007 20383
rect 13369 20213 13403 20247
rect 15209 20213 15243 20247
rect 15853 20213 15887 20247
rect 16037 20213 16071 20247
rect 17141 20213 17175 20247
rect 23029 20213 23063 20247
rect 24869 20213 24903 20247
rect 25421 20213 25455 20247
rect 27261 20213 27295 20247
rect 2329 20009 2363 20043
rect 2881 20009 2915 20043
rect 12265 20009 12299 20043
rect 14841 20009 14875 20043
rect 15025 20009 15059 20043
rect 18337 20009 18371 20043
rect 21373 20009 21407 20043
rect 22293 20009 22327 20043
rect 23581 20009 23615 20043
rect 25881 20009 25915 20043
rect 16773 19941 16807 19975
rect 12817 19873 12851 19907
rect 20637 19873 20671 19907
rect 22477 19873 22511 19907
rect 24501 19873 24535 19907
rect 26525 19873 26559 19907
rect 28181 19873 28215 19907
rect 1501 19805 1535 19839
rect 2973 19805 3007 19839
rect 14197 19805 14231 19839
rect 14381 19805 14415 19839
rect 15669 19805 15703 19839
rect 15761 19805 15795 19839
rect 15945 19805 15979 19839
rect 16957 19805 16991 19839
rect 17581 19805 17615 19839
rect 17785 19805 17819 19839
rect 18429 19805 18463 19839
rect 20269 19805 20303 19839
rect 21281 19805 21315 19839
rect 22017 19805 22051 19839
rect 23213 19805 23247 19839
rect 23397 19805 23431 19839
rect 26341 19805 26375 19839
rect 12633 19737 12667 19771
rect 14289 19737 14323 19771
rect 14993 19737 15027 19771
rect 15209 19737 15243 19771
rect 17499 19737 17533 19771
rect 17693 19737 17727 19771
rect 20453 19737 20487 19771
rect 22109 19737 22143 19771
rect 24768 19737 24802 19771
rect 12725 19669 12759 19703
rect 15669 19669 15703 19703
rect 25145 19465 25179 19499
rect 16957 19397 16991 19431
rect 17173 19397 17207 19431
rect 17969 19397 18003 19431
rect 20637 19397 20671 19431
rect 1409 19329 1443 19363
rect 14841 19329 14875 19363
rect 14933 19329 14967 19363
rect 24501 19329 24535 19363
rect 24685 19329 24719 19363
rect 25329 19329 25363 19363
rect 26433 19329 26467 19363
rect 1593 19261 1627 19295
rect 1869 19261 1903 19295
rect 24317 19261 24351 19295
rect 17141 19125 17175 19159
rect 17325 19125 17359 19159
rect 17877 19125 17911 19159
rect 20545 19125 20579 19159
rect 27445 19125 27479 19159
rect 28089 19125 28123 19159
rect 1869 18921 1903 18955
rect 17509 18921 17543 18955
rect 22017 18921 22051 18955
rect 17141 18785 17175 18819
rect 21373 18785 21407 18819
rect 27353 18785 27387 18819
rect 28181 18785 28215 18819
rect 1961 18717 1995 18751
rect 2421 18717 2455 18751
rect 16497 18717 16531 18751
rect 18153 18717 18187 18751
rect 21189 18717 21223 18751
rect 21925 18717 21959 18751
rect 22201 18717 22235 18751
rect 16313 18649 16347 18683
rect 27997 18649 28031 18683
rect 2605 18581 2639 18615
rect 16681 18581 16715 18615
rect 17509 18581 17543 18615
rect 17693 18581 17727 18615
rect 18337 18581 18371 18615
rect 22385 18581 22419 18615
rect 16681 18377 16715 18411
rect 22937 18377 22971 18411
rect 25329 18377 25363 18411
rect 27813 18377 27847 18411
rect 18328 18309 18362 18343
rect 22845 18309 22879 18343
rect 12357 18241 12391 18275
rect 12449 18241 12483 18275
rect 13277 18241 13311 18275
rect 14381 18241 14415 18275
rect 14657 18241 14691 18275
rect 14841 18241 14875 18275
rect 16865 18241 16899 18275
rect 16957 18241 16991 18275
rect 18061 18241 18095 18275
rect 20821 18241 20855 18275
rect 21005 18241 21039 18275
rect 22017 18241 22051 18275
rect 22201 18241 22235 18275
rect 22753 18241 22787 18275
rect 23857 18241 23891 18275
rect 25421 18241 25455 18275
rect 27169 18241 27203 18275
rect 27721 18241 27755 18275
rect 14473 18173 14507 18207
rect 21097 18173 21131 18207
rect 22293 18173 22327 18207
rect 23213 18173 23247 18207
rect 24041 18173 24075 18207
rect 25145 18173 25179 18207
rect 14565 18105 14599 18139
rect 1409 18037 1443 18071
rect 12173 18037 12207 18071
rect 13369 18037 13403 18071
rect 13737 18037 13771 18071
rect 14197 18037 14231 18071
rect 19441 18037 19475 18071
rect 20637 18037 20671 18071
rect 21833 18037 21867 18071
rect 23673 18037 23707 18071
rect 25789 18037 25823 18071
rect 27077 18037 27111 18071
rect 16129 17833 16163 17867
rect 18613 17833 18647 17867
rect 23397 17833 23431 17867
rect 16497 17765 16531 17799
rect 1409 17697 1443 17731
rect 2789 17697 2823 17731
rect 14473 17697 14507 17731
rect 22017 17697 22051 17731
rect 26525 17697 26559 17731
rect 26801 17697 26835 17731
rect 11253 17629 11287 17663
rect 11897 17629 11931 17663
rect 14105 17629 14139 17663
rect 14381 17629 14415 17663
rect 14565 17629 14599 17663
rect 16957 17629 16991 17663
rect 18337 17629 18371 17663
rect 19809 17629 19843 17663
rect 24409 17629 24443 17663
rect 26341 17629 26375 17663
rect 1593 17561 1627 17595
rect 12142 17561 12176 17595
rect 18613 17561 18647 17595
rect 20076 17561 20110 17595
rect 22284 17561 22318 17595
rect 24654 17561 24688 17595
rect 11437 17493 11471 17527
rect 13277 17493 13311 17527
rect 14197 17493 14231 17527
rect 14841 17493 14875 17527
rect 15945 17493 15979 17527
rect 16129 17493 16163 17527
rect 17141 17493 17175 17527
rect 18429 17493 18463 17527
rect 21189 17493 21223 17527
rect 25789 17493 25823 17527
rect 1685 17289 1719 17323
rect 12265 17289 12299 17323
rect 12633 17289 12667 17323
rect 13921 17289 13955 17323
rect 14657 17289 14691 17323
rect 15485 17289 15519 17323
rect 21005 17289 21039 17323
rect 21925 17289 21959 17323
rect 23489 17289 23523 17323
rect 27537 17289 27571 17323
rect 13461 17221 13495 17255
rect 14866 17221 14900 17255
rect 17049 17221 17083 17255
rect 23949 17221 23983 17255
rect 26157 17221 26191 17255
rect 1777 17153 1811 17187
rect 14381 17153 14415 17187
rect 14749 17153 14783 17187
rect 16681 17153 16715 17187
rect 16865 17153 16899 17187
rect 20177 17153 20211 17187
rect 20821 17153 20855 17187
rect 20913 17153 20947 17187
rect 21833 17153 21867 17187
rect 22109 17153 22143 17187
rect 23857 17153 23891 17187
rect 25697 17153 25731 17187
rect 25789 17153 25823 17187
rect 25973 17153 26007 17187
rect 26985 17153 27019 17187
rect 27077 17153 27111 17187
rect 27261 17153 27295 17187
rect 27353 17153 27387 17187
rect 27997 17153 28031 17187
rect 12725 17085 12759 17119
rect 12909 17085 12943 17119
rect 15945 17085 15979 17119
rect 21281 17085 21315 17119
rect 22293 17085 22327 17119
rect 24041 17085 24075 17119
rect 13737 17017 13771 17051
rect 15577 17017 15611 17051
rect 15025 16949 15059 16983
rect 20269 16949 20303 16983
rect 28089 16949 28123 16983
rect 14657 16745 14691 16779
rect 15761 16745 15795 16779
rect 18061 16745 18095 16779
rect 18245 16745 18279 16779
rect 23765 16745 23799 16779
rect 20545 16677 20579 16711
rect 25605 16677 25639 16711
rect 14197 16609 14231 16643
rect 15301 16609 15335 16643
rect 15485 16609 15519 16643
rect 17601 16609 17635 16643
rect 21005 16609 21039 16643
rect 27997 16609 28031 16643
rect 28181 16609 28215 16643
rect 14105 16541 14139 16575
rect 14381 16541 14415 16575
rect 14473 16541 14507 16575
rect 15393 16541 15427 16575
rect 15577 16541 15611 16575
rect 17334 16541 17368 16575
rect 19257 16541 19291 16575
rect 20361 16541 20395 16575
rect 21189 16541 21223 16575
rect 23581 16541 23615 16575
rect 25053 16541 25087 16575
rect 25513 16541 25547 16575
rect 25697 16541 25731 16575
rect 26341 16541 26375 16575
rect 18213 16473 18247 16507
rect 18429 16473 18463 16507
rect 24961 16473 24995 16507
rect 16221 16405 16255 16439
rect 19349 16405 19383 16439
rect 12817 16201 12851 16235
rect 15669 16201 15703 16235
rect 18061 16201 18095 16235
rect 19809 16201 19843 16235
rect 18429 16133 18463 16167
rect 26985 16133 27019 16167
rect 28089 16133 28123 16167
rect 12725 16065 12759 16099
rect 15485 16065 15519 16099
rect 17141 16065 17175 16099
rect 19165 16065 19199 16099
rect 19349 16065 19383 16099
rect 19441 16065 19475 16099
rect 19533 16065 19567 16099
rect 25697 16065 25731 16099
rect 25789 16065 25823 16099
rect 25973 16065 26007 16099
rect 26065 16065 26099 16099
rect 27261 16065 27295 16099
rect 13001 15997 13035 16031
rect 15301 15997 15335 16031
rect 17601 15997 17635 16031
rect 18220 15997 18254 16031
rect 18337 15997 18371 16031
rect 18705 15997 18739 16031
rect 25053 15997 25087 16031
rect 26985 15997 27019 16031
rect 2697 15861 2731 15895
rect 12357 15861 12391 15895
rect 17417 15861 17451 15895
rect 25513 15861 25547 15895
rect 27169 15861 27203 15895
rect 27997 15861 28031 15895
rect 15117 15657 15151 15691
rect 17969 15657 18003 15691
rect 19257 15657 19291 15691
rect 19717 15657 19751 15691
rect 20729 15657 20763 15691
rect 25237 15657 25271 15691
rect 14197 15589 14231 15623
rect 17417 15589 17451 15623
rect 11989 15521 12023 15555
rect 14105 15521 14139 15555
rect 17049 15521 17083 15555
rect 17509 15521 17543 15555
rect 18245 15521 18279 15555
rect 22661 15521 22695 15555
rect 22845 15521 22879 15555
rect 25881 15521 25915 15555
rect 26341 15521 26375 15555
rect 28181 15521 28215 15555
rect 1501 15453 1535 15487
rect 3985 15453 4019 15487
rect 12173 15453 12207 15487
rect 12357 15453 12391 15487
rect 13001 15453 13035 15487
rect 15025 15453 15059 15487
rect 15669 15453 15703 15487
rect 15853 15453 15887 15487
rect 18337 15453 18371 15487
rect 18429 15453 18463 15487
rect 18705 15453 18739 15487
rect 19441 15453 19475 15487
rect 19533 15453 19567 15487
rect 19809 15453 19843 15487
rect 20269 15453 20303 15487
rect 20545 15453 20579 15487
rect 24777 15453 24811 15487
rect 25421 15453 25455 15487
rect 14565 15385 14599 15419
rect 20361 15385 20395 15419
rect 22937 15385 22971 15419
rect 25513 15385 25547 15419
rect 25605 15385 25639 15419
rect 25743 15385 25777 15419
rect 26525 15385 26559 15419
rect 3893 15317 3927 15351
rect 12817 15317 12851 15351
rect 15669 15317 15703 15351
rect 18613 15317 18647 15351
rect 23305 15317 23339 15351
rect 24593 15317 24627 15351
rect 13369 15113 13403 15147
rect 18889 15113 18923 15147
rect 20637 15113 20671 15147
rect 24133 15113 24167 15147
rect 26341 15113 26375 15147
rect 28089 15113 28123 15147
rect 4169 15045 4203 15079
rect 12256 15045 12290 15079
rect 19349 15045 19383 15079
rect 22998 15045 23032 15079
rect 1961 14977 1995 15011
rect 4353 14977 4387 15011
rect 11989 14977 12023 15011
rect 15025 14977 15059 15011
rect 15209 14977 15243 15011
rect 20545 14977 20579 15011
rect 22109 14977 22143 15011
rect 26249 14977 26283 15011
rect 26433 14977 26467 15011
rect 27353 14977 27387 15011
rect 27997 14977 28031 15011
rect 2789 14909 2823 14943
rect 20729 14909 20763 14943
rect 22753 14909 22787 14943
rect 24961 14909 24995 14943
rect 25237 14909 25271 14943
rect 27169 14909 27203 14943
rect 27261 14909 27295 14943
rect 27445 14909 27479 14943
rect 19073 14841 19107 14875
rect 22293 14841 22327 14875
rect 1869 14773 1903 14807
rect 15117 14773 15151 14807
rect 20177 14773 20211 14807
rect 26985 14773 27019 14807
rect 15301 14569 15335 14603
rect 16037 14569 16071 14603
rect 22845 14569 22879 14603
rect 25145 14569 25179 14603
rect 25881 14569 25915 14603
rect 22385 14501 22419 14535
rect 1409 14433 1443 14467
rect 1593 14433 1627 14467
rect 1869 14433 1903 14467
rect 19809 14433 19843 14467
rect 24501 14433 24535 14467
rect 24685 14433 24719 14467
rect 27537 14433 27571 14467
rect 15945 14365 15979 14399
rect 19993 14365 20027 14399
rect 21005 14365 21039 14399
rect 23029 14365 23063 14399
rect 23213 14365 23247 14399
rect 24777 14365 24811 14399
rect 25605 14365 25639 14399
rect 25881 14365 25915 14399
rect 28181 14365 28215 14399
rect 15269 14297 15303 14331
rect 15485 14297 15519 14331
rect 21272 14297 21306 14331
rect 27997 14297 28031 14331
rect 15117 14229 15151 14263
rect 20177 14229 20211 14263
rect 25697 14229 25731 14263
rect 17259 14025 17293 14059
rect 17969 14025 18003 14059
rect 18705 14025 18739 14059
rect 20913 14025 20947 14059
rect 25329 14025 25363 14059
rect 27905 14025 27939 14059
rect 15577 13957 15611 13991
rect 17049 13957 17083 13991
rect 24961 13957 24995 13991
rect 26985 13957 27019 13991
rect 27353 13957 27387 13991
rect 13369 13889 13403 13923
rect 13636 13889 13670 13923
rect 15393 13889 15427 13923
rect 17877 13889 17911 13923
rect 18061 13889 18095 13923
rect 18613 13889 18647 13923
rect 19533 13889 19567 13923
rect 19800 13889 19834 13923
rect 23305 13889 23339 13923
rect 23397 13889 23431 13923
rect 25145 13889 25179 13923
rect 25789 13889 25823 13923
rect 25973 13889 26007 13923
rect 27169 13889 27203 13923
rect 27813 13889 27847 13923
rect 1501 13821 1535 13855
rect 1685 13821 1719 13855
rect 1961 13821 1995 13855
rect 23121 13821 23155 13855
rect 14749 13753 14783 13787
rect 15761 13685 15795 13719
rect 17233 13685 17267 13719
rect 17417 13685 17451 13719
rect 25973 13685 26007 13719
rect 1961 13481 1995 13515
rect 14105 13481 14139 13515
rect 15577 13481 15611 13515
rect 16313 13481 16347 13515
rect 19901 13481 19935 13515
rect 25697 13481 25731 13515
rect 25881 13481 25915 13515
rect 24869 13413 24903 13447
rect 21557 13345 21591 13379
rect 21741 13345 21775 13379
rect 23121 13345 23155 13379
rect 27537 13345 27571 13379
rect 2053 13277 2087 13311
rect 14289 13277 14323 13311
rect 16221 13277 16255 13311
rect 16405 13277 16439 13311
rect 16957 13277 16991 13311
rect 20085 13277 20119 13311
rect 22845 13277 22879 13311
rect 24777 13277 24811 13311
rect 24961 13277 24995 13311
rect 25421 13277 25455 13311
rect 26341 13277 26375 13311
rect 15393 13209 15427 13243
rect 17224 13209 17258 13243
rect 21465 13209 21499 13243
rect 26525 13209 26559 13243
rect 15593 13141 15627 13175
rect 15761 13141 15795 13175
rect 18337 13141 18371 13175
rect 21097 13141 21131 13175
rect 16129 12937 16163 12971
rect 23213 12937 23247 12971
rect 24317 12937 24351 12971
rect 24685 12937 24719 12971
rect 28089 12937 28123 12971
rect 17509 12869 17543 12903
rect 1593 12801 1627 12835
rect 14749 12801 14783 12835
rect 15016 12801 15050 12835
rect 17693 12801 17727 12835
rect 20821 12801 20855 12835
rect 21005 12801 21039 12835
rect 22100 12801 22134 12835
rect 24225 12801 24259 12835
rect 25605 12801 25639 12835
rect 25881 12801 25915 12835
rect 27169 12801 27203 12835
rect 27445 12801 27479 12835
rect 27997 12801 28031 12835
rect 17325 12733 17359 12767
rect 21833 12733 21867 12767
rect 24133 12733 24167 12767
rect 27353 12733 27387 12767
rect 27261 12665 27295 12699
rect 21189 12597 21223 12631
rect 26985 12597 27019 12631
rect 15577 12393 15611 12427
rect 17233 12393 17267 12427
rect 21281 12393 21315 12427
rect 23857 12393 23891 12427
rect 27721 12393 27755 12427
rect 26893 12325 26927 12359
rect 22477 12257 22511 12291
rect 26433 12257 26467 12291
rect 1501 12189 1535 12223
rect 15761 12189 15795 12223
rect 17417 12189 17451 12223
rect 19257 12189 19291 12223
rect 21097 12189 21131 12223
rect 24593 12189 24627 12223
rect 26893 12189 26927 12223
rect 27169 12189 27203 12223
rect 27629 12189 27663 12223
rect 27813 12189 27847 12223
rect 22744 12121 22778 12155
rect 26249 12121 26283 12155
rect 19349 12053 19383 12087
rect 27077 12053 27111 12087
rect 19165 11849 19199 11883
rect 19625 11849 19659 11883
rect 22845 11849 22879 11883
rect 23489 11849 23523 11883
rect 23949 11849 23983 11883
rect 24961 11849 24995 11883
rect 25973 11849 26007 11883
rect 17693 11781 17727 11815
rect 19809 11781 19843 11815
rect 23857 11781 23891 11815
rect 25605 11781 25639 11815
rect 25789 11781 25823 11815
rect 1501 11713 1535 11747
rect 17325 11713 17359 11747
rect 17785 11713 17819 11747
rect 18705 11713 18739 11747
rect 19993 11713 20027 11747
rect 20545 11713 20579 11747
rect 20637 11713 20671 11747
rect 23029 11713 23063 11747
rect 24869 11713 24903 11747
rect 27997 11713 28031 11747
rect 1685 11645 1719 11679
rect 1961 11645 1995 11679
rect 24041 11645 24075 11679
rect 19073 11577 19107 11611
rect 17509 11509 17543 11543
rect 20821 11509 20855 11543
rect 27353 11509 27387 11543
rect 1869 11305 1903 11339
rect 18705 11305 18739 11339
rect 25881 11305 25915 11339
rect 21189 11237 21223 11271
rect 17325 11169 17359 11203
rect 20729 11169 20763 11203
rect 27537 11169 27571 11203
rect 28181 11169 28215 11203
rect 1961 11101 1995 11135
rect 15393 11101 15427 11135
rect 16497 11101 16531 11135
rect 16681 11101 16715 11135
rect 17592 11101 17626 11135
rect 20473 11101 20507 11135
rect 21373 11101 21407 11135
rect 27997 11033 28031 11067
rect 15577 10965 15611 10999
rect 16313 10965 16347 10999
rect 19349 10965 19383 10999
rect 18061 10761 18095 10795
rect 20545 10761 20579 10795
rect 20913 10761 20947 10795
rect 27813 10761 27847 10795
rect 15945 10625 15979 10659
rect 16681 10625 16715 10659
rect 16937 10625 16971 10659
rect 27721 10625 27755 10659
rect 20269 10557 20303 10591
rect 20453 10557 20487 10591
rect 25973 10557 26007 10591
rect 26249 10557 26283 10591
rect 26433 10557 26467 10591
rect 27077 10557 27111 10591
rect 16129 10489 16163 10523
rect 1501 10421 1535 10455
rect 16773 10217 16807 10251
rect 17417 10081 17451 10115
rect 25329 10081 25363 10115
rect 26801 10081 26835 10115
rect 26985 10081 27019 10115
rect 1777 10013 1811 10047
rect 2421 10013 2455 10047
rect 3065 10013 3099 10047
rect 17141 10013 17175 10047
rect 24685 10013 24719 10047
rect 27445 10013 27479 10047
rect 24593 9945 24627 9979
rect 1685 9877 1719 9911
rect 2329 9877 2363 9911
rect 17233 9877 17267 9911
rect 27537 9877 27571 9911
rect 27169 9673 27203 9707
rect 3617 9605 3651 9639
rect 3801 9537 3835 9571
rect 26433 9537 26467 9571
rect 27261 9537 27295 9571
rect 27721 9537 27755 9571
rect 3249 9469 3283 9503
rect 24869 9469 24903 9503
rect 26249 9469 26283 9503
rect 27813 9401 27847 9435
rect 25237 9129 25271 9163
rect 1409 8993 1443 9027
rect 1593 8993 1627 9027
rect 1869 8993 1903 9027
rect 26341 8993 26375 9027
rect 26525 8993 26559 9027
rect 24685 8925 24719 8959
rect 25145 8925 25179 8959
rect 28181 8857 28215 8891
rect 27353 8449 27387 8483
rect 2973 8381 3007 8415
rect 3157 8381 3191 8415
rect 3433 8381 3467 8415
rect 25973 8381 26007 8415
rect 26249 8381 26283 8415
rect 26433 8381 26467 8415
rect 27261 8313 27295 8347
rect 1593 8245 1627 8279
rect 27997 8245 28031 8279
rect 1961 8041 1995 8075
rect 2973 8041 3007 8075
rect 3893 8041 3927 8075
rect 25789 8041 25823 8075
rect 27537 7905 27571 7939
rect 28181 7905 28215 7939
rect 2053 7837 2087 7871
rect 3985 7837 4019 7871
rect 4629 7837 4663 7871
rect 25697 7837 25731 7871
rect 27997 7769 28031 7803
rect 4537 7701 4571 7735
rect 3985 7429 4019 7463
rect 24777 7429 24811 7463
rect 1501 7361 1535 7395
rect 24593 7361 24627 7395
rect 26985 7361 27019 7395
rect 1685 7293 1719 7327
rect 2881 7293 2915 7327
rect 3801 7293 3835 7327
rect 4261 7293 4295 7327
rect 26157 7293 26191 7327
rect 28089 7157 28123 7191
rect 1961 6953 1995 6987
rect 3801 6953 3835 6987
rect 27537 6817 27571 6851
rect 28181 6817 28215 6851
rect 2053 6749 2087 6783
rect 27997 6681 28031 6715
rect 27813 6409 27847 6443
rect 27721 6273 27755 6307
rect 1685 6205 1719 6239
rect 2145 6205 2179 6239
rect 2329 6205 2363 6239
rect 2605 6205 2639 6239
rect 27077 6069 27111 6103
rect 2237 5865 2271 5899
rect 18429 5729 18463 5763
rect 26341 5729 26375 5763
rect 2329 5661 2363 5695
rect 2973 5661 3007 5695
rect 18245 5661 18279 5695
rect 26525 5593 26559 5627
rect 28181 5593 28215 5627
rect 2881 5525 2915 5559
rect 27537 5321 27571 5355
rect 2697 5253 2731 5287
rect 17877 5185 17911 5219
rect 22753 5185 22787 5219
rect 27629 5185 27663 5219
rect 2053 5117 2087 5151
rect 2513 5117 2547 5151
rect 3157 5117 3191 5151
rect 4997 4981 5031 5015
rect 17693 4981 17727 5015
rect 22845 4981 22879 5015
rect 3249 4641 3283 4675
rect 4445 4641 4479 4675
rect 6285 4641 6319 4675
rect 21373 4641 21407 4675
rect 27445 4641 27479 4675
rect 27997 4641 28031 4675
rect 20729 4573 20763 4607
rect 28181 4573 28215 4607
rect 1409 4505 1443 4539
rect 3065 4505 3099 4539
rect 6101 4505 6135 4539
rect 20913 4505 20947 4539
rect 20913 4233 20947 4267
rect 19717 4165 19751 4199
rect 1777 4097 1811 4131
rect 2421 4097 2455 4131
rect 5273 4097 5307 4131
rect 9229 4097 9263 4131
rect 10517 4097 10551 4131
rect 20821 4097 20855 4131
rect 28089 4097 28123 4131
rect 2881 4029 2915 4063
rect 3065 4029 3099 4063
rect 3341 4029 3375 4063
rect 13001 4029 13035 4063
rect 13185 4029 13219 4063
rect 13553 4029 13587 4063
rect 18061 4029 18095 4063
rect 19901 4029 19935 4063
rect 21833 4029 21867 4063
rect 1685 3961 1719 3995
rect 5365 3893 5399 3927
rect 6377 3893 6411 3927
rect 7481 3893 7515 3927
rect 9321 3893 9355 3927
rect 10609 3893 10643 3927
rect 26433 3893 26467 3927
rect 26985 3893 27019 3927
rect 2881 3689 2915 3723
rect 12633 3689 12667 3723
rect 13185 3689 13219 3723
rect 18337 3689 18371 3723
rect 25421 3621 25455 3655
rect 5365 3553 5399 3587
rect 5917 3553 5951 3587
rect 9321 3553 9355 3587
rect 9689 3553 9723 3587
rect 21925 3553 21959 3587
rect 26341 3553 26375 3587
rect 27537 3553 27571 3587
rect 1593 3485 1627 3519
rect 2237 3485 2271 3519
rect 2789 3485 2823 3519
rect 4353 3485 4387 3519
rect 5181 3485 5215 3519
rect 7481 3485 7515 3519
rect 8401 3485 8435 3519
rect 9137 3485 9171 3519
rect 11621 3485 11655 3519
rect 13093 3485 13127 3519
rect 14657 3485 14691 3519
rect 15117 3485 15151 3519
rect 16313 3485 16347 3519
rect 16957 3485 16991 3519
rect 19533 3485 19567 3519
rect 20637 3485 20671 3519
rect 21281 3485 21315 3519
rect 24409 3485 24443 3519
rect 25513 3485 25547 3519
rect 20729 3417 20763 3451
rect 21465 3417 21499 3451
rect 26525 3417 26559 3451
rect 2145 3349 2179 3383
rect 4261 3349 4295 3383
rect 7573 3349 7607 3383
rect 14565 3349 14599 3383
rect 16405 3349 16439 3383
rect 19625 3349 19659 3383
rect 27077 3145 27111 3179
rect 1869 3077 1903 3111
rect 4169 3077 4203 3111
rect 8861 3077 8895 3111
rect 11713 3077 11747 3111
rect 14473 3077 14507 3111
rect 16865 3077 16899 3111
rect 19625 3077 19659 3111
rect 23489 3077 23523 3111
rect 24225 3077 24259 3111
rect 1685 3009 1719 3043
rect 6377 3009 6411 3043
rect 8677 3009 8711 3043
rect 11529 3009 11563 3043
rect 14289 3009 14323 3043
rect 16681 3009 16715 3043
rect 21833 3009 21867 3043
rect 23397 3009 23431 3043
rect 24041 3009 24075 3043
rect 26985 3009 27019 3043
rect 27813 3009 27847 3043
rect 2789 2941 2823 2975
rect 3985 2941 4019 2975
rect 4537 2941 4571 2975
rect 6561 2941 6595 2975
rect 6837 2941 6871 2975
rect 9137 2941 9171 2975
rect 11989 2941 12023 2975
rect 14749 2941 14783 2975
rect 17141 2941 17175 2975
rect 19441 2941 19475 2975
rect 19993 2941 20027 2975
rect 25145 2941 25179 2975
rect 27721 2805 27755 2839
rect 2881 2601 2915 2635
rect 4077 2601 4111 2635
rect 5273 2601 5307 2635
rect 6469 2601 6503 2635
rect 9505 2601 9539 2635
rect 16865 2601 16899 2635
rect 17509 2601 17543 2635
rect 19441 2601 19475 2635
rect 25973 2465 26007 2499
rect 26249 2465 26283 2499
rect 26433 2465 26467 2499
rect 27445 2465 27479 2499
rect 6377 2397 6411 2431
rect 16681 2397 16715 2431
rect 17693 2397 17727 2431
rect 27169 2397 27203 2431
rect 9413 2329 9447 2363
<< metal1 >>
rect 1104 47354 28888 47376
rect 1104 47302 5582 47354
rect 5634 47302 5646 47354
rect 5698 47302 5710 47354
rect 5762 47302 5774 47354
rect 5826 47302 5838 47354
rect 5890 47302 14846 47354
rect 14898 47302 14910 47354
rect 14962 47302 14974 47354
rect 15026 47302 15038 47354
rect 15090 47302 15102 47354
rect 15154 47302 24110 47354
rect 24162 47302 24174 47354
rect 24226 47302 24238 47354
rect 24290 47302 24302 47354
rect 24354 47302 24366 47354
rect 24418 47302 28888 47354
rect 1104 47280 28888 47302
rect 23198 47104 23204 47116
rect 23159 47076 23204 47104
rect 23198 47064 23204 47076
rect 23256 47064 23262 47116
rect 25961 47107 26019 47113
rect 25961 47073 25973 47107
rect 26007 47104 26019 47107
rect 28350 47104 28356 47116
rect 26007 47076 28356 47104
rect 26007 47073 26019 47076
rect 25961 47067 26019 47073
rect 28350 47064 28356 47076
rect 28408 47064 28414 47116
rect 1670 46996 1676 47048
rect 1728 47036 1734 47048
rect 1765 47039 1823 47045
rect 1765 47036 1777 47039
rect 1728 47008 1777 47036
rect 1728 46996 1734 47008
rect 1765 47005 1777 47008
rect 1811 47005 1823 47039
rect 1765 46999 1823 47005
rect 2961 47039 3019 47045
rect 2961 47005 2973 47039
rect 3007 47036 3019 47039
rect 3602 47036 3608 47048
rect 3007 47008 3608 47036
rect 3007 47005 3019 47008
rect 2961 46999 3019 47005
rect 3602 46996 3608 47008
rect 3660 46996 3666 47048
rect 3786 47036 3792 47048
rect 3747 47008 3792 47036
rect 3786 46996 3792 47008
rect 3844 46996 3850 47048
rect 6086 46996 6092 47048
rect 6144 47036 6150 47048
rect 6365 47039 6423 47045
rect 6365 47036 6377 47039
rect 6144 47008 6377 47036
rect 6144 46996 6150 47008
rect 6365 47005 6377 47008
rect 6411 47005 6423 47039
rect 7101 47039 7159 47045
rect 7101 47036 7113 47039
rect 6365 46999 6423 47005
rect 6886 47008 7113 47036
rect 2590 46860 2596 46912
rect 2648 46900 2654 46912
rect 3050 46900 3056 46912
rect 2648 46872 3056 46900
rect 2648 46860 2654 46872
rect 3050 46860 3056 46872
rect 3108 46860 3114 46912
rect 6546 46900 6552 46912
rect 6507 46872 6552 46900
rect 6546 46860 6552 46872
rect 6604 46860 6610 46912
rect 6638 46860 6644 46912
rect 6696 46900 6702 46912
rect 6886 46900 6914 47008
rect 7101 47005 7113 47008
rect 7147 47005 7159 47039
rect 7834 47036 7840 47048
rect 7795 47008 7840 47036
rect 7101 46999 7159 47005
rect 7834 46996 7840 47008
rect 7892 46996 7898 47048
rect 13814 46996 13820 47048
rect 13872 47036 13878 47048
rect 14093 47039 14151 47045
rect 14093 47036 14105 47039
rect 13872 47008 14105 47036
rect 13872 46996 13878 47008
rect 14093 47005 14105 47008
rect 14139 47005 14151 47039
rect 16666 47036 16672 47048
rect 16627 47008 16672 47036
rect 14093 46999 14151 47005
rect 16666 46996 16672 47008
rect 16724 46996 16730 47048
rect 18138 47036 18144 47048
rect 18099 47008 18144 47036
rect 18138 46996 18144 47008
rect 18196 46996 18202 47048
rect 19334 46996 19340 47048
rect 19392 47036 19398 47048
rect 19429 47039 19487 47045
rect 19429 47036 19441 47039
rect 19392 47008 19441 47036
rect 19392 46996 19398 47008
rect 19429 47005 19441 47008
rect 19475 47005 19487 47039
rect 19429 46999 19487 47005
rect 21910 46996 21916 47048
rect 21968 47036 21974 47048
rect 22005 47039 22063 47045
rect 22005 47036 22017 47039
rect 21968 47008 22017 47036
rect 21968 46996 21974 47008
rect 22005 47005 22017 47008
rect 22051 47005 22063 47039
rect 22005 46999 22063 47005
rect 26421 47039 26479 47045
rect 26421 47005 26433 47039
rect 26467 47036 26479 47039
rect 26973 47039 27031 47045
rect 26973 47036 26985 47039
rect 26467 47008 26985 47036
rect 26467 47005 26479 47008
rect 26421 46999 26479 47005
rect 26973 47005 26985 47008
rect 27019 47005 27031 47039
rect 26973 46999 27031 47005
rect 28077 47039 28135 47045
rect 28077 47005 28089 47039
rect 28123 47036 28135 47039
rect 28166 47036 28172 47048
rect 28123 47008 28172 47036
rect 28123 47005 28135 47008
rect 28077 46999 28135 47005
rect 28166 46996 28172 47008
rect 28224 46996 28230 47048
rect 22189 46971 22247 46977
rect 22189 46937 22201 46971
rect 22235 46968 22247 46971
rect 22738 46968 22744 46980
rect 22235 46940 22744 46968
rect 22235 46937 22247 46940
rect 22189 46931 22247 46937
rect 22738 46928 22744 46940
rect 22796 46928 22802 46980
rect 26234 46928 26240 46980
rect 26292 46968 26298 46980
rect 26292 46940 26337 46968
rect 26292 46928 26298 46940
rect 7282 46900 7288 46912
rect 6696 46872 6914 46900
rect 7243 46872 7288 46900
rect 6696 46860 6702 46872
rect 7282 46860 7288 46872
rect 7340 46860 7346 46912
rect 11606 46860 11612 46912
rect 11664 46900 11670 46912
rect 12526 46900 12532 46912
rect 11664 46872 12532 46900
rect 11664 46860 11670 46872
rect 12526 46860 12532 46872
rect 12584 46860 12590 46912
rect 27062 46860 27068 46912
rect 27120 46900 27126 46912
rect 28074 46900 28080 46912
rect 27120 46872 28080 46900
rect 27120 46860 27126 46872
rect 28074 46860 28080 46872
rect 28132 46860 28138 46912
rect 1104 46810 28888 46832
rect 1104 46758 10214 46810
rect 10266 46758 10278 46810
rect 10330 46758 10342 46810
rect 10394 46758 10406 46810
rect 10458 46758 10470 46810
rect 10522 46758 19478 46810
rect 19530 46758 19542 46810
rect 19594 46758 19606 46810
rect 19658 46758 19670 46810
rect 19722 46758 19734 46810
rect 19786 46758 28888 46810
rect 1104 46736 28888 46758
rect 23842 46696 23848 46708
rect 23216 46668 23848 46696
rect 23216 46637 23244 46668
rect 23842 46656 23848 46668
rect 23900 46656 23906 46708
rect 26234 46656 26240 46708
rect 26292 46696 26298 46708
rect 27065 46699 27123 46705
rect 27065 46696 27077 46699
rect 26292 46668 27077 46696
rect 26292 46656 26298 46668
rect 27065 46665 27077 46668
rect 27111 46665 27123 46699
rect 27065 46659 27123 46665
rect 23201 46631 23259 46637
rect 23201 46597 23213 46631
rect 23247 46597 23259 46631
rect 25590 46628 25596 46640
rect 25551 46600 25596 46628
rect 23201 46591 23259 46597
rect 25590 46588 25596 46600
rect 25648 46588 25654 46640
rect 1670 46560 1676 46572
rect 1631 46532 1676 46560
rect 1670 46520 1676 46532
rect 1728 46520 1734 46572
rect 3602 46520 3608 46572
rect 3660 46560 3666 46572
rect 3973 46563 4031 46569
rect 3973 46560 3985 46563
rect 3660 46532 3985 46560
rect 3660 46520 3666 46532
rect 3973 46529 3985 46532
rect 4019 46529 4031 46563
rect 7834 46560 7840 46572
rect 7795 46532 7840 46560
rect 3973 46523 4031 46529
rect 7834 46520 7840 46532
rect 7892 46520 7898 46572
rect 13814 46560 13820 46572
rect 13775 46532 13820 46560
rect 13814 46520 13820 46532
rect 13872 46520 13878 46572
rect 16666 46560 16672 46572
rect 16627 46532 16672 46560
rect 16666 46520 16672 46532
rect 16724 46520 16730 46572
rect 19334 46520 19340 46572
rect 19392 46560 19398 46572
rect 19429 46563 19487 46569
rect 19429 46560 19441 46563
rect 19392 46532 19441 46560
rect 19392 46520 19398 46532
rect 19429 46529 19441 46532
rect 19475 46529 19487 46563
rect 26970 46560 26976 46572
rect 26931 46532 26976 46560
rect 19429 46523 19487 46529
rect 26970 46520 26976 46532
rect 27028 46520 27034 46572
rect 1857 46495 1915 46501
rect 1857 46461 1869 46495
rect 1903 46492 1915 46495
rect 2130 46492 2136 46504
rect 1903 46464 2136 46492
rect 1903 46461 1915 46464
rect 1857 46455 1915 46461
rect 2130 46452 2136 46464
rect 2188 46452 2194 46504
rect 2225 46495 2283 46501
rect 2225 46461 2237 46495
rect 2271 46461 2283 46495
rect 4154 46492 4160 46504
rect 4115 46464 4160 46492
rect 2225 46455 2283 46461
rect 1302 46384 1308 46436
rect 1360 46424 1366 46436
rect 2240 46424 2268 46455
rect 4154 46452 4160 46464
rect 4212 46452 4218 46504
rect 4433 46495 4491 46501
rect 4433 46461 4445 46495
rect 4479 46461 4491 46495
rect 8018 46492 8024 46504
rect 7979 46464 8024 46492
rect 4433 46455 4491 46461
rect 1360 46396 2268 46424
rect 1360 46384 1366 46396
rect 2314 46384 2320 46436
rect 2372 46424 2378 46436
rect 4448 46424 4476 46455
rect 8018 46452 8024 46464
rect 8076 46452 8082 46504
rect 8386 46492 8392 46504
rect 8347 46464 8392 46492
rect 8386 46452 8392 46464
rect 8444 46452 8450 46504
rect 10965 46495 11023 46501
rect 10965 46461 10977 46495
rect 11011 46492 11023 46495
rect 11517 46495 11575 46501
rect 11517 46492 11529 46495
rect 11011 46464 11529 46492
rect 11011 46461 11023 46464
rect 10965 46455 11023 46461
rect 11517 46461 11529 46464
rect 11563 46461 11575 46495
rect 11698 46492 11704 46504
rect 11659 46464 11704 46492
rect 11517 46455 11575 46461
rect 11698 46452 11704 46464
rect 11756 46452 11762 46504
rect 11977 46495 12035 46501
rect 11977 46461 11989 46495
rect 12023 46461 12035 46495
rect 11977 46455 12035 46461
rect 11992 46424 12020 46455
rect 13446 46452 13452 46504
rect 13504 46492 13510 46504
rect 14001 46495 14059 46501
rect 14001 46492 14013 46495
rect 13504 46464 14013 46492
rect 13504 46452 13510 46464
rect 14001 46461 14013 46464
rect 14047 46461 14059 46495
rect 14001 46455 14059 46461
rect 14277 46495 14335 46501
rect 14277 46461 14289 46495
rect 14323 46461 14335 46495
rect 16850 46492 16856 46504
rect 16811 46464 16856 46492
rect 14277 46455 14335 46461
rect 2372 46396 4476 46424
rect 10980 46396 12020 46424
rect 2372 46384 2378 46396
rect 10980 46368 11008 46396
rect 13538 46384 13544 46436
rect 13596 46424 13602 46436
rect 14292 46424 14320 46455
rect 16850 46452 16856 46464
rect 16908 46452 16914 46504
rect 17129 46495 17187 46501
rect 17129 46461 17141 46495
rect 17175 46461 17187 46495
rect 19613 46495 19671 46501
rect 19613 46492 19625 46495
rect 17129 46455 17187 46461
rect 19352 46464 19625 46492
rect 13596 46396 14320 46424
rect 13596 46384 13602 46396
rect 16758 46384 16764 46436
rect 16816 46424 16822 46436
rect 17144 46424 17172 46455
rect 19352 46436 19380 46464
rect 19613 46461 19625 46464
rect 19659 46461 19671 46495
rect 19978 46492 19984 46504
rect 19939 46464 19984 46492
rect 19613 46455 19671 46461
rect 19978 46452 19984 46464
rect 20036 46452 20042 46504
rect 23750 46492 23756 46504
rect 23711 46464 23756 46492
rect 23750 46452 23756 46464
rect 23808 46452 23814 46504
rect 23934 46492 23940 46504
rect 23895 46464 23940 46492
rect 23934 46452 23940 46464
rect 23992 46452 23998 46504
rect 16816 46396 17172 46424
rect 16816 46384 16822 46396
rect 19334 46384 19340 46436
rect 19392 46384 19398 46436
rect 23017 46427 23075 46433
rect 23017 46424 23029 46427
rect 19444 46396 23029 46424
rect 9582 46316 9588 46368
rect 9640 46356 9646 46368
rect 10137 46359 10195 46365
rect 10137 46356 10149 46359
rect 9640 46328 10149 46356
rect 9640 46316 9646 46328
rect 10137 46325 10149 46328
rect 10183 46325 10195 46359
rect 10137 46319 10195 46325
rect 10962 46316 10968 46368
rect 11020 46316 11026 46368
rect 17586 46316 17592 46368
rect 17644 46356 17650 46368
rect 19444 46356 19472 46396
rect 23017 46393 23029 46396
rect 23063 46393 23075 46427
rect 23017 46387 23075 46393
rect 17644 46328 19472 46356
rect 17644 46316 17650 46328
rect 22002 46316 22008 46368
rect 22060 46356 22066 46368
rect 22097 46359 22155 46365
rect 22097 46356 22109 46359
rect 22060 46328 22109 46356
rect 22060 46316 22066 46328
rect 22097 46325 22109 46328
rect 22143 46325 22155 46359
rect 22097 46319 22155 46325
rect 26329 46359 26387 46365
rect 26329 46325 26341 46359
rect 26375 46356 26387 46359
rect 26418 46356 26424 46368
rect 26375 46328 26424 46356
rect 26375 46325 26387 46328
rect 26329 46319 26387 46325
rect 26418 46316 26424 46328
rect 26476 46316 26482 46368
rect 27890 46356 27896 46368
rect 27851 46328 27896 46356
rect 27890 46316 27896 46328
rect 27948 46316 27954 46368
rect 1104 46266 28888 46288
rect 1104 46214 5582 46266
rect 5634 46214 5646 46266
rect 5698 46214 5710 46266
rect 5762 46214 5774 46266
rect 5826 46214 5838 46266
rect 5890 46214 14846 46266
rect 14898 46214 14910 46266
rect 14962 46214 14974 46266
rect 15026 46214 15038 46266
rect 15090 46214 15102 46266
rect 15154 46214 24110 46266
rect 24162 46214 24174 46266
rect 24226 46214 24238 46266
rect 24290 46214 24302 46266
rect 24354 46214 24366 46266
rect 24418 46214 28888 46266
rect 1104 46192 28888 46214
rect 2130 46152 2136 46164
rect 2091 46124 2136 46152
rect 2130 46112 2136 46124
rect 2188 46112 2194 46164
rect 3145 46155 3203 46161
rect 3145 46121 3157 46155
rect 3191 46152 3203 46155
rect 4154 46152 4160 46164
rect 3191 46124 4160 46152
rect 3191 46121 3203 46124
rect 3145 46115 3203 46121
rect 4154 46112 4160 46124
rect 4212 46112 4218 46164
rect 8018 46152 8024 46164
rect 7979 46124 8024 46152
rect 8018 46112 8024 46124
rect 8076 46112 8082 46164
rect 13446 46152 13452 46164
rect 13407 46124 13452 46152
rect 13446 46112 13452 46124
rect 13504 46112 13510 46164
rect 16669 46155 16727 46161
rect 16669 46121 16681 46155
rect 16715 46152 16727 46155
rect 16850 46152 16856 46164
rect 16715 46124 16856 46152
rect 16715 46121 16727 46124
rect 16669 46115 16727 46121
rect 16850 46112 16856 46124
rect 16908 46112 16914 46164
rect 23750 46112 23756 46164
rect 23808 46152 23814 46164
rect 24397 46155 24455 46161
rect 24397 46152 24409 46155
rect 23808 46124 24409 46152
rect 23808 46112 23814 46124
rect 24397 46121 24409 46124
rect 24443 46121 24455 46155
rect 24397 46115 24455 46121
rect 4982 46084 4988 46096
rect 2240 46056 4988 46084
rect 1578 45948 1584 45960
rect 1539 45920 1584 45948
rect 1578 45908 1584 45920
rect 1636 45908 1642 45960
rect 2240 45957 2268 46056
rect 4982 46044 4988 46056
rect 5040 46044 5046 46096
rect 26970 46084 26976 46096
rect 7944 46056 26976 46084
rect 3786 46016 3792 46028
rect 3747 45988 3792 46016
rect 3786 45976 3792 45988
rect 3844 45976 3850 46028
rect 4062 45976 4068 46028
rect 4120 46016 4126 46028
rect 4249 46019 4307 46025
rect 4249 46016 4261 46019
rect 4120 45988 4261 46016
rect 4120 45976 4126 45988
rect 4249 45985 4261 45988
rect 4295 45985 4307 46019
rect 4249 45979 4307 45985
rect 7944 45957 7972 46056
rect 26970 46044 26976 46056
rect 27028 46044 27034 46096
rect 9582 46016 9588 46028
rect 9543 45988 9588 46016
rect 9582 45976 9588 45988
rect 9640 45976 9646 46028
rect 10134 46016 10140 46028
rect 10095 45988 10140 46016
rect 10134 45976 10140 45988
rect 10192 45976 10198 46028
rect 19705 46019 19763 46025
rect 12406 45988 18276 46016
rect 2225 45951 2283 45957
rect 2225 45917 2237 45951
rect 2271 45917 2283 45951
rect 2225 45911 2283 45917
rect 3237 45951 3295 45957
rect 3237 45917 3249 45951
rect 3283 45917 3295 45951
rect 3237 45911 3295 45917
rect 7929 45951 7987 45957
rect 7929 45917 7941 45951
rect 7975 45917 7987 45951
rect 7929 45911 7987 45917
rect 3252 45812 3280 45911
rect 3973 45883 4031 45889
rect 3973 45849 3985 45883
rect 4019 45880 4031 45883
rect 4522 45880 4528 45892
rect 4019 45852 4528 45880
rect 4019 45849 4031 45852
rect 3973 45843 4031 45849
rect 4522 45840 4528 45852
rect 4580 45840 4586 45892
rect 9769 45883 9827 45889
rect 9769 45849 9781 45883
rect 9815 45880 9827 45883
rect 9858 45880 9864 45892
rect 9815 45852 9864 45880
rect 9815 45849 9827 45852
rect 9769 45843 9827 45849
rect 9858 45840 9864 45852
rect 9916 45840 9922 45892
rect 12406 45812 12434 45988
rect 18248 45960 18276 45988
rect 19705 45985 19717 46019
rect 19751 46016 19763 46019
rect 20162 46016 20168 46028
rect 19751 45988 20168 46016
rect 19751 45985 19763 45988
rect 19705 45979 19763 45985
rect 20162 45976 20168 45988
rect 20220 45976 20226 46028
rect 21266 46016 21272 46028
rect 21227 45988 21272 46016
rect 21266 45976 21272 45988
rect 21324 45976 21330 46028
rect 22002 46016 22008 46028
rect 21963 45988 22008 46016
rect 22002 45976 22008 45988
rect 22060 45976 22066 46028
rect 22554 46016 22560 46028
rect 22515 45988 22560 46016
rect 22554 45976 22560 45988
rect 22612 45976 22618 46028
rect 26142 45976 26148 46028
rect 26200 46016 26206 46028
rect 26329 46019 26387 46025
rect 26329 46016 26341 46019
rect 26200 45988 26341 46016
rect 26200 45976 26206 45988
rect 26329 45985 26341 45988
rect 26375 45985 26387 46019
rect 28166 46016 28172 46028
rect 28127 45988 28172 46016
rect 26329 45979 26387 45985
rect 28166 45976 28172 45988
rect 28224 45976 28230 46028
rect 13541 45951 13599 45957
rect 13541 45917 13553 45951
rect 13587 45917 13599 45951
rect 14274 45948 14280 45960
rect 14235 45920 14280 45948
rect 13541 45911 13599 45917
rect 3252 45784 12434 45812
rect 13556 45812 13584 45911
rect 14274 45908 14280 45920
rect 14332 45908 14338 45960
rect 16577 45951 16635 45957
rect 16577 45917 16589 45951
rect 16623 45917 16635 45951
rect 18230 45948 18236 45960
rect 18143 45920 18236 45948
rect 16577 45911 16635 45917
rect 14458 45880 14464 45892
rect 14419 45852 14464 45880
rect 14458 45840 14464 45852
rect 14516 45840 14522 45892
rect 14734 45840 14740 45892
rect 14792 45880 14798 45892
rect 16117 45883 16175 45889
rect 16117 45880 16129 45883
rect 14792 45852 16129 45880
rect 14792 45840 14798 45852
rect 16117 45849 16129 45852
rect 16163 45849 16175 45883
rect 16592 45880 16620 45911
rect 18230 45908 18236 45920
rect 18288 45908 18294 45960
rect 25774 45908 25780 45960
rect 25832 45948 25838 45960
rect 25869 45951 25927 45957
rect 25869 45948 25881 45951
rect 25832 45920 25881 45948
rect 25832 45908 25838 45920
rect 25869 45917 25881 45920
rect 25915 45917 25927 45951
rect 25869 45911 25927 45917
rect 19886 45880 19892 45892
rect 16592 45852 19380 45880
rect 19847 45852 19892 45880
rect 16117 45843 16175 45849
rect 18046 45812 18052 45824
rect 13556 45784 18052 45812
rect 18046 45772 18052 45784
rect 18104 45772 18110 45824
rect 18322 45812 18328 45824
rect 18283 45784 18328 45812
rect 18322 45772 18328 45784
rect 18380 45772 18386 45824
rect 19352 45812 19380 45852
rect 19886 45840 19892 45852
rect 19944 45840 19950 45892
rect 22186 45880 22192 45892
rect 22147 45852 22192 45880
rect 22186 45840 22192 45852
rect 22244 45840 22250 45892
rect 22296 45852 26924 45880
rect 22296 45812 22324 45852
rect 26896 45824 26924 45852
rect 27522 45840 27528 45892
rect 27580 45880 27586 45892
rect 27985 45883 28043 45889
rect 27985 45880 27997 45883
rect 27580 45852 27997 45880
rect 27580 45840 27586 45852
rect 27985 45849 27997 45852
rect 28031 45849 28043 45883
rect 27985 45843 28043 45849
rect 19352 45784 22324 45812
rect 25777 45815 25835 45821
rect 25777 45781 25789 45815
rect 25823 45812 25835 45815
rect 26234 45812 26240 45824
rect 25823 45784 26240 45812
rect 25823 45781 25835 45784
rect 25777 45775 25835 45781
rect 26234 45772 26240 45784
rect 26292 45772 26298 45824
rect 26878 45772 26884 45824
rect 26936 45812 26942 45824
rect 27430 45812 27436 45824
rect 26936 45784 27436 45812
rect 26936 45772 26942 45784
rect 27430 45772 27436 45784
rect 27488 45772 27494 45824
rect 1104 45722 28888 45744
rect 1104 45670 10214 45722
rect 10266 45670 10278 45722
rect 10330 45670 10342 45722
rect 10394 45670 10406 45722
rect 10458 45670 10470 45722
rect 10522 45670 19478 45722
rect 19530 45670 19542 45722
rect 19594 45670 19606 45722
rect 19658 45670 19670 45722
rect 19722 45670 19734 45722
rect 19786 45670 28888 45722
rect 1104 45648 28888 45670
rect 9858 45608 9864 45620
rect 9819 45580 9864 45608
rect 9858 45568 9864 45580
rect 9916 45568 9922 45620
rect 14458 45608 14464 45620
rect 14419 45580 14464 45608
rect 14458 45568 14464 45580
rect 14516 45568 14522 45620
rect 18046 45568 18052 45620
rect 18104 45608 18110 45620
rect 18104 45580 19564 45608
rect 18104 45568 18110 45580
rect 19536 45552 19564 45580
rect 19886 45568 19892 45620
rect 19944 45608 19950 45620
rect 20533 45611 20591 45617
rect 20533 45608 20545 45611
rect 19944 45580 20545 45608
rect 19944 45568 19950 45580
rect 20533 45577 20545 45580
rect 20579 45577 20591 45611
rect 20533 45571 20591 45577
rect 22097 45611 22155 45617
rect 22097 45577 22109 45611
rect 22143 45608 22155 45611
rect 22186 45608 22192 45620
rect 22143 45580 22192 45608
rect 22143 45577 22155 45580
rect 22097 45571 22155 45577
rect 22186 45568 22192 45580
rect 22244 45568 22250 45620
rect 4522 45540 4528 45552
rect 4483 45512 4528 45540
rect 4522 45500 4528 45512
rect 4580 45500 4586 45552
rect 10689 45543 10747 45549
rect 10689 45509 10701 45543
rect 10735 45540 10747 45543
rect 11698 45540 11704 45552
rect 10735 45512 11704 45540
rect 10735 45509 10747 45512
rect 10689 45503 10747 45509
rect 11698 45500 11704 45512
rect 11756 45500 11762 45552
rect 18322 45540 18328 45552
rect 18283 45512 18328 45540
rect 18322 45500 18328 45512
rect 18380 45500 18386 45552
rect 19518 45500 19524 45552
rect 19576 45500 19582 45552
rect 22738 45540 22744 45552
rect 22699 45512 22744 45540
rect 22738 45500 22744 45512
rect 22796 45500 22802 45552
rect 23385 45543 23443 45549
rect 23385 45509 23397 45543
rect 23431 45540 23443 45543
rect 23934 45540 23940 45552
rect 23431 45512 23940 45540
rect 23431 45509 23443 45512
rect 23385 45503 23443 45509
rect 23934 45500 23940 45512
rect 23992 45500 23998 45552
rect 26234 45500 26240 45552
rect 26292 45540 26298 45552
rect 27522 45540 27528 45552
rect 26292 45512 26337 45540
rect 27483 45512 27528 45540
rect 26292 45500 26298 45512
rect 27522 45500 27528 45512
rect 27580 45500 27586 45552
rect 1578 45472 1584 45484
rect 1539 45444 1584 45472
rect 1578 45432 1584 45444
rect 1636 45432 1642 45484
rect 4617 45475 4675 45481
rect 4617 45441 4629 45475
rect 4663 45472 4675 45475
rect 5442 45472 5448 45484
rect 4663 45444 5448 45472
rect 4663 45441 4675 45444
rect 4617 45435 4675 45441
rect 5442 45432 5448 45444
rect 5500 45432 5506 45484
rect 9950 45472 9956 45484
rect 9911 45444 9956 45472
rect 9950 45432 9956 45444
rect 10008 45472 10014 45484
rect 10597 45475 10655 45481
rect 10597 45472 10609 45475
rect 10008 45444 10609 45472
rect 10008 45432 10014 45444
rect 10597 45441 10609 45444
rect 10643 45441 10655 45475
rect 14366 45472 14372 45484
rect 14327 45444 14372 45472
rect 10597 45435 10655 45441
rect 14366 45432 14372 45444
rect 14424 45432 14430 45484
rect 18138 45472 18144 45484
rect 18099 45444 18144 45472
rect 18138 45432 18144 45444
rect 18196 45432 18202 45484
rect 20438 45472 20444 45484
rect 20399 45444 20444 45472
rect 20438 45432 20444 45444
rect 20496 45432 20502 45484
rect 22002 45472 22008 45484
rect 21963 45444 22008 45472
rect 22002 45432 22008 45444
rect 22060 45432 22066 45484
rect 22833 45475 22891 45481
rect 22833 45441 22845 45475
rect 22879 45441 22891 45475
rect 23290 45472 23296 45484
rect 23251 45444 23296 45472
rect 22833 45435 22891 45441
rect 1765 45407 1823 45413
rect 1765 45373 1777 45407
rect 1811 45404 1823 45407
rect 1946 45404 1952 45416
rect 1811 45376 1952 45404
rect 1811 45373 1823 45376
rect 1765 45367 1823 45373
rect 1946 45364 1952 45376
rect 2004 45364 2010 45416
rect 2041 45407 2099 45413
rect 2041 45373 2053 45407
rect 2087 45373 2099 45407
rect 2041 45367 2099 45373
rect 14 45296 20 45348
rect 72 45336 78 45348
rect 2056 45336 2084 45367
rect 14274 45364 14280 45416
rect 14332 45404 14338 45416
rect 15013 45407 15071 45413
rect 15013 45404 15025 45407
rect 14332 45376 15025 45404
rect 14332 45364 14338 45376
rect 15013 45373 15025 45376
rect 15059 45373 15071 45407
rect 18690 45404 18696 45416
rect 18651 45376 18696 45404
rect 15013 45367 15071 45373
rect 18690 45364 18696 45376
rect 18748 45364 18754 45416
rect 22848 45404 22876 45435
rect 23290 45432 23296 45444
rect 23348 45432 23354 45484
rect 26418 45432 26424 45484
rect 26476 45472 26482 45484
rect 27430 45472 27436 45484
rect 26476 45444 26521 45472
rect 27391 45444 27436 45472
rect 26476 45432 26482 45444
rect 27430 45432 27436 45444
rect 27488 45432 27494 45484
rect 25774 45404 25780 45416
rect 22848 45376 25780 45404
rect 72 45308 2084 45336
rect 72 45296 78 45308
rect 5442 45296 5448 45348
rect 5500 45336 5506 45348
rect 22848 45336 22876 45376
rect 25774 45364 25780 45376
rect 25832 45364 25838 45416
rect 25958 45404 25964 45416
rect 25919 45376 25964 45404
rect 25958 45364 25964 45376
rect 26016 45364 26022 45416
rect 5500 45308 22876 45336
rect 5500 45296 5506 45308
rect 1104 45178 28888 45200
rect 1104 45126 5582 45178
rect 5634 45126 5646 45178
rect 5698 45126 5710 45178
rect 5762 45126 5774 45178
rect 5826 45126 5838 45178
rect 5890 45126 14846 45178
rect 14898 45126 14910 45178
rect 14962 45126 14974 45178
rect 15026 45126 15038 45178
rect 15090 45126 15102 45178
rect 15154 45126 24110 45178
rect 24162 45126 24174 45178
rect 24226 45126 24238 45178
rect 24290 45126 24302 45178
rect 24354 45126 24366 45178
rect 24418 45126 28888 45178
rect 1104 45104 28888 45126
rect 1946 45064 1952 45076
rect 1907 45036 1952 45064
rect 1946 45024 1952 45036
rect 2004 45024 2010 45076
rect 19334 45024 19340 45076
rect 19392 45064 19398 45076
rect 19521 45067 19579 45073
rect 19521 45064 19533 45067
rect 19392 45036 19533 45064
rect 19392 45024 19398 45036
rect 19521 45033 19533 45036
rect 19567 45033 19579 45067
rect 20162 45064 20168 45076
rect 20123 45036 20168 45064
rect 19521 45027 19579 45033
rect 20162 45024 20168 45036
rect 20220 45024 20226 45076
rect 21910 45024 21916 45076
rect 21968 45064 21974 45076
rect 22649 45067 22707 45073
rect 22649 45064 22661 45067
rect 21968 45036 22661 45064
rect 21968 45024 21974 45036
rect 22649 45033 22661 45036
rect 22695 45033 22707 45067
rect 22649 45027 22707 45033
rect 14366 44956 14372 45008
rect 14424 44996 14430 45008
rect 27430 44996 27436 45008
rect 14424 44968 27436 44996
rect 14424 44956 14430 44968
rect 27430 44956 27436 44968
rect 27488 44956 27494 45008
rect 12526 44928 12532 44940
rect 12487 44900 12532 44928
rect 12526 44888 12532 44900
rect 12584 44888 12590 44940
rect 27522 44928 27528 44940
rect 27483 44900 27528 44928
rect 27522 44888 27528 44900
rect 27580 44888 27586 44940
rect 27890 44888 27896 44940
rect 27948 44928 27954 44940
rect 28169 44931 28227 44937
rect 28169 44928 28181 44931
rect 27948 44900 28181 44928
rect 27948 44888 27954 44900
rect 28169 44897 28181 44900
rect 28215 44897 28227 44931
rect 28169 44891 28227 44897
rect 1946 44820 1952 44872
rect 2004 44860 2010 44872
rect 2041 44863 2099 44869
rect 2041 44860 2053 44863
rect 2004 44832 2053 44860
rect 2004 44820 2010 44832
rect 2041 44829 2053 44832
rect 2087 44829 2099 44863
rect 2041 44823 2099 44829
rect 10689 44863 10747 44869
rect 10689 44829 10701 44863
rect 10735 44860 10747 44863
rect 11149 44863 11207 44869
rect 11149 44860 11161 44863
rect 10735 44832 11161 44860
rect 10735 44829 10747 44832
rect 10689 44823 10747 44829
rect 11149 44829 11161 44832
rect 11195 44829 11207 44863
rect 11149 44823 11207 44829
rect 19334 44820 19340 44872
rect 19392 44860 19398 44872
rect 19429 44863 19487 44869
rect 19429 44860 19441 44863
rect 19392 44832 19441 44860
rect 19392 44820 19398 44832
rect 19429 44829 19441 44832
rect 19475 44860 19487 44863
rect 19518 44860 19524 44872
rect 19475 44832 19524 44860
rect 19475 44829 19487 44832
rect 19429 44823 19487 44829
rect 19518 44820 19524 44832
rect 19576 44820 19582 44872
rect 11333 44795 11391 44801
rect 11333 44761 11345 44795
rect 11379 44792 11391 44795
rect 11606 44792 11612 44804
rect 11379 44764 11612 44792
rect 11379 44761 11391 44764
rect 11333 44755 11391 44761
rect 11606 44752 11612 44764
rect 11664 44752 11670 44804
rect 27614 44752 27620 44804
rect 27672 44792 27678 44804
rect 27985 44795 28043 44801
rect 27985 44792 27997 44795
rect 27672 44764 27997 44792
rect 27672 44752 27678 44764
rect 27985 44761 27997 44764
rect 28031 44761 28043 44795
rect 27985 44755 28043 44761
rect 1104 44634 28888 44656
rect 1104 44582 10214 44634
rect 10266 44582 10278 44634
rect 10330 44582 10342 44634
rect 10394 44582 10406 44634
rect 10458 44582 10470 44634
rect 10522 44582 19478 44634
rect 19530 44582 19542 44634
rect 19594 44582 19606 44634
rect 19658 44582 19670 44634
rect 19722 44582 19734 44634
rect 19786 44582 28888 44634
rect 1104 44560 28888 44582
rect 11606 44520 11612 44532
rect 11567 44492 11612 44520
rect 11606 44480 11612 44492
rect 11664 44480 11670 44532
rect 27614 44520 27620 44532
rect 27575 44492 27620 44520
rect 27614 44480 27620 44492
rect 27672 44480 27678 44532
rect 2317 44387 2375 44393
rect 2317 44353 2329 44387
rect 2363 44384 2375 44387
rect 11698 44384 11704 44396
rect 2363 44356 11704 44384
rect 2363 44353 2375 44356
rect 2317 44347 2375 44353
rect 11698 44344 11704 44356
rect 11756 44344 11762 44396
rect 27430 44344 27436 44396
rect 27488 44384 27494 44396
rect 27525 44387 27583 44393
rect 27525 44384 27537 44387
rect 27488 44356 27537 44384
rect 27488 44344 27494 44356
rect 27525 44353 27537 44356
rect 27571 44353 27583 44387
rect 27525 44347 27583 44353
rect 1394 44140 1400 44192
rect 1452 44180 1458 44192
rect 1489 44183 1547 44189
rect 1489 44180 1501 44183
rect 1452 44152 1501 44180
rect 1452 44140 1458 44152
rect 1489 44149 1501 44152
rect 1535 44149 1547 44183
rect 1489 44143 1547 44149
rect 1578 44140 1584 44192
rect 1636 44180 1642 44192
rect 2225 44183 2283 44189
rect 2225 44180 2237 44183
rect 1636 44152 2237 44180
rect 1636 44140 1642 44152
rect 2225 44149 2237 44152
rect 2271 44149 2283 44183
rect 2774 44180 2780 44192
rect 2735 44152 2780 44180
rect 2225 44143 2283 44149
rect 2774 44140 2780 44152
rect 2832 44140 2838 44192
rect 26326 44140 26332 44192
rect 26384 44180 26390 44192
rect 26421 44183 26479 44189
rect 26421 44180 26433 44183
rect 26384 44152 26433 44180
rect 26384 44140 26390 44152
rect 26421 44149 26433 44152
rect 26467 44149 26479 44183
rect 26421 44143 26479 44149
rect 1104 44090 28888 44112
rect 1104 44038 5582 44090
rect 5634 44038 5646 44090
rect 5698 44038 5710 44090
rect 5762 44038 5774 44090
rect 5826 44038 5838 44090
rect 5890 44038 14846 44090
rect 14898 44038 14910 44090
rect 14962 44038 14974 44090
rect 15026 44038 15038 44090
rect 15090 44038 15102 44090
rect 15154 44038 24110 44090
rect 24162 44038 24174 44090
rect 24226 44038 24238 44090
rect 24290 44038 24302 44090
rect 24354 44038 24366 44090
rect 24418 44038 28888 44090
rect 1104 44016 28888 44038
rect 1394 43840 1400 43852
rect 1355 43812 1400 43840
rect 1394 43800 1400 43812
rect 1452 43800 1458 43852
rect 1578 43840 1584 43852
rect 1539 43812 1584 43840
rect 1578 43800 1584 43812
rect 1636 43800 1642 43852
rect 2866 43840 2872 43852
rect 2827 43812 2872 43840
rect 2866 43800 2872 43812
rect 2924 43800 2930 43852
rect 27982 43840 27988 43852
rect 27943 43812 27988 43840
rect 27982 43800 27988 43812
rect 28040 43800 28046 43852
rect 25869 43775 25927 43781
rect 25869 43741 25881 43775
rect 25915 43772 25927 43775
rect 26329 43775 26387 43781
rect 26329 43772 26341 43775
rect 25915 43744 26341 43772
rect 25915 43741 25927 43744
rect 25869 43735 25927 43741
rect 26329 43741 26341 43744
rect 26375 43741 26387 43775
rect 26329 43735 26387 43741
rect 26513 43707 26571 43713
rect 26513 43673 26525 43707
rect 26559 43704 26571 43707
rect 27062 43704 27068 43716
rect 26559 43676 27068 43704
rect 26559 43673 26571 43676
rect 26513 43667 26571 43673
rect 27062 43664 27068 43676
rect 27120 43664 27126 43716
rect 1104 43546 28888 43568
rect 1104 43494 10214 43546
rect 10266 43494 10278 43546
rect 10330 43494 10342 43546
rect 10394 43494 10406 43546
rect 10458 43494 10470 43546
rect 10522 43494 19478 43546
rect 19530 43494 19542 43546
rect 19594 43494 19606 43546
rect 19658 43494 19670 43546
rect 19722 43494 19734 43546
rect 19786 43494 28888 43546
rect 1104 43472 28888 43494
rect 27062 43432 27068 43444
rect 27023 43404 27068 43432
rect 27062 43392 27068 43404
rect 27120 43392 27126 43444
rect 2774 43364 2780 43376
rect 2516 43336 2780 43364
rect 2516 43305 2544 43336
rect 2774 43324 2780 43336
rect 2832 43324 2838 43376
rect 2501 43299 2559 43305
rect 2501 43265 2513 43299
rect 2547 43265 2559 43299
rect 2501 43259 2559 43265
rect 27157 43299 27215 43305
rect 27157 43265 27169 43299
rect 27203 43296 27215 43299
rect 27801 43299 27859 43305
rect 27801 43296 27813 43299
rect 27203 43268 27813 43296
rect 27203 43265 27215 43268
rect 27157 43259 27215 43265
rect 27801 43265 27813 43268
rect 27847 43296 27859 43299
rect 28258 43296 28264 43308
rect 27847 43268 28264 43296
rect 27847 43265 27859 43268
rect 27801 43259 27859 43265
rect 28258 43256 28264 43268
rect 28316 43256 28322 43308
rect 2685 43231 2743 43237
rect 2685 43197 2697 43231
rect 2731 43228 2743 43231
rect 2958 43228 2964 43240
rect 2731 43200 2964 43228
rect 2731 43197 2743 43200
rect 2685 43191 2743 43197
rect 2958 43188 2964 43200
rect 3016 43188 3022 43240
rect 3050 43188 3056 43240
rect 3108 43228 3114 43240
rect 3108 43200 3153 43228
rect 3108 43188 3114 43200
rect 26510 43052 26516 43104
rect 26568 43092 26574 43104
rect 27709 43095 27767 43101
rect 27709 43092 27721 43095
rect 26568 43064 27721 43092
rect 26568 43052 26574 43064
rect 27709 43061 27721 43064
rect 27755 43061 27767 43095
rect 27709 43055 27767 43061
rect 1104 43002 28888 43024
rect 1104 42950 5582 43002
rect 5634 42950 5646 43002
rect 5698 42950 5710 43002
rect 5762 42950 5774 43002
rect 5826 42950 5838 43002
rect 5890 42950 14846 43002
rect 14898 42950 14910 43002
rect 14962 42950 14974 43002
rect 15026 42950 15038 43002
rect 15090 42950 15102 43002
rect 15154 42950 24110 43002
rect 24162 42950 24174 43002
rect 24226 42950 24238 43002
rect 24290 42950 24302 43002
rect 24354 42950 24366 43002
rect 24418 42950 28888 43002
rect 1104 42928 28888 42950
rect 2958 42752 2964 42764
rect 2919 42724 2964 42752
rect 2958 42712 2964 42724
rect 3016 42712 3022 42764
rect 26326 42752 26332 42764
rect 26287 42724 26332 42752
rect 26326 42712 26332 42724
rect 26384 42712 26390 42764
rect 26510 42752 26516 42764
rect 26471 42724 26516 42752
rect 26510 42712 26516 42724
rect 26568 42712 26574 42764
rect 28169 42755 28227 42761
rect 28169 42721 28181 42755
rect 28215 42752 28227 42755
rect 28810 42752 28816 42764
rect 28215 42724 28816 42752
rect 28215 42721 28227 42724
rect 28169 42715 28227 42721
rect 28810 42712 28816 42724
rect 28868 42712 28874 42764
rect 1762 42684 1768 42696
rect 1723 42656 1768 42684
rect 1762 42644 1768 42656
rect 1820 42644 1826 42696
rect 3053 42687 3111 42693
rect 3053 42653 3065 42687
rect 3099 42684 3111 42687
rect 3142 42684 3148 42696
rect 3099 42656 3148 42684
rect 3099 42653 3111 42656
rect 3053 42647 3111 42653
rect 3142 42644 3148 42656
rect 3200 42684 3206 42696
rect 3200 42656 6914 42684
rect 3200 42644 3206 42656
rect 6886 42548 6914 42656
rect 27706 42548 27712 42560
rect 6886 42520 27712 42548
rect 27706 42508 27712 42520
rect 27764 42508 27770 42560
rect 1104 42458 28888 42480
rect 1104 42406 10214 42458
rect 10266 42406 10278 42458
rect 10330 42406 10342 42458
rect 10394 42406 10406 42458
rect 10458 42406 10470 42458
rect 10522 42406 19478 42458
rect 19530 42406 19542 42458
rect 19594 42406 19606 42458
rect 19658 42406 19670 42458
rect 19722 42406 19734 42458
rect 19786 42406 28888 42458
rect 1104 42384 28888 42406
rect 27706 42208 27712 42220
rect 27667 42180 27712 42208
rect 27706 42168 27712 42180
rect 27764 42168 27770 42220
rect 2774 42140 2780 42152
rect 2735 42112 2780 42140
rect 2774 42100 2780 42112
rect 2832 42100 2838 42152
rect 3878 42100 3884 42152
rect 3936 42140 3942 42152
rect 4433 42143 4491 42149
rect 4433 42140 4445 42143
rect 3936 42112 4445 42140
rect 3936 42100 3942 42112
rect 4433 42109 4445 42112
rect 4479 42109 4491 42143
rect 4614 42140 4620 42152
rect 4575 42112 4620 42140
rect 4433 42103 4491 42109
rect 4614 42100 4620 42112
rect 4672 42100 4678 42152
rect 1578 42004 1584 42016
rect 1539 41976 1584 42004
rect 1578 41964 1584 41976
rect 1636 41964 1642 42016
rect 26418 42004 26424 42016
rect 26379 41976 26424 42004
rect 26418 41964 26424 41976
rect 26476 41964 26482 42016
rect 27062 42004 27068 42016
rect 27023 41976 27068 42004
rect 27062 41964 27068 41976
rect 27120 41964 27126 42016
rect 27798 42004 27804 42016
rect 27759 41976 27804 42004
rect 27798 41964 27804 41976
rect 27856 41964 27862 42016
rect 1104 41914 28888 41936
rect 1104 41862 5582 41914
rect 5634 41862 5646 41914
rect 5698 41862 5710 41914
rect 5762 41862 5774 41914
rect 5826 41862 5838 41914
rect 5890 41862 14846 41914
rect 14898 41862 14910 41914
rect 14962 41862 14974 41914
rect 15026 41862 15038 41914
rect 15090 41862 15102 41914
rect 15154 41862 24110 41914
rect 24162 41862 24174 41914
rect 24226 41862 24238 41914
rect 24290 41862 24302 41914
rect 24354 41862 24366 41914
rect 24418 41862 28888 41914
rect 1104 41840 28888 41862
rect 3878 41800 3884 41812
rect 3839 41772 3884 41800
rect 3878 41760 3884 41772
rect 3936 41760 3942 41812
rect 4614 41800 4620 41812
rect 4575 41772 4620 41800
rect 4614 41760 4620 41772
rect 4672 41760 4678 41812
rect 1394 41664 1400 41676
rect 1355 41636 1400 41664
rect 1394 41624 1400 41636
rect 1452 41624 1458 41676
rect 1762 41624 1768 41676
rect 1820 41664 1826 41676
rect 3237 41667 3295 41673
rect 3237 41664 3249 41667
rect 1820 41636 3249 41664
rect 1820 41624 1826 41636
rect 3237 41633 3249 41636
rect 3283 41633 3295 41667
rect 3237 41627 3295 41633
rect 26329 41667 26387 41673
rect 26329 41633 26341 41667
rect 26375 41664 26387 41667
rect 27062 41664 27068 41676
rect 26375 41636 27068 41664
rect 26375 41633 26387 41636
rect 26329 41627 26387 41633
rect 27062 41624 27068 41636
rect 27120 41624 27126 41676
rect 28166 41664 28172 41676
rect 28127 41636 28172 41664
rect 28166 41624 28172 41636
rect 28224 41624 28230 41676
rect 3973 41599 4031 41605
rect 3973 41565 3985 41599
rect 4019 41596 4031 41599
rect 9950 41596 9956 41608
rect 4019 41568 9956 41596
rect 4019 41565 4031 41568
rect 3973 41559 4031 41565
rect 9950 41556 9956 41568
rect 10008 41596 10014 41608
rect 10594 41596 10600 41608
rect 10008 41568 10600 41596
rect 10008 41556 10014 41568
rect 10594 41556 10600 41568
rect 10652 41556 10658 41608
rect 3050 41528 3056 41540
rect 3011 41500 3056 41528
rect 3050 41488 3056 41500
rect 3108 41488 3114 41540
rect 26513 41531 26571 41537
rect 26513 41497 26525 41531
rect 26559 41528 26571 41531
rect 27798 41528 27804 41540
rect 26559 41500 27804 41528
rect 26559 41497 26571 41500
rect 26513 41491 26571 41497
rect 27798 41488 27804 41500
rect 27856 41488 27862 41540
rect 1104 41370 28888 41392
rect 1104 41318 10214 41370
rect 10266 41318 10278 41370
rect 10330 41318 10342 41370
rect 10394 41318 10406 41370
rect 10458 41318 10470 41370
rect 10522 41318 19478 41370
rect 19530 41318 19542 41370
rect 19594 41318 19606 41370
rect 19658 41318 19670 41370
rect 19722 41318 19734 41370
rect 19786 41318 28888 41370
rect 1104 41296 28888 41318
rect 1578 41120 1584 41132
rect 1539 41092 1584 41120
rect 1578 41080 1584 41092
rect 1636 41080 1642 41132
rect 26418 41080 26424 41132
rect 26476 41120 26482 41132
rect 27157 41123 27215 41129
rect 26476 41092 26521 41120
rect 26476 41080 26482 41092
rect 27157 41089 27169 41123
rect 27203 41120 27215 41123
rect 27338 41120 27344 41132
rect 27203 41092 27344 41120
rect 27203 41089 27215 41092
rect 27157 41083 27215 41089
rect 27338 41080 27344 41092
rect 27396 41080 27402 41132
rect 1765 41055 1823 41061
rect 1765 41021 1777 41055
rect 1811 41052 1823 41055
rect 2038 41052 2044 41064
rect 1811 41024 2044 41052
rect 1811 41021 1823 41024
rect 1765 41015 1823 41021
rect 2038 41012 2044 41024
rect 2096 41012 2102 41064
rect 3234 41052 3240 41064
rect 3195 41024 3240 41052
rect 3234 41012 3240 41024
rect 3292 41012 3298 41064
rect 25958 41052 25964 41064
rect 25919 41024 25964 41052
rect 25958 41012 25964 41024
rect 26016 41012 26022 41064
rect 26237 41055 26295 41061
rect 26237 41021 26249 41055
rect 26283 41052 26295 41055
rect 27065 41055 27123 41061
rect 27065 41052 27077 41055
rect 26283 41024 27077 41052
rect 26283 41021 26295 41024
rect 26237 41015 26295 41021
rect 27065 41021 27077 41024
rect 27111 41021 27123 41055
rect 27065 41015 27123 41021
rect 28077 40919 28135 40925
rect 28077 40885 28089 40919
rect 28123 40916 28135 40919
rect 28166 40916 28172 40928
rect 28123 40888 28172 40916
rect 28123 40885 28135 40888
rect 28077 40879 28135 40885
rect 28166 40876 28172 40888
rect 28224 40876 28230 40928
rect 1104 40826 28888 40848
rect 1104 40774 5582 40826
rect 5634 40774 5646 40826
rect 5698 40774 5710 40826
rect 5762 40774 5774 40826
rect 5826 40774 5838 40826
rect 5890 40774 14846 40826
rect 14898 40774 14910 40826
rect 14962 40774 14974 40826
rect 15026 40774 15038 40826
rect 15090 40774 15102 40826
rect 15154 40774 24110 40826
rect 24162 40774 24174 40826
rect 24226 40774 24238 40826
rect 24290 40774 24302 40826
rect 24354 40774 24366 40826
rect 24418 40774 28888 40826
rect 1104 40752 28888 40774
rect 2038 40712 2044 40724
rect 1999 40684 2044 40712
rect 2038 40672 2044 40684
rect 2096 40672 2102 40724
rect 2685 40715 2743 40721
rect 2685 40681 2697 40715
rect 2731 40712 2743 40715
rect 3050 40712 3056 40724
rect 2731 40684 3056 40712
rect 2731 40681 2743 40684
rect 2685 40675 2743 40681
rect 3050 40672 3056 40684
rect 3108 40672 3114 40724
rect 27522 40576 27528 40588
rect 27483 40548 27528 40576
rect 27522 40536 27528 40548
rect 27580 40536 27586 40588
rect 28166 40576 28172 40588
rect 28127 40548 28172 40576
rect 28166 40536 28172 40548
rect 28224 40536 28230 40588
rect 2133 40511 2191 40517
rect 2133 40477 2145 40511
rect 2179 40508 2191 40511
rect 2777 40511 2835 40517
rect 2777 40508 2789 40511
rect 2179 40480 2789 40508
rect 2179 40477 2191 40480
rect 2133 40471 2191 40477
rect 2777 40477 2789 40480
rect 2823 40508 2835 40511
rect 2823 40480 6914 40508
rect 2823 40477 2835 40480
rect 2777 40471 2835 40477
rect 6886 40372 6914 40480
rect 27982 40440 27988 40452
rect 27943 40412 27988 40440
rect 27982 40400 27988 40412
rect 28040 40400 28046 40452
rect 27614 40372 27620 40384
rect 6886 40344 27620 40372
rect 27614 40332 27620 40344
rect 27672 40332 27678 40384
rect 1104 40282 28888 40304
rect 1104 40230 10214 40282
rect 10266 40230 10278 40282
rect 10330 40230 10342 40282
rect 10394 40230 10406 40282
rect 10458 40230 10470 40282
rect 10522 40230 19478 40282
rect 19530 40230 19542 40282
rect 19594 40230 19606 40282
rect 19658 40230 19670 40282
rect 19722 40230 19734 40282
rect 19786 40230 28888 40282
rect 1104 40208 28888 40230
rect 27801 40171 27859 40177
rect 27801 40137 27813 40171
rect 27847 40168 27859 40171
rect 27982 40168 27988 40180
rect 27847 40140 27988 40168
rect 27847 40137 27859 40140
rect 27801 40131 27859 40137
rect 27982 40128 27988 40140
rect 28040 40128 28046 40180
rect 19334 40060 19340 40112
rect 19392 40100 19398 40112
rect 27338 40100 27344 40112
rect 19392 40072 27344 40100
rect 19392 40060 19398 40072
rect 27338 40060 27344 40072
rect 27396 40060 27402 40112
rect 27706 40032 27712 40044
rect 27667 40004 27712 40032
rect 27706 39992 27712 40004
rect 27764 39992 27770 40044
rect 26326 39788 26332 39840
rect 26384 39828 26390 39840
rect 27065 39831 27123 39837
rect 27065 39828 27077 39831
rect 26384 39800 27077 39828
rect 26384 39788 26390 39800
rect 27065 39797 27077 39800
rect 27111 39797 27123 39831
rect 27065 39791 27123 39797
rect 1104 39738 28888 39760
rect 1104 39686 5582 39738
rect 5634 39686 5646 39738
rect 5698 39686 5710 39738
rect 5762 39686 5774 39738
rect 5826 39686 5838 39738
rect 5890 39686 14846 39738
rect 14898 39686 14910 39738
rect 14962 39686 14974 39738
rect 15026 39686 15038 39738
rect 15090 39686 15102 39738
rect 15154 39686 24110 39738
rect 24162 39686 24174 39738
rect 24226 39686 24238 39738
rect 24290 39686 24302 39738
rect 24354 39686 24366 39738
rect 24418 39686 28888 39738
rect 1104 39664 28888 39686
rect 21453 39559 21511 39565
rect 21453 39525 21465 39559
rect 21499 39556 21511 39559
rect 21818 39556 21824 39568
rect 21499 39528 21824 39556
rect 21499 39525 21511 39528
rect 21453 39519 21511 39525
rect 21818 39516 21824 39528
rect 21876 39516 21882 39568
rect 20717 39491 20775 39497
rect 20717 39457 20729 39491
rect 20763 39488 20775 39491
rect 26326 39488 26332 39500
rect 20763 39460 21312 39488
rect 26287 39460 26332 39488
rect 20763 39457 20775 39460
rect 20717 39451 20775 39457
rect 21284 39432 21312 39460
rect 26326 39448 26332 39460
rect 26384 39448 26390 39500
rect 28166 39488 28172 39500
rect 28127 39460 28172 39488
rect 28166 39448 28172 39460
rect 28224 39448 28230 39500
rect 20441 39423 20499 39429
rect 20441 39389 20453 39423
rect 20487 39389 20499 39423
rect 20441 39383 20499 39389
rect 20533 39423 20591 39429
rect 20533 39389 20545 39423
rect 20579 39420 20591 39423
rect 20806 39420 20812 39432
rect 20579 39392 20812 39420
rect 20579 39389 20591 39392
rect 20533 39383 20591 39389
rect 20456 39352 20484 39383
rect 20806 39380 20812 39392
rect 20864 39380 20870 39432
rect 21174 39420 21180 39432
rect 21135 39392 21180 39420
rect 21174 39380 21180 39392
rect 21232 39380 21238 39432
rect 21266 39380 21272 39432
rect 21324 39420 21330 39432
rect 21453 39423 21511 39429
rect 21453 39420 21465 39423
rect 21324 39392 21465 39420
rect 21324 39380 21330 39392
rect 21453 39389 21465 39392
rect 21499 39389 21511 39423
rect 21453 39383 21511 39389
rect 26510 39352 26516 39364
rect 20456 39324 21312 39352
rect 26471 39324 26516 39352
rect 20548 39296 20576 39324
rect 20530 39244 20536 39296
rect 20588 39244 20594 39296
rect 20717 39287 20775 39293
rect 20717 39253 20729 39287
rect 20763 39284 20775 39287
rect 20898 39284 20904 39296
rect 20763 39256 20904 39284
rect 20763 39253 20775 39256
rect 20717 39247 20775 39253
rect 20898 39244 20904 39256
rect 20956 39244 20962 39296
rect 21284 39293 21312 39324
rect 26510 39312 26516 39324
rect 26568 39312 26574 39364
rect 21269 39287 21327 39293
rect 21269 39253 21281 39287
rect 21315 39253 21327 39287
rect 21269 39247 21327 39253
rect 1104 39194 28888 39216
rect 1104 39142 10214 39194
rect 10266 39142 10278 39194
rect 10330 39142 10342 39194
rect 10394 39142 10406 39194
rect 10458 39142 10470 39194
rect 10522 39142 19478 39194
rect 19530 39142 19542 39194
rect 19594 39142 19606 39194
rect 19658 39142 19670 39194
rect 19722 39142 19734 39194
rect 19786 39142 28888 39194
rect 1104 39120 28888 39142
rect 26510 39040 26516 39092
rect 26568 39080 26574 39092
rect 27617 39083 27675 39089
rect 27617 39080 27629 39083
rect 26568 39052 27629 39080
rect 26568 39040 26574 39052
rect 27617 39049 27629 39052
rect 27663 39049 27675 39083
rect 27617 39043 27675 39049
rect 20806 38972 20812 39024
rect 20864 38972 20870 39024
rect 19334 38904 19340 38956
rect 19392 38944 19398 38956
rect 19429 38947 19487 38953
rect 19429 38944 19441 38947
rect 19392 38916 19441 38944
rect 19392 38904 19398 38916
rect 19429 38913 19441 38916
rect 19475 38913 19487 38947
rect 19429 38907 19487 38913
rect 19613 38947 19671 38953
rect 19613 38913 19625 38947
rect 19659 38944 19671 38947
rect 19886 38944 19892 38956
rect 19659 38916 19892 38944
rect 19659 38913 19671 38916
rect 19613 38907 19671 38913
rect 19886 38904 19892 38916
rect 19944 38904 19950 38956
rect 20824 38944 20852 38972
rect 20901 38947 20959 38953
rect 20901 38944 20913 38947
rect 20824 38916 20913 38944
rect 20901 38913 20913 38916
rect 20947 38913 20959 38947
rect 21818 38944 21824 38956
rect 21779 38916 21824 38944
rect 20901 38907 20959 38913
rect 21818 38904 21824 38916
rect 21876 38904 21882 38956
rect 22189 38947 22247 38953
rect 22189 38913 22201 38947
rect 22235 38944 22247 38947
rect 22370 38944 22376 38956
rect 22235 38916 22376 38944
rect 22235 38913 22247 38916
rect 22189 38907 22247 38913
rect 22370 38904 22376 38916
rect 22428 38904 22434 38956
rect 27709 38947 27767 38953
rect 27709 38913 27721 38947
rect 27755 38944 27767 38947
rect 27798 38944 27804 38956
rect 27755 38916 27804 38944
rect 27755 38913 27767 38916
rect 27709 38907 27767 38913
rect 27798 38904 27804 38916
rect 27856 38944 27862 38956
rect 28258 38944 28264 38956
rect 27856 38916 28264 38944
rect 27856 38904 27862 38916
rect 28258 38904 28264 38916
rect 28316 38904 28322 38956
rect 20809 38879 20867 38885
rect 20809 38845 20821 38879
rect 20855 38876 20867 38879
rect 21266 38876 21272 38888
rect 20855 38848 21272 38876
rect 20855 38845 20867 38848
rect 20809 38839 20867 38845
rect 21266 38836 21272 38848
rect 21324 38836 21330 38888
rect 22094 38836 22100 38888
rect 22152 38876 22158 38888
rect 22152 38848 22197 38876
rect 22152 38836 22158 38848
rect 20533 38811 20591 38817
rect 20533 38777 20545 38811
rect 20579 38808 20591 38811
rect 20990 38808 20996 38820
rect 20579 38780 20996 38808
rect 20579 38777 20591 38780
rect 20533 38771 20591 38777
rect 20990 38768 20996 38780
rect 21048 38768 21054 38820
rect 1670 38740 1676 38752
rect 1631 38712 1676 38740
rect 1670 38700 1676 38712
rect 1728 38700 1734 38752
rect 19429 38743 19487 38749
rect 19429 38709 19441 38743
rect 19475 38740 19487 38743
rect 19518 38740 19524 38752
rect 19475 38712 19524 38740
rect 19475 38709 19487 38712
rect 19429 38703 19487 38709
rect 19518 38700 19524 38712
rect 19576 38700 19582 38752
rect 20806 38740 20812 38752
rect 20767 38712 20812 38740
rect 20806 38700 20812 38712
rect 20864 38700 20870 38752
rect 21358 38700 21364 38752
rect 21416 38740 21422 38752
rect 21913 38743 21971 38749
rect 21913 38740 21925 38743
rect 21416 38712 21925 38740
rect 21416 38700 21422 38712
rect 21913 38709 21925 38712
rect 21959 38709 21971 38743
rect 22278 38740 22284 38752
rect 22239 38712 22284 38740
rect 21913 38703 21971 38709
rect 22278 38700 22284 38712
rect 22336 38700 22342 38752
rect 26326 38700 26332 38752
rect 26384 38740 26390 38752
rect 26421 38743 26479 38749
rect 26421 38740 26433 38743
rect 26384 38712 26433 38740
rect 26384 38700 26390 38712
rect 26421 38709 26433 38712
rect 26467 38709 26479 38743
rect 26421 38703 26479 38709
rect 1104 38650 28888 38672
rect 1104 38598 5582 38650
rect 5634 38598 5646 38650
rect 5698 38598 5710 38650
rect 5762 38598 5774 38650
rect 5826 38598 5838 38650
rect 5890 38598 14846 38650
rect 14898 38598 14910 38650
rect 14962 38598 14974 38650
rect 15026 38598 15038 38650
rect 15090 38598 15102 38650
rect 15154 38598 24110 38650
rect 24162 38598 24174 38650
rect 24226 38598 24238 38650
rect 24290 38598 24302 38650
rect 24354 38598 24366 38650
rect 24418 38598 28888 38650
rect 1104 38576 28888 38598
rect 20625 38471 20683 38477
rect 20625 38437 20637 38471
rect 20671 38437 20683 38471
rect 20625 38431 20683 38437
rect 1397 38403 1455 38409
rect 1397 38369 1409 38403
rect 1443 38400 1455 38403
rect 1670 38400 1676 38412
rect 1443 38372 1676 38400
rect 1443 38369 1455 38372
rect 1397 38363 1455 38369
rect 1670 38360 1676 38372
rect 1728 38360 1734 38412
rect 2774 38400 2780 38412
rect 2735 38372 2780 38400
rect 2774 38360 2780 38372
rect 2832 38360 2838 38412
rect 20640 38400 20668 38431
rect 20806 38400 20812 38412
rect 20640 38372 20812 38400
rect 20806 38360 20812 38372
rect 20864 38400 20870 38412
rect 21085 38403 21143 38409
rect 21085 38400 21097 38403
rect 20864 38372 21097 38400
rect 20864 38360 20870 38372
rect 21085 38369 21097 38372
rect 21131 38369 21143 38403
rect 26326 38400 26332 38412
rect 26287 38372 26332 38400
rect 21085 38363 21143 38369
rect 26326 38360 26332 38372
rect 26384 38360 26390 38412
rect 28169 38403 28227 38409
rect 28169 38369 28181 38403
rect 28215 38400 28227 38403
rect 28718 38400 28724 38412
rect 28215 38372 28724 38400
rect 28215 38369 28227 38372
rect 28169 38363 28227 38369
rect 28718 38360 28724 38372
rect 28776 38360 28782 38412
rect 18782 38292 18788 38344
rect 18840 38332 18846 38344
rect 19518 38341 19524 38344
rect 19245 38335 19303 38341
rect 19245 38332 19257 38335
rect 18840 38304 19257 38332
rect 18840 38292 18846 38304
rect 19245 38301 19257 38304
rect 19291 38301 19303 38335
rect 19512 38332 19524 38341
rect 19479 38304 19524 38332
rect 19245 38295 19303 38301
rect 19512 38295 19524 38304
rect 19518 38292 19524 38295
rect 19576 38292 19582 38344
rect 20530 38292 20536 38344
rect 20588 38332 20594 38344
rect 21361 38335 21419 38341
rect 21361 38332 21373 38335
rect 20588 38304 21373 38332
rect 20588 38292 20594 38304
rect 21361 38301 21373 38304
rect 21407 38301 21419 38335
rect 23750 38332 23756 38344
rect 23711 38304 23756 38332
rect 21361 38295 21419 38301
rect 23750 38292 23756 38304
rect 23808 38292 23814 38344
rect 1581 38267 1639 38273
rect 1581 38233 1593 38267
rect 1627 38264 1639 38267
rect 2130 38264 2136 38276
rect 1627 38236 2136 38264
rect 1627 38233 1639 38236
rect 1581 38227 1639 38233
rect 2130 38224 2136 38236
rect 2188 38224 2194 38276
rect 22830 38224 22836 38276
rect 22888 38264 22894 38276
rect 23486 38267 23544 38273
rect 23486 38264 23498 38267
rect 22888 38236 23498 38264
rect 22888 38224 22894 38236
rect 23486 38233 23498 38236
rect 23532 38233 23544 38267
rect 23486 38227 23544 38233
rect 26513 38267 26571 38273
rect 26513 38233 26525 38267
rect 26559 38264 26571 38267
rect 27706 38264 27712 38276
rect 26559 38236 27712 38264
rect 26559 38233 26571 38236
rect 26513 38227 26571 38233
rect 27706 38224 27712 38236
rect 27764 38224 27770 38276
rect 22373 38199 22431 38205
rect 22373 38165 22385 38199
rect 22419 38196 22431 38199
rect 22554 38196 22560 38208
rect 22419 38168 22560 38196
rect 22419 38165 22431 38168
rect 22373 38159 22431 38165
rect 22554 38156 22560 38168
rect 22612 38156 22618 38208
rect 1104 38106 28888 38128
rect 1104 38054 10214 38106
rect 10266 38054 10278 38106
rect 10330 38054 10342 38106
rect 10394 38054 10406 38106
rect 10458 38054 10470 38106
rect 10522 38054 19478 38106
rect 19530 38054 19542 38106
rect 19594 38054 19606 38106
rect 19658 38054 19670 38106
rect 19722 38054 19734 38106
rect 19786 38054 28888 38106
rect 1104 38032 28888 38054
rect 2130 37992 2136 38004
rect 2091 37964 2136 37992
rect 2130 37952 2136 37964
rect 2188 37952 2194 38004
rect 19334 37952 19340 38004
rect 19392 37992 19398 38004
rect 19889 37995 19947 38001
rect 19889 37992 19901 37995
rect 19392 37964 19901 37992
rect 19392 37952 19398 37964
rect 19889 37961 19901 37964
rect 19935 37961 19947 37995
rect 19889 37955 19947 37961
rect 21069 37995 21127 38001
rect 21069 37961 21081 37995
rect 21115 37992 21127 37995
rect 21174 37992 21180 38004
rect 21115 37964 21180 37992
rect 21115 37961 21127 37964
rect 21069 37955 21127 37961
rect 21174 37952 21180 37964
rect 21232 37952 21238 38004
rect 22830 37992 22836 38004
rect 22791 37964 22836 37992
rect 22830 37952 22836 37964
rect 22888 37952 22894 38004
rect 27706 37992 27712 38004
rect 27667 37964 27712 37992
rect 27706 37952 27712 37964
rect 27764 37952 27770 38004
rect 20530 37924 20536 37936
rect 20272 37896 20536 37924
rect 2222 37856 2228 37868
rect 2183 37828 2228 37856
rect 2222 37816 2228 37828
rect 2280 37816 2286 37868
rect 20162 37856 20168 37868
rect 20123 37828 20168 37856
rect 20162 37816 20168 37828
rect 20220 37816 20226 37868
rect 20272 37865 20300 37896
rect 20530 37884 20536 37896
rect 20588 37884 20594 37936
rect 21266 37884 21272 37936
rect 21324 37924 21330 37936
rect 21324 37896 22600 37924
rect 21324 37884 21330 37896
rect 22572 37868 22600 37896
rect 20257 37859 20315 37865
rect 20257 37825 20269 37859
rect 20303 37825 20315 37859
rect 20257 37819 20315 37825
rect 22189 37859 22247 37865
rect 22189 37825 22201 37859
rect 22235 37825 22247 37859
rect 22189 37819 22247 37825
rect 20070 37788 20076 37800
rect 20031 37760 20076 37788
rect 20070 37748 20076 37760
rect 20128 37748 20134 37800
rect 20346 37748 20352 37800
rect 20404 37788 20410 37800
rect 20404 37760 20449 37788
rect 20404 37748 20410 37760
rect 20530 37680 20536 37732
rect 20588 37720 20594 37732
rect 20588 37692 21128 37720
rect 20588 37680 20594 37692
rect 1581 37655 1639 37661
rect 1581 37621 1593 37655
rect 1627 37652 1639 37655
rect 3234 37652 3240 37664
rect 1627 37624 3240 37652
rect 1627 37621 1639 37624
rect 1581 37615 1639 37621
rect 3234 37612 3240 37624
rect 3292 37612 3298 37664
rect 20806 37612 20812 37664
rect 20864 37652 20870 37664
rect 21100 37661 21128 37692
rect 20901 37655 20959 37661
rect 20901 37652 20913 37655
rect 20864 37624 20913 37652
rect 20864 37612 20870 37624
rect 20901 37621 20913 37624
rect 20947 37621 20959 37655
rect 20901 37615 20959 37621
rect 21085 37655 21143 37661
rect 21085 37621 21097 37655
rect 21131 37621 21143 37655
rect 22204 37652 22232 37819
rect 22278 37816 22284 37868
rect 22336 37856 22342 37868
rect 22373 37859 22431 37865
rect 22373 37856 22385 37859
rect 22336 37828 22385 37856
rect 22336 37816 22342 37828
rect 22373 37825 22385 37828
rect 22419 37825 22431 37859
rect 22373 37819 22431 37825
rect 22465 37859 22523 37865
rect 22465 37825 22477 37859
rect 22511 37825 22523 37859
rect 22465 37819 22523 37825
rect 22370 37680 22376 37732
rect 22428 37720 22434 37732
rect 22480 37720 22508 37819
rect 22554 37816 22560 37868
rect 22612 37856 22618 37868
rect 22612 37828 22657 37856
rect 22612 37816 22618 37828
rect 27706 37816 27712 37868
rect 27764 37856 27770 37868
rect 27801 37859 27859 37865
rect 27801 37856 27813 37859
rect 27764 37828 27813 37856
rect 27764 37816 27770 37828
rect 27801 37825 27813 37828
rect 27847 37825 27859 37859
rect 27801 37819 27859 37825
rect 22428 37692 22508 37720
rect 22428 37680 22434 37692
rect 22738 37652 22744 37664
rect 22204 37624 22744 37652
rect 21085 37615 21143 37621
rect 22738 37612 22744 37624
rect 22796 37612 22802 37664
rect 1104 37562 28888 37584
rect 1104 37510 5582 37562
rect 5634 37510 5646 37562
rect 5698 37510 5710 37562
rect 5762 37510 5774 37562
rect 5826 37510 5838 37562
rect 5890 37510 14846 37562
rect 14898 37510 14910 37562
rect 14962 37510 14974 37562
rect 15026 37510 15038 37562
rect 15090 37510 15102 37562
rect 15154 37510 24110 37562
rect 24162 37510 24174 37562
rect 24226 37510 24238 37562
rect 24290 37510 24302 37562
rect 24354 37510 24366 37562
rect 24418 37510 28888 37562
rect 1104 37488 28888 37510
rect 19886 37448 19892 37460
rect 19847 37420 19892 37448
rect 19886 37408 19892 37420
rect 19944 37408 19950 37460
rect 21361 37451 21419 37457
rect 21361 37417 21373 37451
rect 21407 37448 21419 37451
rect 22094 37448 22100 37460
rect 21407 37420 22100 37448
rect 21407 37417 21419 37420
rect 21361 37411 21419 37417
rect 22094 37408 22100 37420
rect 22152 37408 22158 37460
rect 27433 37315 27491 37321
rect 27433 37281 27445 37315
rect 27479 37312 27491 37315
rect 27890 37312 27896 37324
rect 27479 37284 27896 37312
rect 27479 37281 27491 37284
rect 27433 37275 27491 37281
rect 27890 37272 27896 37284
rect 27948 37272 27954 37324
rect 28077 37315 28135 37321
rect 28077 37281 28089 37315
rect 28123 37312 28135 37315
rect 28166 37312 28172 37324
rect 28123 37284 28172 37312
rect 28123 37281 28135 37284
rect 28077 37275 28135 37281
rect 28166 37272 28172 37284
rect 28224 37272 28230 37324
rect 1394 37244 1400 37256
rect 1355 37216 1400 37244
rect 1394 37204 1400 37216
rect 1452 37204 1458 37256
rect 3234 37204 3240 37256
rect 3292 37244 3298 37256
rect 20162 37244 20168 37256
rect 3292 37216 3337 37244
rect 20123 37216 20168 37244
rect 3292 37204 3298 37216
rect 20162 37204 20168 37216
rect 20220 37204 20226 37256
rect 20898 37244 20904 37256
rect 20859 37216 20904 37244
rect 20898 37204 20904 37216
rect 20956 37204 20962 37256
rect 21177 37247 21235 37253
rect 21177 37213 21189 37247
rect 21223 37244 21235 37247
rect 22554 37244 22560 37256
rect 21223 37216 22560 37244
rect 21223 37213 21235 37216
rect 21177 37207 21235 37213
rect 22554 37204 22560 37216
rect 22612 37204 22618 37256
rect 26786 37244 26792 37256
rect 26747 37216 26792 37244
rect 26786 37204 26792 37216
rect 26844 37204 26850 37256
rect 2774 37136 2780 37188
rect 2832 37176 2838 37188
rect 3053 37179 3111 37185
rect 3053 37176 3065 37179
rect 2832 37148 3065 37176
rect 2832 37136 2838 37148
rect 3053 37145 3065 37148
rect 3099 37145 3111 37179
rect 3053 37139 3111 37145
rect 19889 37179 19947 37185
rect 19889 37145 19901 37179
rect 19935 37176 19947 37179
rect 20530 37176 20536 37188
rect 19935 37148 20536 37176
rect 19935 37145 19947 37148
rect 19889 37139 19947 37145
rect 20530 37136 20536 37148
rect 20588 37136 20594 37188
rect 21913 37179 21971 37185
rect 21913 37176 21925 37179
rect 20824 37148 21925 37176
rect 20073 37111 20131 37117
rect 20073 37077 20085 37111
rect 20119 37108 20131 37111
rect 20254 37108 20260 37120
rect 20119 37080 20260 37108
rect 20119 37077 20131 37080
rect 20073 37071 20131 37077
rect 20254 37068 20260 37080
rect 20312 37108 20318 37120
rect 20824 37108 20852 37148
rect 21913 37145 21925 37148
rect 21959 37145 21971 37179
rect 21913 37139 21971 37145
rect 22097 37179 22155 37185
rect 22097 37145 22109 37179
rect 22143 37176 22155 37179
rect 22370 37176 22376 37188
rect 22143 37148 22376 37176
rect 22143 37145 22155 37148
rect 22097 37139 22155 37145
rect 22370 37136 22376 37148
rect 22428 37136 22434 37188
rect 20990 37108 20996 37120
rect 20312 37080 20852 37108
rect 20903 37080 20996 37108
rect 20312 37068 20318 37080
rect 20990 37068 20996 37080
rect 21048 37108 21054 37120
rect 21450 37108 21456 37120
rect 21048 37080 21456 37108
rect 21048 37068 21054 37080
rect 21450 37068 21456 37080
rect 21508 37068 21514 37120
rect 26602 37108 26608 37120
rect 26563 37080 26608 37108
rect 26602 37068 26608 37080
rect 26660 37068 26666 37120
rect 1104 37018 28888 37040
rect 1104 36966 10214 37018
rect 10266 36966 10278 37018
rect 10330 36966 10342 37018
rect 10394 36966 10406 37018
rect 10458 36966 10470 37018
rect 10522 36966 19478 37018
rect 19530 36966 19542 37018
rect 19594 36966 19606 37018
rect 19658 36966 19670 37018
rect 19722 36966 19734 37018
rect 19786 36966 28888 37018
rect 1104 36944 28888 36966
rect 2774 36904 2780 36916
rect 2735 36876 2780 36904
rect 2774 36864 2780 36876
rect 2832 36864 2838 36916
rect 1854 36768 1860 36780
rect 1815 36740 1860 36768
rect 1854 36728 1860 36740
rect 1912 36728 1918 36780
rect 2038 36728 2044 36780
rect 2096 36768 2102 36780
rect 2685 36771 2743 36777
rect 2685 36768 2697 36771
rect 2096 36740 2697 36768
rect 2096 36728 2102 36740
rect 2685 36737 2697 36740
rect 2731 36737 2743 36771
rect 17954 36768 17960 36780
rect 17915 36740 17960 36768
rect 2685 36731 2743 36737
rect 17954 36728 17960 36740
rect 18012 36728 18018 36780
rect 22646 36768 22652 36780
rect 22607 36740 22652 36768
rect 22646 36728 22652 36740
rect 22704 36728 22710 36780
rect 27614 36728 27620 36780
rect 27672 36768 27678 36780
rect 27801 36771 27859 36777
rect 27801 36768 27813 36771
rect 27672 36740 27813 36768
rect 27672 36728 27678 36740
rect 27801 36737 27813 36740
rect 27847 36737 27859 36771
rect 27801 36731 27859 36737
rect 18233 36703 18291 36709
rect 18233 36669 18245 36703
rect 18279 36700 18291 36703
rect 18414 36700 18420 36712
rect 18279 36672 18420 36700
rect 18279 36669 18291 36672
rect 18233 36663 18291 36669
rect 18414 36660 18420 36672
rect 18472 36700 18478 36712
rect 23290 36700 23296 36712
rect 18472 36672 23296 36700
rect 18472 36660 18478 36672
rect 23290 36660 23296 36672
rect 23348 36660 23354 36712
rect 2133 36567 2191 36573
rect 2133 36533 2145 36567
rect 2179 36564 2191 36567
rect 2314 36564 2320 36576
rect 2179 36536 2320 36564
rect 2179 36533 2191 36536
rect 2133 36527 2191 36533
rect 2314 36524 2320 36536
rect 2372 36564 2378 36576
rect 16942 36564 16948 36576
rect 2372 36536 16948 36564
rect 2372 36524 2378 36536
rect 16942 36524 16948 36536
rect 17000 36524 17006 36576
rect 22462 36524 22468 36576
rect 22520 36564 22526 36576
rect 22557 36567 22615 36573
rect 22557 36564 22569 36567
rect 22520 36536 22569 36564
rect 22520 36524 22526 36536
rect 22557 36533 22569 36536
rect 22603 36533 22615 36567
rect 22557 36527 22615 36533
rect 27893 36567 27951 36573
rect 27893 36533 27905 36567
rect 27939 36564 27951 36567
rect 27982 36564 27988 36576
rect 27939 36536 27988 36564
rect 27939 36533 27951 36536
rect 27893 36527 27951 36533
rect 27982 36524 27988 36536
rect 28040 36524 28046 36576
rect 1104 36474 28888 36496
rect 1104 36422 5582 36474
rect 5634 36422 5646 36474
rect 5698 36422 5710 36474
rect 5762 36422 5774 36474
rect 5826 36422 5838 36474
rect 5890 36422 14846 36474
rect 14898 36422 14910 36474
rect 14962 36422 14974 36474
rect 15026 36422 15038 36474
rect 15090 36422 15102 36474
rect 15154 36422 24110 36474
rect 24162 36422 24174 36474
rect 24226 36422 24238 36474
rect 24290 36422 24302 36474
rect 24354 36422 24366 36474
rect 24418 36422 28888 36474
rect 1104 36400 28888 36422
rect 20070 36360 20076 36372
rect 20031 36332 20076 36360
rect 20070 36320 20076 36332
rect 20128 36320 20134 36372
rect 22462 36252 22468 36304
rect 22520 36292 22526 36304
rect 22520 36264 23152 36292
rect 22520 36252 22526 36264
rect 22370 36224 22376 36236
rect 22020 36196 22376 36224
rect 17954 36116 17960 36168
rect 18012 36156 18018 36168
rect 18049 36159 18107 36165
rect 18049 36156 18061 36159
rect 18012 36128 18061 36156
rect 18012 36116 18018 36128
rect 18049 36125 18061 36128
rect 18095 36125 18107 36159
rect 18049 36119 18107 36125
rect 20349 36159 20407 36165
rect 20349 36125 20361 36159
rect 20395 36156 20407 36159
rect 20714 36156 20720 36168
rect 20395 36128 20720 36156
rect 20395 36125 20407 36128
rect 20349 36119 20407 36125
rect 20714 36116 20720 36128
rect 20772 36116 20778 36168
rect 20898 36156 20904 36168
rect 20824 36128 20904 36156
rect 18322 36048 18328 36100
rect 18380 36088 18386 36100
rect 18417 36091 18475 36097
rect 18417 36088 18429 36091
rect 18380 36060 18429 36088
rect 18380 36048 18386 36060
rect 18417 36057 18429 36060
rect 18463 36088 18475 36091
rect 19334 36088 19340 36100
rect 18463 36060 19340 36088
rect 18463 36057 18475 36060
rect 18417 36051 18475 36057
rect 19334 36048 19340 36060
rect 19392 36048 19398 36100
rect 19886 36048 19892 36100
rect 19944 36088 19950 36100
rect 20073 36091 20131 36097
rect 20073 36088 20085 36091
rect 19944 36060 20085 36088
rect 19944 36048 19950 36060
rect 20073 36057 20085 36060
rect 20119 36057 20131 36091
rect 20073 36051 20131 36057
rect 20257 36091 20315 36097
rect 20257 36057 20269 36091
rect 20303 36088 20315 36091
rect 20824 36088 20852 36128
rect 20898 36116 20904 36128
rect 20956 36116 20962 36168
rect 22020 36165 22048 36196
rect 22370 36184 22376 36196
rect 22428 36184 22434 36236
rect 22005 36159 22063 36165
rect 22005 36125 22017 36159
rect 22051 36125 22063 36159
rect 22186 36156 22192 36168
rect 22147 36128 22192 36156
rect 22005 36119 22063 36125
rect 22186 36116 22192 36128
rect 22244 36116 22250 36168
rect 22649 36159 22707 36165
rect 22649 36125 22661 36159
rect 22695 36156 22707 36159
rect 22738 36156 22744 36168
rect 22695 36128 22744 36156
rect 22695 36125 22707 36128
rect 22649 36119 22707 36125
rect 22738 36116 22744 36128
rect 22796 36116 22802 36168
rect 22833 36159 22891 36165
rect 22833 36125 22845 36159
rect 22879 36125 22891 36159
rect 22833 36119 22891 36125
rect 22925 36159 22983 36165
rect 22925 36125 22937 36159
rect 22971 36125 22983 36159
rect 22925 36119 22983 36125
rect 23017 36159 23075 36165
rect 23017 36125 23029 36159
rect 23063 36156 23075 36159
rect 23124 36156 23152 36264
rect 27890 36252 27896 36304
rect 27948 36292 27954 36304
rect 27948 36264 28212 36292
rect 27948 36252 27954 36264
rect 27522 36224 27528 36236
rect 27483 36196 27528 36224
rect 27522 36184 27528 36196
rect 27580 36184 27586 36236
rect 27982 36224 27988 36236
rect 27943 36196 27988 36224
rect 27982 36184 27988 36196
rect 28040 36184 28046 36236
rect 28184 36233 28212 36264
rect 28169 36227 28227 36233
rect 28169 36193 28181 36227
rect 28215 36193 28227 36227
rect 28169 36187 28227 36193
rect 25222 36156 25228 36168
rect 23063 36128 23152 36156
rect 25135 36128 25228 36156
rect 23063 36125 23075 36128
rect 23017 36119 23075 36125
rect 20990 36088 20996 36100
rect 20303 36060 20852 36088
rect 20951 36060 20996 36088
rect 20303 36057 20315 36060
rect 20257 36051 20315 36057
rect 20990 36048 20996 36060
rect 21048 36048 21054 36100
rect 22097 36091 22155 36097
rect 22097 36057 22109 36091
rect 22143 36088 22155 36091
rect 22848 36088 22876 36119
rect 22143 36060 22876 36088
rect 22143 36057 22155 36060
rect 22097 36051 22155 36057
rect 20901 36023 20959 36029
rect 20901 35989 20913 36023
rect 20947 36020 20959 36023
rect 21266 36020 21272 36032
rect 20947 35992 21272 36020
rect 20947 35989 20959 35992
rect 20901 35983 20959 35989
rect 21266 35980 21272 35992
rect 21324 35980 21330 36032
rect 22370 35980 22376 36032
rect 22428 36020 22434 36032
rect 22940 36020 22968 36119
rect 25222 36116 25228 36128
rect 25280 36156 25286 36168
rect 26786 36156 26792 36168
rect 25280 36128 26792 36156
rect 25280 36116 25286 36128
rect 26786 36116 26792 36128
rect 26844 36116 26850 36168
rect 25409 36091 25467 36097
rect 25409 36057 25421 36091
rect 25455 36088 25467 36091
rect 25590 36088 25596 36100
rect 25455 36060 25596 36088
rect 25455 36057 25467 36060
rect 25409 36051 25467 36057
rect 25590 36048 25596 36060
rect 25648 36048 25654 36100
rect 22428 35992 22968 36020
rect 23293 36023 23351 36029
rect 22428 35980 22434 35992
rect 23293 35989 23305 36023
rect 23339 36020 23351 36023
rect 24394 36020 24400 36032
rect 23339 35992 24400 36020
rect 23339 35989 23351 35992
rect 23293 35983 23351 35989
rect 24394 35980 24400 35992
rect 24452 35980 24458 36032
rect 1104 35930 28888 35952
rect 1104 35878 10214 35930
rect 10266 35878 10278 35930
rect 10330 35878 10342 35930
rect 10394 35878 10406 35930
rect 10458 35878 10470 35930
rect 10522 35878 19478 35930
rect 19530 35878 19542 35930
rect 19594 35878 19606 35930
rect 19658 35878 19670 35930
rect 19722 35878 19734 35930
rect 19786 35878 28888 35930
rect 1104 35856 28888 35878
rect 20165 35819 20223 35825
rect 16960 35788 20116 35816
rect 16960 35760 16988 35788
rect 16942 35748 16948 35760
rect 16903 35720 16948 35748
rect 16942 35708 16948 35720
rect 17000 35708 17006 35760
rect 18230 35748 18236 35760
rect 18191 35720 18236 35748
rect 18230 35708 18236 35720
rect 18288 35748 18294 35760
rect 18690 35748 18696 35760
rect 18288 35720 18696 35748
rect 18288 35708 18294 35720
rect 18690 35708 18696 35720
rect 18748 35708 18754 35760
rect 17129 35683 17187 35689
rect 17129 35649 17141 35683
rect 17175 35680 17187 35683
rect 17681 35683 17739 35689
rect 17681 35680 17693 35683
rect 17175 35652 17693 35680
rect 17175 35649 17187 35652
rect 17129 35643 17187 35649
rect 17681 35649 17693 35652
rect 17727 35680 17739 35683
rect 17954 35680 17960 35692
rect 17727 35652 17960 35680
rect 17727 35649 17739 35652
rect 17681 35643 17739 35649
rect 17954 35640 17960 35652
rect 18012 35640 18018 35692
rect 18782 35680 18788 35692
rect 18743 35652 18788 35680
rect 18782 35640 18788 35652
rect 18840 35640 18846 35692
rect 19052 35683 19110 35689
rect 19052 35649 19064 35683
rect 19098 35680 19110 35683
rect 19334 35680 19340 35692
rect 19098 35652 19340 35680
rect 19098 35649 19110 35652
rect 19052 35643 19110 35649
rect 19334 35640 19340 35652
rect 19392 35640 19398 35692
rect 20088 35680 20116 35788
rect 20165 35785 20177 35819
rect 20211 35816 20223 35819
rect 20990 35816 20996 35828
rect 20211 35788 20996 35816
rect 20211 35785 20223 35788
rect 20165 35779 20223 35785
rect 20990 35776 20996 35788
rect 21048 35776 21054 35828
rect 25222 35816 25228 35828
rect 21100 35788 25228 35816
rect 20714 35708 20720 35760
rect 20772 35748 20778 35760
rect 20809 35751 20867 35757
rect 20809 35748 20821 35751
rect 20772 35720 20821 35748
rect 20772 35708 20778 35720
rect 20809 35717 20821 35720
rect 20855 35717 20867 35751
rect 21100 35748 21128 35788
rect 25222 35776 25228 35788
rect 25280 35776 25286 35828
rect 20809 35711 20867 35717
rect 20916 35720 21128 35748
rect 20916 35680 20944 35720
rect 21542 35708 21548 35760
rect 21600 35748 21606 35760
rect 21600 35720 24348 35748
rect 21600 35708 21606 35720
rect 21082 35689 21088 35692
rect 20088 35652 20944 35680
rect 21053 35683 21088 35689
rect 21053 35649 21065 35683
rect 21053 35643 21088 35649
rect 21082 35640 21088 35643
rect 21140 35640 21146 35692
rect 21177 35683 21235 35689
rect 21177 35649 21189 35683
rect 21223 35680 21235 35683
rect 22462 35680 22468 35692
rect 21223 35652 22324 35680
rect 22423 35652 22468 35680
rect 21223 35649 21235 35652
rect 21177 35643 21235 35649
rect 22296 35624 22324 35652
rect 22462 35640 22468 35652
rect 22520 35640 22526 35692
rect 24320 35680 24348 35720
rect 24394 35708 24400 35760
rect 24452 35757 24458 35760
rect 24452 35748 24464 35757
rect 24452 35720 24497 35748
rect 24452 35711 24464 35720
rect 24452 35708 24458 35711
rect 25590 35680 25596 35692
rect 24320 35652 24808 35680
rect 25551 35652 25596 35680
rect 21275 35615 21333 35621
rect 21275 35581 21287 35615
rect 21321 35581 21333 35615
rect 21275 35575 21333 35581
rect 21284 35544 21312 35575
rect 22278 35572 22284 35624
rect 22336 35612 22342 35624
rect 22373 35615 22431 35621
rect 22373 35612 22385 35615
rect 22336 35584 22385 35612
rect 22336 35572 22342 35584
rect 22373 35581 22385 35584
rect 22419 35581 22431 35615
rect 22373 35575 22431 35581
rect 24673 35615 24731 35621
rect 24673 35581 24685 35615
rect 24719 35581 24731 35615
rect 24780 35612 24808 35652
rect 25590 35640 25596 35652
rect 25648 35640 25654 35692
rect 27246 35640 27252 35692
rect 27304 35680 27310 35692
rect 27617 35683 27675 35689
rect 27617 35680 27629 35683
rect 27304 35652 27629 35680
rect 27304 35640 27310 35652
rect 27617 35649 27629 35652
rect 27663 35649 27675 35683
rect 27617 35643 27675 35649
rect 25866 35612 25872 35624
rect 24780 35584 25872 35612
rect 24673 35575 24731 35581
rect 22646 35544 22652 35556
rect 21284 35516 22652 35544
rect 22646 35504 22652 35516
rect 22704 35544 22710 35556
rect 22704 35516 23336 35544
rect 22704 35504 22710 35516
rect 23308 35488 23336 35516
rect 24688 35488 24716 35575
rect 25866 35572 25872 35584
rect 25924 35612 25930 35624
rect 26145 35615 26203 35621
rect 26145 35612 26157 35615
rect 25924 35584 26157 35612
rect 25924 35572 25930 35584
rect 26145 35581 26157 35584
rect 26191 35612 26203 35615
rect 27706 35612 27712 35624
rect 26191 35584 27712 35612
rect 26191 35581 26203 35584
rect 26145 35575 26203 35581
rect 27706 35572 27712 35584
rect 27764 35572 27770 35624
rect 1394 35436 1400 35488
rect 1452 35476 1458 35488
rect 1489 35479 1547 35485
rect 1489 35476 1501 35479
rect 1452 35448 1501 35476
rect 1452 35436 1458 35448
rect 1489 35445 1501 35448
rect 1535 35445 1547 35479
rect 1489 35439 1547 35445
rect 2317 35479 2375 35485
rect 2317 35445 2329 35479
rect 2363 35476 2375 35479
rect 3602 35476 3608 35488
rect 2363 35448 3608 35476
rect 2363 35445 2375 35448
rect 2317 35439 2375 35445
rect 3602 35436 3608 35448
rect 3660 35436 3666 35488
rect 11698 35436 11704 35488
rect 11756 35476 11762 35488
rect 21542 35476 21548 35488
rect 11756 35448 21548 35476
rect 11756 35436 11762 35448
rect 21542 35436 21548 35448
rect 21600 35436 21606 35488
rect 22833 35479 22891 35485
rect 22833 35445 22845 35479
rect 22879 35476 22891 35479
rect 23106 35476 23112 35488
rect 22879 35448 23112 35476
rect 22879 35445 22891 35448
rect 22833 35439 22891 35445
rect 23106 35436 23112 35448
rect 23164 35436 23170 35488
rect 23290 35476 23296 35488
rect 23251 35448 23296 35476
rect 23290 35436 23296 35448
rect 23348 35436 23354 35488
rect 23474 35436 23480 35488
rect 23532 35476 23538 35488
rect 23750 35476 23756 35488
rect 23532 35448 23756 35476
rect 23532 35436 23538 35448
rect 23750 35436 23756 35448
rect 23808 35476 23814 35488
rect 24670 35476 24676 35488
rect 23808 35448 24676 35476
rect 23808 35436 23814 35448
rect 24670 35436 24676 35448
rect 24728 35436 24734 35488
rect 26326 35436 26332 35488
rect 26384 35476 26390 35488
rect 26973 35479 27031 35485
rect 26973 35476 26985 35479
rect 26384 35448 26985 35476
rect 26384 35436 26390 35448
rect 26973 35445 26985 35448
rect 27019 35445 27031 35479
rect 26973 35439 27031 35445
rect 1104 35386 28888 35408
rect 1104 35334 5582 35386
rect 5634 35334 5646 35386
rect 5698 35334 5710 35386
rect 5762 35334 5774 35386
rect 5826 35334 5838 35386
rect 5890 35334 14846 35386
rect 14898 35334 14910 35386
rect 14962 35334 14974 35386
rect 15026 35334 15038 35386
rect 15090 35334 15102 35386
rect 15154 35334 24110 35386
rect 24162 35334 24174 35386
rect 24226 35334 24238 35386
rect 24290 35334 24302 35386
rect 24354 35334 24366 35386
rect 24418 35334 28888 35386
rect 1104 35312 28888 35334
rect 20625 35275 20683 35281
rect 20625 35241 20637 35275
rect 20671 35272 20683 35275
rect 20714 35272 20720 35284
rect 20671 35244 20720 35272
rect 20671 35241 20683 35244
rect 20625 35235 20683 35241
rect 20640 35204 20668 35235
rect 20714 35232 20720 35244
rect 20772 35272 20778 35284
rect 21174 35272 21180 35284
rect 20772 35244 21180 35272
rect 20772 35232 20778 35244
rect 21174 35232 21180 35244
rect 21232 35232 21238 35284
rect 22186 35232 22192 35284
rect 22244 35272 22250 35284
rect 22465 35275 22523 35281
rect 22465 35272 22477 35275
rect 22244 35244 22477 35272
rect 22244 35232 22250 35244
rect 22465 35241 22477 35244
rect 22511 35241 22523 35275
rect 27246 35272 27252 35284
rect 27207 35244 27252 35272
rect 22465 35235 22523 35241
rect 27246 35232 27252 35244
rect 27304 35232 27310 35284
rect 22741 35207 22799 35213
rect 22741 35204 22753 35207
rect 19812 35176 20668 35204
rect 22066 35176 22753 35204
rect 1394 35136 1400 35148
rect 1355 35108 1400 35136
rect 1394 35096 1400 35108
rect 1452 35096 1458 35148
rect 2774 35136 2780 35148
rect 2735 35108 2780 35136
rect 2774 35096 2780 35108
rect 2832 35096 2838 35148
rect 18322 35136 18328 35148
rect 18283 35108 18328 35136
rect 18322 35096 18328 35108
rect 18380 35096 18386 35148
rect 17954 35028 17960 35080
rect 18012 35068 18018 35080
rect 19812 35077 19840 35176
rect 20257 35139 20315 35145
rect 20257 35105 20269 35139
rect 20303 35136 20315 35139
rect 20990 35136 20996 35148
rect 20303 35108 20996 35136
rect 20303 35105 20315 35108
rect 20257 35099 20315 35105
rect 20990 35096 20996 35108
rect 21048 35096 21054 35148
rect 22066 35136 22094 35176
rect 22741 35173 22753 35176
rect 22787 35204 22799 35207
rect 23566 35204 23572 35216
rect 22787 35176 23572 35204
rect 22787 35173 22799 35176
rect 22741 35167 22799 35173
rect 23566 35164 23572 35176
rect 23624 35164 23630 35216
rect 21468 35108 22094 35136
rect 21468 35077 21496 35108
rect 22554 35096 22560 35148
rect 22612 35136 22618 35148
rect 22833 35139 22891 35145
rect 22612 35108 22784 35136
rect 22612 35096 22618 35108
rect 18049 35071 18107 35077
rect 18049 35068 18061 35071
rect 18012 35040 18061 35068
rect 18012 35028 18018 35040
rect 18049 35037 18061 35040
rect 18095 35037 18107 35071
rect 18049 35031 18107 35037
rect 19613 35071 19671 35077
rect 19613 35037 19625 35071
rect 19659 35037 19671 35071
rect 19613 35031 19671 35037
rect 19797 35071 19855 35077
rect 19797 35037 19809 35071
rect 19843 35037 19855 35071
rect 19797 35031 19855 35037
rect 20441 35071 20499 35077
rect 20441 35037 20453 35071
rect 20487 35068 20499 35071
rect 21453 35071 21511 35077
rect 21453 35068 21465 35071
rect 20487 35040 21465 35068
rect 20487 35037 20499 35040
rect 20441 35031 20499 35037
rect 21453 35037 21465 35040
rect 21499 35037 21511 35071
rect 21453 35031 21511 35037
rect 22649 35071 22707 35077
rect 22649 35037 22661 35071
rect 22695 35037 22707 35071
rect 22756 35068 22784 35108
rect 22833 35105 22845 35139
rect 22879 35136 22891 35139
rect 23658 35136 23664 35148
rect 22879 35108 23664 35136
rect 22879 35105 22891 35108
rect 22833 35099 22891 35105
rect 23658 35096 23664 35108
rect 23716 35096 23722 35148
rect 24670 35096 24676 35148
rect 24728 35136 24734 35148
rect 25869 35139 25927 35145
rect 25869 35136 25881 35139
rect 24728 35108 25881 35136
rect 24728 35096 24734 35108
rect 25869 35105 25881 35108
rect 25915 35105 25927 35139
rect 25869 35099 25927 35105
rect 22925 35071 22983 35077
rect 22925 35068 22937 35071
rect 22756 35040 22937 35068
rect 22649 35031 22707 35037
rect 22925 35037 22937 35040
rect 22971 35037 22983 35071
rect 23106 35068 23112 35080
rect 23067 35040 23112 35068
rect 22925 35031 22983 35037
rect 1581 35003 1639 35009
rect 1581 35000 1593 35003
rect 1504 34972 1593 35000
rect 1504 34944 1532 34972
rect 1581 34969 1593 34972
rect 1627 34969 1639 35003
rect 19628 35000 19656 35031
rect 19628 34972 21220 35000
rect 1581 34963 1639 34969
rect 1486 34892 1492 34944
rect 1544 34892 1550 34944
rect 19705 34935 19763 34941
rect 19705 34901 19717 34935
rect 19751 34932 19763 34935
rect 19886 34932 19892 34944
rect 19751 34904 19892 34932
rect 19751 34901 19763 34904
rect 19705 34895 19763 34901
rect 19886 34892 19892 34904
rect 19944 34892 19950 34944
rect 21082 34932 21088 34944
rect 21043 34904 21088 34932
rect 21082 34892 21088 34904
rect 21140 34892 21146 34944
rect 21192 34932 21220 34972
rect 21266 34960 21272 35012
rect 21324 35000 21330 35012
rect 21324 34972 21369 35000
rect 21324 34960 21330 34972
rect 22094 34932 22100 34944
rect 21192 34904 22100 34932
rect 22094 34892 22100 34904
rect 22152 34932 22158 34944
rect 22664 34932 22692 35031
rect 23106 35028 23112 35040
rect 23164 35028 23170 35080
rect 25317 35071 25375 35077
rect 25317 35037 25329 35071
rect 25363 35037 25375 35071
rect 25317 35031 25375 35037
rect 26136 35071 26194 35077
rect 26136 35037 26148 35071
rect 26182 35068 26194 35071
rect 26602 35068 26608 35080
rect 26182 35040 26608 35068
rect 26182 35037 26194 35040
rect 26136 35031 26194 35037
rect 24949 35003 25007 35009
rect 24949 34969 24961 35003
rect 24995 34969 25007 35003
rect 25332 35000 25360 35031
rect 26602 35028 26608 35040
rect 26660 35028 26666 35080
rect 27706 35068 27712 35080
rect 27667 35040 27712 35068
rect 27706 35028 27712 35040
rect 27764 35028 27770 35080
rect 25590 35000 25596 35012
rect 25332 34972 25596 35000
rect 24949 34963 25007 34969
rect 22152 34904 22692 34932
rect 22152 34892 22158 34904
rect 24854 34892 24860 34944
rect 24912 34932 24918 34944
rect 24964 34932 24992 34963
rect 25590 34960 25596 34972
rect 25648 35000 25654 35012
rect 27724 35000 27752 35028
rect 25648 34972 27752 35000
rect 25648 34960 25654 34972
rect 27798 34960 27804 35012
rect 27856 35000 27862 35012
rect 27985 35003 28043 35009
rect 27985 35000 27997 35003
rect 27856 34972 27997 35000
rect 27856 34960 27862 34972
rect 27985 34969 27997 34972
rect 28031 35000 28043 35003
rect 28810 35000 28816 35012
rect 28031 34972 28816 35000
rect 28031 34969 28043 34972
rect 27985 34963 28043 34969
rect 28810 34960 28816 34972
rect 28868 34960 28874 35012
rect 27430 34932 27436 34944
rect 24912 34904 27436 34932
rect 24912 34892 24918 34904
rect 27430 34892 27436 34904
rect 27488 34892 27494 34944
rect 1104 34842 28888 34864
rect 1104 34790 10214 34842
rect 10266 34790 10278 34842
rect 10330 34790 10342 34842
rect 10394 34790 10406 34842
rect 10458 34790 10470 34842
rect 10522 34790 19478 34842
rect 19530 34790 19542 34842
rect 19594 34790 19606 34842
rect 19658 34790 19670 34842
rect 19722 34790 19734 34842
rect 19786 34790 28888 34842
rect 1104 34768 28888 34790
rect 2222 34688 2228 34740
rect 2280 34728 2286 34740
rect 2280 34700 27476 34728
rect 2280 34688 2286 34700
rect 27448 34672 27476 34700
rect 1762 34660 1768 34672
rect 1723 34632 1768 34660
rect 1762 34620 1768 34632
rect 1820 34620 1826 34672
rect 1946 34620 1952 34672
rect 2004 34660 2010 34672
rect 18601 34663 18659 34669
rect 18601 34660 18613 34663
rect 2004 34632 18613 34660
rect 2004 34620 2010 34632
rect 18601 34629 18613 34632
rect 18647 34660 18659 34663
rect 20438 34660 20444 34672
rect 18647 34632 20444 34660
rect 18647 34629 18659 34632
rect 18601 34623 18659 34629
rect 20438 34620 20444 34632
rect 20496 34620 20502 34672
rect 20990 34660 20996 34672
rect 20951 34632 20996 34660
rect 20990 34620 20996 34632
rect 21048 34620 21054 34672
rect 21082 34620 21088 34672
rect 21140 34669 21146 34672
rect 21140 34663 21169 34669
rect 21157 34629 21169 34663
rect 21140 34623 21169 34629
rect 21140 34620 21146 34623
rect 21266 34620 21272 34672
rect 21324 34660 21330 34672
rect 21324 34632 22048 34660
rect 21324 34620 21330 34632
rect 3602 34552 3608 34604
rect 3660 34592 3666 34604
rect 3660 34564 3705 34592
rect 3660 34552 3666 34564
rect 17954 34552 17960 34604
rect 18012 34592 18018 34604
rect 18049 34595 18107 34601
rect 18049 34592 18061 34595
rect 18012 34564 18061 34592
rect 18012 34552 18018 34564
rect 18049 34561 18061 34564
rect 18095 34561 18107 34595
rect 18049 34555 18107 34561
rect 19886 34552 19892 34604
rect 19944 34592 19950 34604
rect 20809 34595 20867 34601
rect 19944 34564 20760 34592
rect 19944 34552 19950 34564
rect 3418 34524 3424 34536
rect 3379 34496 3424 34524
rect 3418 34484 3424 34496
rect 3476 34484 3482 34536
rect 20622 34524 20628 34536
rect 20583 34496 20628 34524
rect 20622 34484 20628 34496
rect 20680 34484 20686 34536
rect 20732 34456 20760 34564
rect 20809 34561 20821 34595
rect 20855 34561 20867 34595
rect 20809 34555 20867 34561
rect 20824 34524 20852 34555
rect 20898 34552 20904 34604
rect 20956 34592 20962 34604
rect 22020 34601 22048 34632
rect 24670 34620 24676 34672
rect 24728 34660 24734 34672
rect 27430 34660 27436 34672
rect 24728 34632 26464 34660
rect 27343 34632 27436 34660
rect 24728 34620 24734 34632
rect 22005 34595 22063 34601
rect 20956 34564 21001 34592
rect 21100 34564 21864 34592
rect 20956 34552 20962 34564
rect 21100 34524 21128 34564
rect 21269 34527 21327 34533
rect 21269 34524 21281 34527
rect 20824 34496 21128 34524
rect 21192 34496 21281 34524
rect 21192 34456 21220 34496
rect 21269 34493 21281 34496
rect 21315 34493 21327 34527
rect 21269 34487 21327 34493
rect 21836 34465 21864 34564
rect 22005 34561 22017 34595
rect 22051 34561 22063 34595
rect 22186 34592 22192 34604
rect 22147 34564 22192 34592
rect 22005 34555 22063 34561
rect 22186 34552 22192 34564
rect 22244 34552 22250 34604
rect 26165 34595 26223 34601
rect 26165 34561 26177 34595
rect 26211 34592 26223 34595
rect 26326 34592 26332 34604
rect 26211 34564 26332 34592
rect 26211 34561 26223 34564
rect 26165 34555 26223 34561
rect 26326 34552 26332 34564
rect 26384 34552 26390 34604
rect 26436 34601 26464 34632
rect 27430 34620 27436 34632
rect 27488 34620 27494 34672
rect 26421 34595 26479 34601
rect 26421 34561 26433 34595
rect 26467 34561 26479 34595
rect 26421 34555 26479 34561
rect 27065 34595 27123 34601
rect 27065 34561 27077 34595
rect 27111 34592 27123 34595
rect 27706 34592 27712 34604
rect 27111 34564 27712 34592
rect 27111 34561 27123 34564
rect 27065 34555 27123 34561
rect 27706 34552 27712 34564
rect 27764 34552 27770 34604
rect 20732 34428 21220 34456
rect 21821 34459 21879 34465
rect 21821 34425 21833 34459
rect 21867 34425 21879 34459
rect 21821 34419 21879 34425
rect 22189 34391 22247 34397
rect 22189 34357 22201 34391
rect 22235 34388 22247 34391
rect 23290 34388 23296 34400
rect 22235 34360 23296 34388
rect 22235 34357 22247 34360
rect 22189 34351 22247 34357
rect 23290 34348 23296 34360
rect 23348 34348 23354 34400
rect 25038 34388 25044 34400
rect 24999 34360 25044 34388
rect 25038 34348 25044 34360
rect 25096 34348 25102 34400
rect 1104 34298 28888 34320
rect 1104 34246 5582 34298
rect 5634 34246 5646 34298
rect 5698 34246 5710 34298
rect 5762 34246 5774 34298
rect 5826 34246 5838 34298
rect 5890 34246 14846 34298
rect 14898 34246 14910 34298
rect 14962 34246 14974 34298
rect 15026 34246 15038 34298
rect 15090 34246 15102 34298
rect 15154 34246 24110 34298
rect 24162 34246 24174 34298
rect 24226 34246 24238 34298
rect 24290 34246 24302 34298
rect 24354 34246 24366 34298
rect 24418 34246 28888 34298
rect 1104 34224 28888 34246
rect 2593 34187 2651 34193
rect 2593 34153 2605 34187
rect 2639 34184 2651 34187
rect 3418 34184 3424 34196
rect 2639 34156 3424 34184
rect 2639 34153 2651 34156
rect 2593 34147 2651 34153
rect 3418 34144 3424 34156
rect 3476 34144 3482 34196
rect 20162 34184 20168 34196
rect 20123 34156 20168 34184
rect 20162 34144 20168 34156
rect 20220 34144 20226 34196
rect 20364 34156 20668 34184
rect 20364 34116 20392 34156
rect 19444 34088 20392 34116
rect 2682 33980 2688 33992
rect 2643 33952 2688 33980
rect 2682 33940 2688 33952
rect 2740 33940 2746 33992
rect 19444 33989 19472 34088
rect 20438 34076 20444 34128
rect 20496 34076 20502 34128
rect 20456 33989 20484 34076
rect 19245 33983 19303 33989
rect 19245 33949 19257 33983
rect 19291 33949 19303 33983
rect 19245 33943 19303 33949
rect 19429 33983 19487 33989
rect 19429 33949 19441 33983
rect 19475 33949 19487 33983
rect 19429 33943 19487 33949
rect 20349 33983 20407 33989
rect 20349 33949 20361 33983
rect 20395 33949 20407 33983
rect 20349 33943 20407 33949
rect 20441 33983 20499 33989
rect 20441 33949 20453 33983
rect 20487 33949 20499 33983
rect 20441 33943 20499 33949
rect 19260 33912 19288 33943
rect 19886 33912 19892 33924
rect 19260 33884 19892 33912
rect 19886 33872 19892 33884
rect 19944 33872 19950 33924
rect 19337 33847 19395 33853
rect 19337 33813 19349 33847
rect 19383 33844 19395 33847
rect 20162 33844 20168 33856
rect 19383 33816 20168 33844
rect 19383 33813 19395 33816
rect 19337 33807 19395 33813
rect 20162 33804 20168 33816
rect 20220 33804 20226 33856
rect 20364 33844 20392 33943
rect 20530 33912 20536 33924
rect 20491 33884 20536 33912
rect 20530 33872 20536 33884
rect 20588 33872 20594 33924
rect 20640 33912 20668 34156
rect 20898 34144 20904 34196
rect 20956 34184 20962 34196
rect 21361 34187 21419 34193
rect 21361 34184 21373 34187
rect 20956 34156 21373 34184
rect 20956 34144 20962 34156
rect 21361 34153 21373 34156
rect 21407 34153 21419 34187
rect 21361 34147 21419 34153
rect 23477 34187 23535 34193
rect 23477 34153 23489 34187
rect 23523 34184 23535 34187
rect 23566 34184 23572 34196
rect 23523 34156 23572 34184
rect 23523 34153 23535 34156
rect 23477 34147 23535 34153
rect 23566 34144 23572 34156
rect 23624 34144 23630 34196
rect 23661 34187 23719 34193
rect 23661 34153 23673 34187
rect 23707 34153 23719 34187
rect 23661 34147 23719 34153
rect 23290 34076 23296 34128
rect 23348 34116 23354 34128
rect 23676 34116 23704 34147
rect 23348 34088 23704 34116
rect 23348 34076 23354 34088
rect 21082 34008 21088 34060
rect 21140 34048 21146 34060
rect 21266 34048 21272 34060
rect 21140 34020 21272 34048
rect 21140 34008 21146 34020
rect 21266 34008 21272 34020
rect 21324 34008 21330 34060
rect 21453 34051 21511 34057
rect 21453 34017 21465 34051
rect 21499 34048 21511 34051
rect 22186 34048 22192 34060
rect 21499 34020 22192 34048
rect 21499 34017 21511 34020
rect 21453 34011 21511 34017
rect 22186 34008 22192 34020
rect 22244 34048 22250 34060
rect 22646 34048 22652 34060
rect 22244 34020 22652 34048
rect 22244 34008 22250 34020
rect 22646 34008 22652 34020
rect 22704 34048 22710 34060
rect 24397 34051 24455 34057
rect 24397 34048 24409 34051
rect 22704 34020 24409 34048
rect 22704 34008 22710 34020
rect 24397 34017 24409 34020
rect 24443 34017 24455 34051
rect 27522 34048 27528 34060
rect 27483 34020 27528 34048
rect 24397 34011 24455 34017
rect 27522 34008 27528 34020
rect 27580 34008 27586 34060
rect 28166 34048 28172 34060
rect 28127 34020 28172 34048
rect 28166 34008 28172 34020
rect 28224 34008 28230 34060
rect 20714 33940 20720 33992
rect 20772 33980 20778 33992
rect 21545 33983 21603 33989
rect 20772 33952 20817 33980
rect 20772 33940 20778 33952
rect 21545 33949 21557 33983
rect 21591 33980 21603 33983
rect 21818 33980 21824 33992
rect 21591 33952 21824 33980
rect 21591 33949 21603 33952
rect 21545 33943 21603 33949
rect 21818 33940 21824 33952
rect 21876 33980 21882 33992
rect 22462 33980 22468 33992
rect 21876 33952 22468 33980
rect 21876 33940 21882 33952
rect 22462 33940 22468 33952
rect 22520 33980 22526 33992
rect 23382 33980 23388 33992
rect 22520 33952 23388 33980
rect 22520 33940 22526 33952
rect 23382 33940 23388 33952
rect 23440 33940 23446 33992
rect 25038 33980 25044 33992
rect 23676 33952 25044 33980
rect 23676 33912 23704 33952
rect 25038 33940 25044 33952
rect 25096 33980 25102 33992
rect 25777 33983 25835 33989
rect 25777 33980 25789 33983
rect 25096 33952 25789 33980
rect 25096 33940 25102 33952
rect 25777 33949 25789 33952
rect 25823 33949 25835 33983
rect 25777 33943 25835 33949
rect 23842 33912 23848 33924
rect 20640 33884 23704 33912
rect 23803 33884 23848 33912
rect 23842 33872 23848 33884
rect 23900 33872 23906 33924
rect 24578 33912 24584 33924
rect 24320 33884 24584 33912
rect 20898 33844 20904 33856
rect 20364 33816 20904 33844
rect 20898 33804 20904 33816
rect 20956 33804 20962 33856
rect 23645 33847 23703 33853
rect 23645 33813 23657 33847
rect 23691 33844 23703 33847
rect 24320 33844 24348 33884
rect 24578 33872 24584 33884
rect 24636 33872 24642 33924
rect 27154 33872 27160 33924
rect 27212 33912 27218 33924
rect 27985 33915 28043 33921
rect 27985 33912 27997 33915
rect 27212 33884 27997 33912
rect 27212 33872 27218 33884
rect 27985 33881 27997 33884
rect 28031 33881 28043 33915
rect 27985 33875 28043 33881
rect 25130 33844 25136 33856
rect 23691 33816 24348 33844
rect 25091 33816 25136 33844
rect 23691 33813 23703 33816
rect 23645 33807 23703 33813
rect 25130 33804 25136 33816
rect 25188 33804 25194 33856
rect 1104 33754 28888 33776
rect 1104 33702 10214 33754
rect 10266 33702 10278 33754
rect 10330 33702 10342 33754
rect 10394 33702 10406 33754
rect 10458 33702 10470 33754
rect 10522 33702 19478 33754
rect 19530 33702 19542 33754
rect 19594 33702 19606 33754
rect 19658 33702 19670 33754
rect 19722 33702 19734 33754
rect 19786 33702 28888 33754
rect 1104 33680 28888 33702
rect 19337 33643 19395 33649
rect 19337 33609 19349 33643
rect 19383 33609 19395 33643
rect 24578 33640 24584 33652
rect 24539 33612 24584 33640
rect 19337 33603 19395 33609
rect 18322 33572 18328 33584
rect 17972 33544 18328 33572
rect 17972 33513 18000 33544
rect 18322 33532 18328 33544
rect 18380 33572 18386 33584
rect 18782 33572 18788 33584
rect 18380 33544 18788 33572
rect 18380 33532 18386 33544
rect 18782 33532 18788 33544
rect 18840 33532 18846 33584
rect 19352 33572 19380 33603
rect 24578 33600 24584 33612
rect 24636 33600 24642 33652
rect 27154 33640 27160 33652
rect 27115 33612 27160 33640
rect 27154 33600 27160 33612
rect 27212 33600 27218 33652
rect 22646 33572 22652 33584
rect 19352 33544 20116 33572
rect 22607 33544 22652 33572
rect 17957 33507 18015 33513
rect 17957 33473 17969 33507
rect 18003 33473 18015 33507
rect 17957 33467 18015 33473
rect 18224 33507 18282 33513
rect 18224 33473 18236 33507
rect 18270 33504 18282 33507
rect 19797 33507 19855 33513
rect 18270 33476 19748 33504
rect 18270 33473 18282 33476
rect 18224 33467 18282 33473
rect 19720 33436 19748 33476
rect 19797 33473 19809 33507
rect 19843 33504 19855 33507
rect 19886 33504 19892 33516
rect 19843 33476 19892 33504
rect 19843 33473 19855 33476
rect 19797 33467 19855 33473
rect 19886 33464 19892 33476
rect 19944 33464 19950 33516
rect 20088 33513 20116 33544
rect 22646 33532 22652 33544
rect 22704 33532 22710 33584
rect 23468 33575 23526 33581
rect 23468 33541 23480 33575
rect 23514 33572 23526 33575
rect 23566 33572 23572 33584
rect 23514 33544 23572 33572
rect 23514 33541 23526 33544
rect 23468 33535 23526 33541
rect 23566 33532 23572 33544
rect 23624 33532 23630 33584
rect 27614 33532 27620 33584
rect 27672 33572 27678 33584
rect 27890 33572 27896 33584
rect 27672 33544 27896 33572
rect 27672 33532 27678 33544
rect 27890 33532 27896 33544
rect 27948 33572 27954 33584
rect 27985 33575 28043 33581
rect 27985 33572 27997 33575
rect 27948 33544 27997 33572
rect 27948 33532 27954 33544
rect 27985 33541 27997 33544
rect 28031 33541 28043 33575
rect 27985 33535 28043 33541
rect 20073 33507 20131 33513
rect 20073 33473 20085 33507
rect 20119 33473 20131 33507
rect 20073 33467 20131 33473
rect 20162 33464 20168 33516
rect 20220 33504 20226 33516
rect 25130 33504 25136 33516
rect 20220 33476 20265 33504
rect 23124 33476 25136 33504
rect 20220 33464 20226 33476
rect 23124 33436 23152 33476
rect 25130 33464 25136 33476
rect 25188 33464 25194 33516
rect 26970 33464 26976 33516
rect 27028 33504 27034 33516
rect 27065 33507 27123 33513
rect 27065 33504 27077 33507
rect 27028 33476 27077 33504
rect 27028 33464 27034 33476
rect 27065 33473 27077 33476
rect 27111 33473 27123 33507
rect 27706 33504 27712 33516
rect 27667 33476 27712 33504
rect 27065 33467 27123 33473
rect 27706 33464 27712 33476
rect 27764 33464 27770 33516
rect 19720 33408 23152 33436
rect 23201 33439 23259 33445
rect 23201 33405 23213 33439
rect 23247 33405 23259 33439
rect 23201 33399 23259 33405
rect 19889 33371 19947 33377
rect 19889 33337 19901 33371
rect 19935 33368 19947 33371
rect 20530 33368 20536 33380
rect 19935 33340 20536 33368
rect 19935 33337 19947 33340
rect 19889 33331 19947 33337
rect 20530 33328 20536 33340
rect 20588 33328 20594 33380
rect 19978 33260 19984 33312
rect 20036 33300 20042 33312
rect 20349 33303 20407 33309
rect 20349 33300 20361 33303
rect 20036 33272 20361 33300
rect 20036 33260 20042 33272
rect 20349 33269 20361 33272
rect 20395 33269 20407 33303
rect 20349 33263 20407 33269
rect 22557 33303 22615 33309
rect 22557 33269 22569 33303
rect 22603 33300 22615 33303
rect 22738 33300 22744 33312
rect 22603 33272 22744 33300
rect 22603 33269 22615 33272
rect 22557 33263 22615 33269
rect 22738 33260 22744 33272
rect 22796 33260 22802 33312
rect 23216 33300 23244 33399
rect 23474 33300 23480 33312
rect 23216 33272 23480 33300
rect 23474 33260 23480 33272
rect 23532 33260 23538 33312
rect 25777 33303 25835 33309
rect 25777 33269 25789 33303
rect 25823 33300 25835 33303
rect 26234 33300 26240 33312
rect 25823 33272 26240 33300
rect 25823 33269 25835 33272
rect 25777 33263 25835 33269
rect 26234 33260 26240 33272
rect 26292 33260 26298 33312
rect 26326 33260 26332 33312
rect 26384 33300 26390 33312
rect 26421 33303 26479 33309
rect 26421 33300 26433 33303
rect 26384 33272 26433 33300
rect 26384 33260 26390 33272
rect 26421 33269 26433 33272
rect 26467 33269 26479 33303
rect 26421 33263 26479 33269
rect 1104 33210 28888 33232
rect 1104 33158 5582 33210
rect 5634 33158 5646 33210
rect 5698 33158 5710 33210
rect 5762 33158 5774 33210
rect 5826 33158 5838 33210
rect 5890 33158 14846 33210
rect 14898 33158 14910 33210
rect 14962 33158 14974 33210
rect 15026 33158 15038 33210
rect 15090 33158 15102 33210
rect 15154 33158 24110 33210
rect 24162 33158 24174 33210
rect 24226 33158 24238 33210
rect 24290 33158 24302 33210
rect 24354 33158 24366 33210
rect 24418 33158 28888 33210
rect 1104 33136 28888 33158
rect 19334 33056 19340 33108
rect 19392 33096 19398 33108
rect 19705 33099 19763 33105
rect 19705 33096 19717 33099
rect 19392 33068 19717 33096
rect 19392 33056 19398 33068
rect 19705 33065 19717 33068
rect 19751 33065 19763 33099
rect 19705 33059 19763 33065
rect 23017 33099 23075 33105
rect 23017 33065 23029 33099
rect 23063 33096 23075 33099
rect 23566 33096 23572 33108
rect 23063 33068 23572 33096
rect 23063 33065 23075 33068
rect 23017 33059 23075 33065
rect 23566 33056 23572 33068
rect 23624 33056 23630 33108
rect 19978 33028 19984 33040
rect 19939 33000 19984 33028
rect 19978 32988 19984 33000
rect 20036 32988 20042 33040
rect 20073 33031 20131 33037
rect 20073 32997 20085 33031
rect 20119 33028 20131 33031
rect 20622 33028 20628 33040
rect 20119 33000 20628 33028
rect 20119 32997 20131 33000
rect 20073 32991 20131 32997
rect 20622 32988 20628 33000
rect 20680 32988 20686 33040
rect 22370 32988 22376 33040
rect 22428 33028 22434 33040
rect 23477 33031 23535 33037
rect 22428 33000 22692 33028
rect 22428 32988 22434 33000
rect 19889 32895 19947 32901
rect 19889 32861 19901 32895
rect 19935 32861 19947 32895
rect 19889 32855 19947 32861
rect 19904 32824 19932 32855
rect 20162 32852 20168 32904
rect 20220 32892 20226 32904
rect 20349 32895 20407 32901
rect 20220 32864 20265 32892
rect 20220 32852 20226 32864
rect 20349 32861 20361 32895
rect 20395 32892 20407 32895
rect 21726 32892 21732 32904
rect 20395 32864 21732 32892
rect 20395 32861 20407 32864
rect 20349 32855 20407 32861
rect 21726 32852 21732 32864
rect 21784 32852 21790 32904
rect 22370 32892 22376 32904
rect 22331 32864 22376 32892
rect 22370 32852 22376 32864
rect 22428 32852 22434 32904
rect 22554 32892 22560 32904
rect 22515 32864 22560 32892
rect 22554 32852 22560 32864
rect 22612 32852 22618 32904
rect 22664 32901 22692 33000
rect 23477 32997 23489 33031
rect 23523 33028 23535 33031
rect 23658 33028 23664 33040
rect 23523 33000 23664 33028
rect 23523 32997 23535 33000
rect 23477 32991 23535 32997
rect 23658 32988 23664 33000
rect 23716 32988 23722 33040
rect 26970 33028 26976 33040
rect 25884 33000 26976 33028
rect 22649 32895 22707 32901
rect 22649 32861 22661 32895
rect 22695 32861 22707 32895
rect 22649 32855 22707 32861
rect 22738 32852 22744 32904
rect 22796 32892 22802 32904
rect 25884 32901 25912 33000
rect 26970 32988 26976 33000
rect 27028 32988 27034 33040
rect 26326 32960 26332 32972
rect 26287 32932 26332 32960
rect 26326 32920 26332 32932
rect 26384 32920 26390 32972
rect 28074 32960 28080 32972
rect 28035 32932 28080 32960
rect 28074 32920 28080 32932
rect 28132 32920 28138 32972
rect 23753 32895 23811 32901
rect 23753 32892 23765 32895
rect 22796 32864 23765 32892
rect 22796 32852 22802 32864
rect 23753 32861 23765 32864
rect 23799 32861 23811 32895
rect 23753 32855 23811 32861
rect 25869 32895 25927 32901
rect 25869 32861 25881 32895
rect 25915 32861 25927 32895
rect 25869 32855 25927 32861
rect 20714 32824 20720 32836
rect 19904 32796 20720 32824
rect 20714 32784 20720 32796
rect 20772 32784 20778 32836
rect 23382 32784 23388 32836
rect 23440 32824 23446 32836
rect 23477 32827 23535 32833
rect 23477 32824 23489 32827
rect 23440 32796 23489 32824
rect 23440 32784 23446 32796
rect 23477 32793 23489 32796
rect 23523 32793 23535 32827
rect 23477 32787 23535 32793
rect 25777 32827 25835 32833
rect 25777 32793 25789 32827
rect 25823 32824 25835 32827
rect 26513 32827 26571 32833
rect 26513 32824 26525 32827
rect 25823 32796 26525 32824
rect 25823 32793 25835 32796
rect 25777 32787 25835 32793
rect 26513 32793 26525 32796
rect 26559 32793 26571 32827
rect 26513 32787 26571 32793
rect 23658 32756 23664 32768
rect 23619 32728 23664 32756
rect 23658 32716 23664 32728
rect 23716 32716 23722 32768
rect 1104 32666 28888 32688
rect 1104 32614 10214 32666
rect 10266 32614 10278 32666
rect 10330 32614 10342 32666
rect 10394 32614 10406 32666
rect 10458 32614 10470 32666
rect 10522 32614 19478 32666
rect 19530 32614 19542 32666
rect 19594 32614 19606 32666
rect 19658 32614 19670 32666
rect 19722 32614 19734 32666
rect 19786 32614 28888 32666
rect 1104 32592 28888 32614
rect 20162 32512 20168 32564
rect 20220 32552 20226 32564
rect 20809 32555 20867 32561
rect 20809 32552 20821 32555
rect 20220 32524 20821 32552
rect 20220 32512 20226 32524
rect 20809 32521 20821 32524
rect 20855 32521 20867 32555
rect 20809 32515 20867 32521
rect 18322 32484 18328 32496
rect 16684 32456 18328 32484
rect 16684 32425 16712 32456
rect 18322 32444 18328 32456
rect 18380 32444 18386 32496
rect 20254 32444 20260 32496
rect 20312 32484 20318 32496
rect 20349 32487 20407 32493
rect 20349 32484 20361 32487
rect 20312 32456 20361 32484
rect 20312 32444 20318 32456
rect 20349 32453 20361 32456
rect 20395 32484 20407 32487
rect 26237 32487 26295 32493
rect 20395 32456 21220 32484
rect 20395 32453 20407 32456
rect 20349 32447 20407 32453
rect 21192 32428 21220 32456
rect 26237 32453 26249 32487
rect 26283 32484 26295 32487
rect 27801 32487 27859 32493
rect 27801 32484 27813 32487
rect 26283 32456 27813 32484
rect 26283 32453 26295 32456
rect 26237 32447 26295 32453
rect 27801 32453 27813 32456
rect 27847 32453 27859 32487
rect 27801 32447 27859 32453
rect 16669 32419 16727 32425
rect 16669 32385 16681 32419
rect 16715 32385 16727 32419
rect 16669 32379 16727 32385
rect 16758 32376 16764 32428
rect 16816 32416 16822 32428
rect 16925 32419 16983 32425
rect 16925 32416 16937 32419
rect 16816 32388 16937 32416
rect 16816 32376 16822 32388
rect 16925 32385 16937 32388
rect 16971 32385 16983 32419
rect 16925 32379 16983 32385
rect 19981 32419 20039 32425
rect 19981 32385 19993 32419
rect 20027 32385 20039 32419
rect 19981 32379 20039 32385
rect 19996 32348 20024 32379
rect 20070 32376 20076 32428
rect 20128 32416 20134 32428
rect 20165 32419 20223 32425
rect 20165 32416 20177 32419
rect 20128 32388 20177 32416
rect 20128 32376 20134 32388
rect 20165 32385 20177 32388
rect 20211 32385 20223 32419
rect 20165 32379 20223 32385
rect 20993 32419 21051 32425
rect 20993 32385 21005 32419
rect 21039 32416 21051 32419
rect 21082 32416 21088 32428
rect 21039 32388 21088 32416
rect 21039 32385 21051 32388
rect 20993 32379 21051 32385
rect 21082 32376 21088 32388
rect 21140 32376 21146 32428
rect 21174 32376 21180 32428
rect 21232 32416 21238 32428
rect 21232 32388 21277 32416
rect 21232 32376 21238 32388
rect 21542 32376 21548 32428
rect 21600 32416 21606 32428
rect 22005 32419 22063 32425
rect 22005 32416 22017 32419
rect 21600 32388 22017 32416
rect 21600 32376 21606 32388
rect 22005 32385 22017 32388
rect 22051 32416 22063 32419
rect 23658 32416 23664 32428
rect 22051 32388 23664 32416
rect 22051 32385 22063 32388
rect 22005 32379 22063 32385
rect 23658 32376 23664 32388
rect 23716 32376 23722 32428
rect 26970 32416 26976 32428
rect 26931 32388 26976 32416
rect 26970 32376 26976 32388
rect 27028 32376 27034 32428
rect 27709 32419 27767 32425
rect 27709 32385 27721 32419
rect 27755 32416 27767 32419
rect 28442 32416 28448 32428
rect 27755 32388 28448 32416
rect 27755 32385 27767 32388
rect 27709 32379 27767 32385
rect 28442 32376 28448 32388
rect 28500 32376 28506 32428
rect 20714 32348 20720 32360
rect 19996 32320 20720 32348
rect 20714 32308 20720 32320
rect 20772 32308 20778 32360
rect 21266 32308 21272 32360
rect 21324 32348 21330 32360
rect 22097 32351 22155 32357
rect 22097 32348 22109 32351
rect 21324 32320 22109 32348
rect 21324 32308 21330 32320
rect 22097 32317 22109 32320
rect 22143 32348 22155 32351
rect 22462 32348 22468 32360
rect 22143 32320 22468 32348
rect 22143 32317 22155 32320
rect 22097 32311 22155 32317
rect 22462 32308 22468 32320
rect 22520 32348 22526 32360
rect 22738 32348 22744 32360
rect 22520 32320 22744 32348
rect 22520 32308 22526 32320
rect 22738 32308 22744 32320
rect 22796 32308 22802 32360
rect 25958 32348 25964 32360
rect 25919 32320 25964 32348
rect 25958 32308 25964 32320
rect 26016 32308 26022 32360
rect 26234 32308 26240 32360
rect 26292 32348 26298 32360
rect 26421 32351 26479 32357
rect 26421 32348 26433 32351
rect 26292 32320 26433 32348
rect 26292 32308 26298 32320
rect 26421 32317 26433 32320
rect 26467 32317 26479 32351
rect 26421 32311 26479 32317
rect 1394 32172 1400 32224
rect 1452 32212 1458 32224
rect 1489 32215 1547 32221
rect 1489 32212 1501 32215
rect 1452 32184 1501 32212
rect 1452 32172 1458 32184
rect 1489 32181 1501 32184
rect 1535 32181 1547 32215
rect 1489 32175 1547 32181
rect 17678 32172 17684 32224
rect 17736 32212 17742 32224
rect 18049 32215 18107 32221
rect 18049 32212 18061 32215
rect 17736 32184 18061 32212
rect 17736 32172 17742 32184
rect 18049 32181 18061 32184
rect 18095 32181 18107 32215
rect 18049 32175 18107 32181
rect 19610 32172 19616 32224
rect 19668 32212 19674 32224
rect 21726 32212 21732 32224
rect 19668 32184 21732 32212
rect 19668 32172 19674 32184
rect 21726 32172 21732 32184
rect 21784 32172 21790 32224
rect 22278 32212 22284 32224
rect 22239 32184 22284 32212
rect 22278 32172 22284 32184
rect 22336 32172 22342 32224
rect 27065 32215 27123 32221
rect 27065 32181 27077 32215
rect 27111 32212 27123 32215
rect 27246 32212 27252 32224
rect 27111 32184 27252 32212
rect 27111 32181 27123 32184
rect 27065 32175 27123 32181
rect 27246 32172 27252 32184
rect 27304 32172 27310 32224
rect 1104 32122 28888 32144
rect 1104 32070 5582 32122
rect 5634 32070 5646 32122
rect 5698 32070 5710 32122
rect 5762 32070 5774 32122
rect 5826 32070 5838 32122
rect 5890 32070 14846 32122
rect 14898 32070 14910 32122
rect 14962 32070 14974 32122
rect 15026 32070 15038 32122
rect 15090 32070 15102 32122
rect 15154 32070 24110 32122
rect 24162 32070 24174 32122
rect 24226 32070 24238 32122
rect 24290 32070 24302 32122
rect 24354 32070 24366 32122
rect 24418 32070 28888 32122
rect 1104 32048 28888 32070
rect 3326 31968 3332 32020
rect 3384 32008 3390 32020
rect 22281 32011 22339 32017
rect 3384 31980 6914 32008
rect 3384 31968 3390 31980
rect 6886 31940 6914 31980
rect 12406 31980 22094 32008
rect 12406 31940 12434 31980
rect 6886 31912 12434 31940
rect 16669 31943 16727 31949
rect 16669 31909 16681 31943
rect 16715 31940 16727 31943
rect 16758 31940 16764 31952
rect 16715 31912 16764 31940
rect 16715 31909 16727 31912
rect 16669 31903 16727 31909
rect 16758 31900 16764 31912
rect 16816 31900 16822 31952
rect 20257 31943 20315 31949
rect 20257 31909 20269 31943
rect 20303 31940 20315 31943
rect 20530 31940 20536 31952
rect 20303 31912 20536 31940
rect 20303 31909 20315 31912
rect 20257 31903 20315 31909
rect 20530 31900 20536 31912
rect 20588 31900 20594 31952
rect 22066 31940 22094 31980
rect 22281 31977 22293 32011
rect 22327 32008 22339 32011
rect 22554 32008 22560 32020
rect 22327 31980 22560 32008
rect 22327 31977 22339 31980
rect 22281 31971 22339 31977
rect 22554 31968 22560 31980
rect 22612 31968 22618 32020
rect 23477 32011 23535 32017
rect 23477 31977 23489 32011
rect 23523 32008 23535 32011
rect 23658 32008 23664 32020
rect 23523 31980 23664 32008
rect 23523 31977 23535 31980
rect 23477 31971 23535 31977
rect 23658 31968 23664 31980
rect 23716 31968 23722 32020
rect 22066 31912 25636 31940
rect 1394 31872 1400 31884
rect 1355 31844 1400 31872
rect 1394 31832 1400 31844
rect 1452 31832 1458 31884
rect 1854 31872 1860 31884
rect 1815 31844 1860 31872
rect 1854 31832 1860 31844
rect 1912 31832 1918 31884
rect 17586 31872 17592 31884
rect 17547 31844 17592 31872
rect 17586 31832 17592 31844
rect 17644 31832 17650 31884
rect 17773 31875 17831 31881
rect 17773 31841 17785 31875
rect 17819 31872 17831 31875
rect 17862 31872 17868 31884
rect 17819 31844 17868 31872
rect 17819 31841 17831 31844
rect 17773 31835 17831 31841
rect 17862 31832 17868 31844
rect 17920 31832 17926 31884
rect 20714 31872 20720 31884
rect 19444 31844 20720 31872
rect 16485 31807 16543 31813
rect 16485 31773 16497 31807
rect 16531 31804 16543 31807
rect 16850 31804 16856 31816
rect 16531 31776 16856 31804
rect 16531 31773 16543 31776
rect 16485 31767 16543 31773
rect 16850 31764 16856 31776
rect 16908 31764 16914 31816
rect 19444 31813 19472 31844
rect 20714 31832 20720 31844
rect 20772 31832 20778 31884
rect 22373 31875 22431 31881
rect 22373 31841 22385 31875
rect 22419 31872 22431 31875
rect 22646 31872 22652 31884
rect 22419 31844 22652 31872
rect 22419 31841 22431 31844
rect 22373 31835 22431 31841
rect 22646 31832 22652 31844
rect 22704 31872 22710 31884
rect 23106 31872 23112 31884
rect 22704 31844 23112 31872
rect 22704 31832 22710 31844
rect 23106 31832 23112 31844
rect 23164 31832 23170 31884
rect 25608 31881 25636 31912
rect 25593 31875 25651 31881
rect 25593 31841 25605 31875
rect 25639 31841 25651 31875
rect 27246 31872 27252 31884
rect 27207 31844 27252 31872
rect 25593 31835 25651 31841
rect 27246 31832 27252 31844
rect 27304 31832 27310 31884
rect 18693 31807 18751 31813
rect 18693 31773 18705 31807
rect 18739 31804 18751 31807
rect 19245 31807 19303 31813
rect 19245 31804 19257 31807
rect 18739 31776 19257 31804
rect 18739 31773 18751 31776
rect 18693 31767 18751 31773
rect 19245 31773 19257 31776
rect 19291 31773 19303 31807
rect 19245 31767 19303 31773
rect 19429 31807 19487 31813
rect 19429 31773 19441 31807
rect 19475 31773 19487 31807
rect 19610 31804 19616 31816
rect 19571 31776 19616 31804
rect 19429 31767 19487 31773
rect 19610 31764 19616 31776
rect 19668 31764 19674 31816
rect 20070 31804 20076 31816
rect 20031 31776 20076 31804
rect 20070 31764 20076 31776
rect 20128 31764 20134 31816
rect 20257 31807 20315 31813
rect 20257 31773 20269 31807
rect 20303 31804 20315 31807
rect 20438 31804 20444 31816
rect 20303 31776 20444 31804
rect 20303 31773 20315 31776
rect 20257 31767 20315 31773
rect 20438 31764 20444 31776
rect 20496 31764 20502 31816
rect 21174 31764 21180 31816
rect 21232 31804 21238 31816
rect 21913 31807 21971 31813
rect 21913 31804 21925 31807
rect 21232 31776 21925 31804
rect 21232 31764 21238 31776
rect 21913 31773 21925 31776
rect 21959 31773 21971 31807
rect 22094 31804 22100 31816
rect 22055 31776 22100 31804
rect 21913 31767 21971 31773
rect 22094 31764 22100 31776
rect 22152 31764 22158 31816
rect 22247 31807 22305 31813
rect 22247 31782 22259 31807
rect 22204 31773 22259 31782
rect 22293 31804 22305 31807
rect 22462 31804 22468 31816
rect 22293 31773 22324 31804
rect 22423 31776 22468 31804
rect 22204 31754 22324 31773
rect 22462 31764 22468 31776
rect 22520 31764 22526 31816
rect 23569 31807 23627 31813
rect 23569 31773 23581 31807
rect 23615 31804 23627 31807
rect 23842 31804 23848 31816
rect 23615 31776 23848 31804
rect 23615 31773 23627 31776
rect 23569 31767 23627 31773
rect 23842 31764 23848 31776
rect 23900 31764 23906 31816
rect 27430 31764 27436 31816
rect 27488 31804 27494 31816
rect 28077 31807 28135 31813
rect 27488 31776 27533 31804
rect 27488 31764 27494 31776
rect 28077 31773 28089 31807
rect 28123 31804 28135 31807
rect 28166 31804 28172 31816
rect 28123 31776 28172 31804
rect 28123 31773 28135 31776
rect 28077 31767 28135 31773
rect 28166 31764 28172 31776
rect 28224 31764 28230 31816
rect 22204 31748 22291 31754
rect 1578 31736 1584 31748
rect 1539 31708 1584 31736
rect 1578 31696 1584 31708
rect 1636 31696 1642 31748
rect 22186 31696 22192 31748
rect 22244 31726 22291 31748
rect 22244 31696 22250 31726
rect 17126 31668 17132 31680
rect 17087 31640 17132 31668
rect 17126 31628 17132 31640
rect 17184 31628 17190 31680
rect 17497 31671 17555 31677
rect 17497 31637 17509 31671
rect 17543 31668 17555 31671
rect 17586 31668 17592 31680
rect 17543 31640 17592 31668
rect 17543 31637 17555 31640
rect 17497 31631 17555 31637
rect 17586 31628 17592 31640
rect 17644 31628 17650 31680
rect 18506 31668 18512 31680
rect 18467 31640 18512 31668
rect 18506 31628 18512 31640
rect 18564 31628 18570 31680
rect 1104 31578 28888 31600
rect 1104 31526 10214 31578
rect 10266 31526 10278 31578
rect 10330 31526 10342 31578
rect 10394 31526 10406 31578
rect 10458 31526 10470 31578
rect 10522 31526 19478 31578
rect 19530 31526 19542 31578
rect 19594 31526 19606 31578
rect 19658 31526 19670 31578
rect 19722 31526 19734 31578
rect 19786 31526 28888 31578
rect 1104 31504 28888 31526
rect 1578 31424 1584 31476
rect 1636 31464 1642 31476
rect 1857 31467 1915 31473
rect 1857 31464 1869 31467
rect 1636 31436 1869 31464
rect 1636 31424 1642 31436
rect 1857 31433 1869 31436
rect 1903 31433 1915 31467
rect 16850 31464 16856 31476
rect 16811 31436 16856 31464
rect 1857 31427 1915 31433
rect 16850 31424 16856 31436
rect 16908 31424 16914 31476
rect 23842 31424 23848 31476
rect 23900 31464 23906 31476
rect 23937 31467 23995 31473
rect 23937 31464 23949 31467
rect 23900 31436 23949 31464
rect 23900 31424 23906 31436
rect 23937 31433 23949 31436
rect 23983 31433 23995 31467
rect 23937 31427 23995 31433
rect 17126 31356 17132 31408
rect 17184 31396 17190 31408
rect 18506 31405 18512 31408
rect 17221 31399 17279 31405
rect 17221 31396 17233 31399
rect 17184 31368 17233 31396
rect 17184 31356 17190 31368
rect 17221 31365 17233 31368
rect 17267 31365 17279 31399
rect 17221 31359 17279 31365
rect 18500 31359 18512 31405
rect 18564 31396 18570 31408
rect 18564 31368 18600 31396
rect 18506 31356 18512 31359
rect 18564 31356 18570 31368
rect 1949 31331 2007 31337
rect 1949 31297 1961 31331
rect 1995 31328 2007 31331
rect 2222 31328 2228 31340
rect 1995 31300 2228 31328
rect 1995 31297 2007 31300
rect 1949 31291 2007 31297
rect 2222 31288 2228 31300
rect 2280 31288 2286 31340
rect 17037 31331 17095 31337
rect 17037 31297 17049 31331
rect 17083 31328 17095 31331
rect 17083 31300 17264 31328
rect 17083 31297 17095 31300
rect 17037 31291 17095 31297
rect 17236 31272 17264 31300
rect 18322 31288 18328 31340
rect 18380 31288 18386 31340
rect 20162 31288 20168 31340
rect 20220 31328 20226 31340
rect 21821 31331 21879 31337
rect 21821 31328 21833 31331
rect 20220 31300 21833 31328
rect 20220 31288 20226 31300
rect 21821 31297 21833 31300
rect 21867 31297 21879 31331
rect 21821 31291 21879 31297
rect 22005 31331 22063 31337
rect 22005 31297 22017 31331
rect 22051 31328 22063 31331
rect 22094 31328 22100 31340
rect 22051 31300 22100 31328
rect 22051 31297 22063 31300
rect 22005 31291 22063 31297
rect 22094 31288 22100 31300
rect 22152 31288 22158 31340
rect 22462 31288 22468 31340
rect 22520 31328 22526 31340
rect 22813 31331 22871 31337
rect 22813 31328 22825 31331
rect 22520 31300 22825 31328
rect 22520 31288 22526 31300
rect 22813 31297 22825 31300
rect 22859 31297 22871 31331
rect 27798 31328 27804 31340
rect 27759 31300 27804 31328
rect 22813 31291 22871 31297
rect 27798 31288 27804 31300
rect 27856 31288 27862 31340
rect 17218 31220 17224 31272
rect 17276 31220 17282 31272
rect 18233 31263 18291 31269
rect 18233 31229 18245 31263
rect 18279 31260 18291 31263
rect 18340 31260 18368 31288
rect 18279 31232 18368 31260
rect 22557 31263 22615 31269
rect 18279 31229 18291 31232
rect 18233 31223 18291 31229
rect 22557 31229 22569 31263
rect 22603 31229 22615 31263
rect 22557 31223 22615 31229
rect 18248 31124 18276 31223
rect 19242 31124 19248 31136
rect 18248 31096 19248 31124
rect 19242 31084 19248 31096
rect 19300 31084 19306 31136
rect 19613 31127 19671 31133
rect 19613 31093 19625 31127
rect 19659 31124 19671 31127
rect 20070 31124 20076 31136
rect 19659 31096 20076 31124
rect 19659 31093 19671 31096
rect 19613 31087 19671 31093
rect 20070 31084 20076 31096
rect 20128 31084 20134 31136
rect 21821 31127 21879 31133
rect 21821 31093 21833 31127
rect 21867 31124 21879 31127
rect 21910 31124 21916 31136
rect 21867 31096 21916 31124
rect 21867 31093 21879 31096
rect 21821 31087 21879 31093
rect 21910 31084 21916 31096
rect 21968 31084 21974 31136
rect 22572 31124 22600 31223
rect 23474 31124 23480 31136
rect 22572 31096 23480 31124
rect 23474 31084 23480 31096
rect 23532 31084 23538 31136
rect 27893 31127 27951 31133
rect 27893 31093 27905 31127
rect 27939 31124 27951 31127
rect 27982 31124 27988 31136
rect 27939 31096 27988 31124
rect 27939 31093 27951 31096
rect 27893 31087 27951 31093
rect 27982 31084 27988 31096
rect 28040 31084 28046 31136
rect 1104 31034 28888 31056
rect 1104 30982 5582 31034
rect 5634 30982 5646 31034
rect 5698 30982 5710 31034
rect 5762 30982 5774 31034
rect 5826 30982 5838 31034
rect 5890 30982 14846 31034
rect 14898 30982 14910 31034
rect 14962 30982 14974 31034
rect 15026 30982 15038 31034
rect 15090 30982 15102 31034
rect 15154 30982 24110 31034
rect 24162 30982 24174 31034
rect 24226 30982 24238 31034
rect 24290 30982 24302 31034
rect 24354 30982 24366 31034
rect 24418 30982 28888 31034
rect 1104 30960 28888 30982
rect 21269 30923 21327 30929
rect 21269 30889 21281 30923
rect 21315 30920 21327 30923
rect 21358 30920 21364 30932
rect 21315 30892 21364 30920
rect 21315 30889 21327 30892
rect 21269 30883 21327 30889
rect 21358 30880 21364 30892
rect 21416 30880 21422 30932
rect 19334 30812 19340 30864
rect 19392 30852 19398 30864
rect 20165 30855 20223 30861
rect 20165 30852 20177 30855
rect 19392 30824 20177 30852
rect 19392 30812 19398 30824
rect 20165 30821 20177 30824
rect 20211 30821 20223 30855
rect 20165 30815 20223 30821
rect 20898 30812 20904 30864
rect 20956 30852 20962 30864
rect 22005 30855 22063 30861
rect 22005 30852 22017 30855
rect 20956 30824 22017 30852
rect 20956 30812 20962 30824
rect 22005 30821 22017 30824
rect 22051 30852 22063 30855
rect 22094 30852 22100 30864
rect 22051 30824 22100 30852
rect 22051 30821 22063 30824
rect 22005 30815 22063 30821
rect 22094 30812 22100 30824
rect 22152 30812 22158 30864
rect 21910 30784 21916 30796
rect 20456 30756 21916 30784
rect 14366 30676 14372 30728
rect 14424 30716 14430 30728
rect 14829 30719 14887 30725
rect 14829 30716 14841 30719
rect 14424 30688 14841 30716
rect 14424 30676 14430 30688
rect 14829 30685 14841 30688
rect 14875 30685 14887 30719
rect 14829 30679 14887 30685
rect 15013 30719 15071 30725
rect 15013 30685 15025 30719
rect 15059 30716 15071 30719
rect 15657 30719 15715 30725
rect 15657 30716 15669 30719
rect 15059 30688 15669 30716
rect 15059 30685 15071 30688
rect 15013 30679 15071 30685
rect 15657 30685 15669 30688
rect 15703 30685 15715 30719
rect 15657 30679 15715 30685
rect 17129 30719 17187 30725
rect 17129 30685 17141 30719
rect 17175 30716 17187 30719
rect 17218 30716 17224 30728
rect 17175 30688 17224 30716
rect 17175 30685 17187 30688
rect 17129 30679 17187 30685
rect 17218 30676 17224 30688
rect 17276 30676 17282 30728
rect 20456 30725 20484 30756
rect 21910 30744 21916 30756
rect 21968 30744 21974 30796
rect 27522 30784 27528 30796
rect 27483 30756 27528 30784
rect 27522 30744 27528 30756
rect 27580 30744 27586 30796
rect 27982 30784 27988 30796
rect 27943 30756 27988 30784
rect 27982 30744 27988 30756
rect 28040 30744 28046 30796
rect 28166 30784 28172 30796
rect 28127 30756 28172 30784
rect 28166 30744 28172 30756
rect 28224 30744 28230 30796
rect 20441 30719 20499 30725
rect 20441 30685 20453 30719
rect 20487 30685 20499 30719
rect 20441 30679 20499 30685
rect 20806 30676 20812 30728
rect 20864 30716 20870 30728
rect 20901 30719 20959 30725
rect 20901 30716 20913 30719
rect 20864 30688 20913 30716
rect 20864 30676 20870 30688
rect 20901 30685 20913 30688
rect 20947 30685 20959 30719
rect 20901 30679 20959 30685
rect 24854 30676 24860 30728
rect 24912 30716 24918 30728
rect 24949 30719 25007 30725
rect 24949 30716 24961 30719
rect 24912 30688 24961 30716
rect 24912 30676 24918 30688
rect 24949 30685 24961 30688
rect 24995 30685 25007 30719
rect 24949 30679 25007 30685
rect 25133 30719 25191 30725
rect 25133 30685 25145 30719
rect 25179 30716 25191 30719
rect 26142 30716 26148 30728
rect 25179 30688 26148 30716
rect 25179 30685 25191 30688
rect 25133 30679 25191 30685
rect 26142 30676 26148 30688
rect 26200 30676 26206 30728
rect 14642 30648 14648 30660
rect 14603 30620 14648 30648
rect 14642 30608 14648 30620
rect 14700 30608 14706 30660
rect 17310 30648 17316 30660
rect 17271 30620 17316 30648
rect 17310 30608 17316 30620
rect 17368 30608 17374 30660
rect 19242 30648 19248 30660
rect 19203 30620 19248 30648
rect 19242 30608 19248 30620
rect 19300 30608 19306 30660
rect 19429 30651 19487 30657
rect 19429 30617 19441 30651
rect 19475 30648 19487 30651
rect 19978 30648 19984 30660
rect 19475 30620 19984 30648
rect 19475 30617 19487 30620
rect 19429 30611 19487 30617
rect 19978 30608 19984 30620
rect 20036 30608 20042 30660
rect 20165 30651 20223 30657
rect 20165 30617 20177 30651
rect 20211 30648 20223 30651
rect 20254 30648 20260 30660
rect 20211 30620 20260 30648
rect 20211 30617 20223 30620
rect 20165 30611 20223 30617
rect 20254 30608 20260 30620
rect 20312 30608 20318 30660
rect 20349 30651 20407 30657
rect 20349 30617 20361 30651
rect 20395 30648 20407 30651
rect 20824 30648 20852 30676
rect 20395 30620 20852 30648
rect 21085 30651 21143 30657
rect 20395 30617 20407 30620
rect 20349 30611 20407 30617
rect 21085 30617 21097 30651
rect 21131 30648 21143 30651
rect 21634 30648 21640 30660
rect 21131 30620 21640 30648
rect 21131 30617 21143 30620
rect 21085 30611 21143 30617
rect 21634 30608 21640 30620
rect 21692 30648 21698 30660
rect 21821 30651 21879 30657
rect 21821 30648 21833 30651
rect 21692 30620 21833 30648
rect 21692 30608 21698 30620
rect 21821 30617 21833 30620
rect 21867 30617 21879 30651
rect 21821 30611 21879 30617
rect 15470 30580 15476 30592
rect 15431 30552 15476 30580
rect 15470 30540 15476 30552
rect 15528 30540 15534 30592
rect 16666 30540 16672 30592
rect 16724 30580 16730 30592
rect 16945 30583 17003 30589
rect 16945 30580 16957 30583
rect 16724 30552 16957 30580
rect 16724 30540 16730 30552
rect 16945 30549 16957 30552
rect 16991 30549 17003 30583
rect 16945 30543 17003 30549
rect 25041 30583 25099 30589
rect 25041 30549 25053 30583
rect 25087 30580 25099 30583
rect 25130 30580 25136 30592
rect 25087 30552 25136 30580
rect 25087 30549 25099 30552
rect 25041 30543 25099 30549
rect 25130 30540 25136 30552
rect 25188 30540 25194 30592
rect 1104 30490 28888 30512
rect 1104 30438 10214 30490
rect 10266 30438 10278 30490
rect 10330 30438 10342 30490
rect 10394 30438 10406 30490
rect 10458 30438 10470 30490
rect 10522 30438 19478 30490
rect 19530 30438 19542 30490
rect 19594 30438 19606 30490
rect 19658 30438 19670 30490
rect 19722 30438 19734 30490
rect 19786 30438 28888 30490
rect 1104 30416 28888 30438
rect 17310 30376 17316 30388
rect 17271 30348 17316 30376
rect 17310 30336 17316 30348
rect 17368 30336 17374 30388
rect 19978 30336 19984 30388
rect 20036 30376 20042 30388
rect 22462 30376 22468 30388
rect 20036 30348 21096 30376
rect 22423 30348 22468 30376
rect 20036 30336 20042 30348
rect 14912 30311 14970 30317
rect 14912 30277 14924 30311
rect 14958 30308 14970 30311
rect 15470 30308 15476 30320
rect 14958 30280 15476 30308
rect 14958 30277 14970 30280
rect 14912 30271 14970 30277
rect 15470 30268 15476 30280
rect 15528 30268 15534 30320
rect 17681 30311 17739 30317
rect 17681 30277 17693 30311
rect 17727 30308 17739 30311
rect 17770 30308 17776 30320
rect 17727 30280 17776 30308
rect 17727 30277 17739 30280
rect 17681 30271 17739 30277
rect 17770 30268 17776 30280
rect 17828 30268 17834 30320
rect 21068 30308 21096 30348
rect 22462 30336 22468 30348
rect 22520 30336 22526 30388
rect 23017 30311 23075 30317
rect 23017 30308 23029 30311
rect 21068 30280 23029 30308
rect 23017 30277 23029 30280
rect 23063 30277 23075 30311
rect 23017 30271 23075 30277
rect 1394 30240 1400 30252
rect 1355 30212 1400 30240
rect 1394 30200 1400 30212
rect 1452 30200 1458 30252
rect 16666 30240 16672 30252
rect 16627 30212 16672 30240
rect 16666 30200 16672 30212
rect 16724 30200 16730 30252
rect 19245 30243 19303 30249
rect 19245 30209 19257 30243
rect 19291 30240 19303 30243
rect 19334 30240 19340 30252
rect 19291 30212 19340 30240
rect 19291 30209 19303 30212
rect 19245 30203 19303 30209
rect 19334 30200 19340 30212
rect 19392 30200 19398 30252
rect 19705 30243 19763 30249
rect 19705 30209 19717 30243
rect 19751 30209 19763 30243
rect 19705 30203 19763 30209
rect 13998 30132 14004 30184
rect 14056 30172 14062 30184
rect 14645 30175 14703 30181
rect 14645 30172 14657 30175
rect 14056 30144 14657 30172
rect 14056 30132 14062 30144
rect 14645 30141 14657 30144
rect 14691 30141 14703 30175
rect 14645 30135 14703 30141
rect 17773 30175 17831 30181
rect 17773 30141 17785 30175
rect 17819 30141 17831 30175
rect 17773 30135 17831 30141
rect 17788 30104 17816 30135
rect 17862 30132 17868 30184
rect 17920 30172 17926 30184
rect 18966 30172 18972 30184
rect 17920 30144 17965 30172
rect 18927 30144 18972 30172
rect 17920 30132 17926 30144
rect 18966 30132 18972 30144
rect 19024 30132 19030 30184
rect 19720 30172 19748 30203
rect 19794 30200 19800 30252
rect 19852 30240 19858 30252
rect 19981 30243 20039 30249
rect 19852 30212 19897 30240
rect 19852 30200 19858 30212
rect 19981 30209 19993 30243
rect 20027 30240 20039 30243
rect 20162 30240 20168 30252
rect 20027 30212 20168 30240
rect 20027 30209 20039 30212
rect 19981 30203 20039 30209
rect 20162 30200 20168 30212
rect 20220 30200 20226 30252
rect 20254 30200 20260 30252
rect 20312 30240 20318 30252
rect 20671 30243 20729 30249
rect 20671 30240 20683 30243
rect 20312 30212 20683 30240
rect 20312 30200 20318 30212
rect 20671 30209 20683 30212
rect 20717 30209 20729 30243
rect 20806 30240 20812 30252
rect 20767 30212 20812 30240
rect 20671 30203 20729 30209
rect 20806 30200 20812 30212
rect 20864 30200 20870 30252
rect 20901 30243 20959 30249
rect 20901 30209 20913 30243
rect 20947 30209 20959 30243
rect 20901 30203 20959 30209
rect 21085 30243 21143 30249
rect 21085 30209 21097 30243
rect 21131 30240 21143 30243
rect 21818 30240 21824 30252
rect 21131 30212 21588 30240
rect 21779 30212 21824 30240
rect 21131 30209 21143 30212
rect 21085 30203 21143 30209
rect 20905 30172 20933 30203
rect 21358 30172 21364 30184
rect 19720 30144 20852 30172
rect 20905 30144 21364 30172
rect 20824 30116 20852 30144
rect 21358 30132 21364 30144
rect 21416 30132 21422 30184
rect 19058 30104 19064 30116
rect 17788 30076 19064 30104
rect 19058 30064 19064 30076
rect 19116 30064 19122 30116
rect 19153 30107 19211 30113
rect 19153 30073 19165 30107
rect 19199 30104 19211 30107
rect 20441 30107 20499 30113
rect 20441 30104 20453 30107
rect 19199 30076 20453 30104
rect 19199 30073 19211 30076
rect 19153 30067 19211 30073
rect 20441 30073 20453 30076
rect 20487 30073 20499 30107
rect 20441 30067 20499 30073
rect 20806 30064 20812 30116
rect 20864 30064 20870 30116
rect 1581 30039 1639 30045
rect 1581 30005 1593 30039
rect 1627 30036 1639 30039
rect 14550 30036 14556 30048
rect 1627 30008 14556 30036
rect 1627 30005 1639 30008
rect 1581 29999 1639 30005
rect 14550 29996 14556 30008
rect 14608 29996 14614 30048
rect 16025 30039 16083 30045
rect 16025 30005 16037 30039
rect 16071 30036 16083 30039
rect 16114 30036 16120 30048
rect 16071 30008 16120 30036
rect 16071 30005 16083 30008
rect 16025 29999 16083 30005
rect 16114 29996 16120 30008
rect 16172 29996 16178 30048
rect 16853 30039 16911 30045
rect 16853 30005 16865 30039
rect 16899 30036 16911 30039
rect 16942 30036 16948 30048
rect 16899 30008 16948 30036
rect 16899 30005 16911 30008
rect 16853 29999 16911 30005
rect 16942 29996 16948 30008
rect 17000 29996 17006 30048
rect 19245 30039 19303 30045
rect 19245 30005 19257 30039
rect 19291 30036 19303 30039
rect 19334 30036 19340 30048
rect 19291 30008 19340 30036
rect 19291 30005 19303 30008
rect 19245 29999 19303 30005
rect 19334 29996 19340 30008
rect 19392 29996 19398 30048
rect 19981 30039 20039 30045
rect 19981 30005 19993 30039
rect 20027 30036 20039 30039
rect 21560 30036 21588 30212
rect 21818 30200 21824 30212
rect 21876 30200 21882 30252
rect 22002 30240 22008 30252
rect 21963 30212 22008 30240
rect 22002 30200 22008 30212
rect 22060 30200 22066 30252
rect 25130 30249 25136 30252
rect 22097 30243 22155 30249
rect 22097 30209 22109 30243
rect 22143 30209 22155 30243
rect 22097 30203 22155 30209
rect 22189 30243 22247 30249
rect 22189 30209 22201 30243
rect 22235 30209 22247 30243
rect 25124 30240 25136 30249
rect 25091 30212 25136 30240
rect 22189 30203 22247 30209
rect 25124 30203 25136 30212
rect 21910 30132 21916 30184
rect 21968 30172 21974 30184
rect 22112 30172 22140 30203
rect 21968 30144 22140 30172
rect 21968 30132 21974 30144
rect 21726 30064 21732 30116
rect 21784 30104 21790 30116
rect 22204 30104 22232 30203
rect 25130 30200 25136 30203
rect 25188 30200 25194 30252
rect 26970 30200 26976 30252
rect 27028 30240 27034 30252
rect 27157 30243 27215 30249
rect 27157 30240 27169 30243
rect 27028 30212 27169 30240
rect 27028 30200 27034 30212
rect 27157 30209 27169 30212
rect 27203 30240 27215 30243
rect 27614 30240 27620 30252
rect 27203 30212 27620 30240
rect 27203 30209 27215 30212
rect 27157 30203 27215 30209
rect 27614 30200 27620 30212
rect 27672 30200 27678 30252
rect 27798 30200 27804 30252
rect 27856 30240 27862 30252
rect 27985 30243 28043 30249
rect 27985 30240 27997 30243
rect 27856 30212 27997 30240
rect 27856 30200 27862 30212
rect 27985 30209 27997 30212
rect 28031 30209 28043 30243
rect 27985 30203 28043 30209
rect 24857 30175 24915 30181
rect 24857 30172 24869 30175
rect 24044 30144 24869 30172
rect 24044 30116 24072 30144
rect 24857 30141 24869 30144
rect 24903 30141 24915 30175
rect 24857 30135 24915 30141
rect 21784 30076 22232 30104
rect 23201 30107 23259 30113
rect 21784 30064 21790 30076
rect 23201 30073 23213 30107
rect 23247 30104 23259 30107
rect 23474 30104 23480 30116
rect 23247 30076 23480 30104
rect 23247 30073 23259 30076
rect 23201 30067 23259 30073
rect 23474 30064 23480 30076
rect 23532 30104 23538 30116
rect 24026 30104 24032 30116
rect 23532 30076 24032 30104
rect 23532 30064 23538 30076
rect 24026 30064 24032 30076
rect 24084 30064 24090 30116
rect 20027 30008 21588 30036
rect 20027 30005 20039 30008
rect 19981 29999 20039 30005
rect 26142 29996 26148 30048
rect 26200 30036 26206 30048
rect 26237 30039 26295 30045
rect 26237 30036 26249 30039
rect 26200 30008 26249 30036
rect 26200 29996 26206 30008
rect 26237 30005 26249 30008
rect 26283 30005 26295 30039
rect 26237 29999 26295 30005
rect 26510 29996 26516 30048
rect 26568 30036 26574 30048
rect 27065 30039 27123 30045
rect 27065 30036 27077 30039
rect 26568 30008 27077 30036
rect 26568 29996 26574 30008
rect 27065 30005 27077 30008
rect 27111 30005 27123 30039
rect 27065 29999 27123 30005
rect 27893 30039 27951 30045
rect 27893 30005 27905 30039
rect 27939 30036 27951 30039
rect 28534 30036 28540 30048
rect 27939 30008 28540 30036
rect 27939 30005 27951 30008
rect 27893 29999 27951 30005
rect 28534 29996 28540 30008
rect 28592 29996 28598 30048
rect 1104 29946 28888 29968
rect 1104 29894 5582 29946
rect 5634 29894 5646 29946
rect 5698 29894 5710 29946
rect 5762 29894 5774 29946
rect 5826 29894 5838 29946
rect 5890 29894 14846 29946
rect 14898 29894 14910 29946
rect 14962 29894 14974 29946
rect 15026 29894 15038 29946
rect 15090 29894 15102 29946
rect 15154 29894 24110 29946
rect 24162 29894 24174 29946
rect 24226 29894 24238 29946
rect 24290 29894 24302 29946
rect 24354 29894 24366 29946
rect 24418 29894 28888 29946
rect 1104 29872 28888 29894
rect 14642 29792 14648 29844
rect 14700 29832 14706 29844
rect 14737 29835 14795 29841
rect 14737 29832 14749 29835
rect 14700 29804 14749 29832
rect 14700 29792 14706 29804
rect 14737 29801 14749 29804
rect 14783 29801 14795 29835
rect 14737 29795 14795 29801
rect 16117 29835 16175 29841
rect 16117 29801 16129 29835
rect 16163 29832 16175 29835
rect 16574 29832 16580 29844
rect 16163 29804 16580 29832
rect 16163 29801 16175 29804
rect 16117 29795 16175 29801
rect 16574 29792 16580 29804
rect 16632 29832 16638 29844
rect 17862 29832 17868 29844
rect 16632 29804 17868 29832
rect 16632 29792 16638 29804
rect 17862 29792 17868 29804
rect 17920 29792 17926 29844
rect 20162 29792 20168 29844
rect 20220 29832 20226 29844
rect 21637 29835 21695 29841
rect 21637 29832 21649 29835
rect 20220 29804 21649 29832
rect 20220 29792 20226 29804
rect 21637 29801 21649 29804
rect 21683 29801 21695 29835
rect 21637 29795 21695 29801
rect 22002 29792 22008 29844
rect 22060 29832 22066 29844
rect 22097 29835 22155 29841
rect 22097 29832 22109 29835
rect 22060 29804 22109 29832
rect 22060 29792 22066 29804
rect 22097 29801 22109 29804
rect 22143 29801 22155 29835
rect 22097 29795 22155 29801
rect 14458 29724 14464 29776
rect 14516 29764 14522 29776
rect 14516 29736 15976 29764
rect 14516 29724 14522 29736
rect 14550 29656 14556 29708
rect 14608 29696 14614 29708
rect 15304 29705 15332 29736
rect 15197 29699 15255 29705
rect 15197 29696 15209 29699
rect 14608 29668 15209 29696
rect 14608 29656 14614 29668
rect 15197 29665 15209 29668
rect 15243 29665 15255 29699
rect 15197 29659 15255 29665
rect 15289 29699 15347 29705
rect 15289 29665 15301 29699
rect 15335 29665 15347 29699
rect 15289 29659 15347 29665
rect 15948 29637 15976 29736
rect 20806 29724 20812 29776
rect 20864 29764 20870 29776
rect 21450 29764 21456 29776
rect 20864 29736 21456 29764
rect 20864 29724 20870 29736
rect 21450 29724 21456 29736
rect 21508 29724 21514 29776
rect 20990 29656 20996 29708
rect 21048 29696 21054 29708
rect 21818 29696 21824 29708
rect 21048 29668 21824 29696
rect 21048 29656 21054 29668
rect 21818 29656 21824 29668
rect 21876 29656 21882 29708
rect 23014 29656 23020 29708
rect 23072 29696 23078 29708
rect 23658 29696 23664 29708
rect 23072 29668 23244 29696
rect 23072 29656 23078 29668
rect 15933 29631 15991 29637
rect 15933 29597 15945 29631
rect 15979 29597 15991 29631
rect 15933 29591 15991 29597
rect 16853 29631 16911 29637
rect 16853 29597 16865 29631
rect 16899 29597 16911 29631
rect 16853 29591 16911 29597
rect 13998 29520 14004 29572
rect 14056 29560 14062 29572
rect 16868 29560 16896 29591
rect 16942 29588 16948 29640
rect 17000 29628 17006 29640
rect 17120 29631 17178 29637
rect 17120 29628 17132 29631
rect 17000 29600 17132 29628
rect 17000 29588 17006 29600
rect 17120 29597 17132 29600
rect 17166 29597 17178 29631
rect 19242 29628 19248 29640
rect 17120 29591 17178 29597
rect 17236 29600 19248 29628
rect 14056 29532 16896 29560
rect 14056 29520 14062 29532
rect 15105 29495 15163 29501
rect 15105 29461 15117 29495
rect 15151 29492 15163 29495
rect 16114 29492 16120 29504
rect 15151 29464 16120 29492
rect 15151 29461 15163 29464
rect 15105 29455 15163 29461
rect 16114 29452 16120 29464
rect 16172 29452 16178 29504
rect 16868 29492 16896 29532
rect 17236 29492 17264 29600
rect 19242 29588 19248 29600
rect 19300 29588 19306 29640
rect 19334 29588 19340 29640
rect 19392 29628 19398 29640
rect 19501 29631 19559 29637
rect 19501 29628 19513 29631
rect 19392 29600 19513 29628
rect 19392 29588 19398 29600
rect 19501 29597 19513 29600
rect 19547 29597 19559 29631
rect 19501 29591 19559 29597
rect 19794 29588 19800 29640
rect 19852 29628 19858 29640
rect 20438 29628 20444 29640
rect 19852 29600 20444 29628
rect 19852 29588 19858 29600
rect 20438 29588 20444 29600
rect 20496 29628 20502 29640
rect 21450 29628 21456 29640
rect 20496 29600 21456 29628
rect 20496 29588 20502 29600
rect 21450 29588 21456 29600
rect 21508 29588 21514 29640
rect 21545 29631 21603 29637
rect 21545 29597 21557 29631
rect 21591 29628 21603 29631
rect 21726 29628 21732 29640
rect 21591 29600 21732 29628
rect 21591 29597 21603 29600
rect 21545 29591 21603 29597
rect 21726 29588 21732 29600
rect 21784 29588 21790 29640
rect 22554 29628 22560 29640
rect 22515 29600 22560 29628
rect 22554 29588 22560 29600
rect 22612 29588 22618 29640
rect 22741 29631 22799 29637
rect 22741 29597 22753 29631
rect 22787 29628 22799 29631
rect 23106 29628 23112 29640
rect 22787 29600 23112 29628
rect 22787 29597 22799 29600
rect 22741 29591 22799 29597
rect 23106 29588 23112 29600
rect 23164 29588 23170 29640
rect 23216 29637 23244 29668
rect 23400 29668 23664 29696
rect 23400 29637 23428 29668
rect 23658 29656 23664 29668
rect 23716 29656 23722 29708
rect 26510 29696 26516 29708
rect 26471 29668 26516 29696
rect 26510 29656 26516 29668
rect 26568 29656 26574 29708
rect 28169 29699 28227 29705
rect 28169 29665 28181 29699
rect 28215 29696 28227 29699
rect 28718 29696 28724 29708
rect 28215 29668 28724 29696
rect 28215 29665 28227 29668
rect 28169 29659 28227 29665
rect 28718 29656 28724 29668
rect 28776 29656 28782 29708
rect 23201 29631 23259 29637
rect 23201 29597 23213 29631
rect 23247 29597 23259 29631
rect 23201 29591 23259 29597
rect 23385 29631 23443 29637
rect 23385 29597 23397 29631
rect 23431 29597 23443 29631
rect 23385 29591 23443 29597
rect 23477 29631 23535 29637
rect 23477 29597 23489 29631
rect 23523 29597 23535 29631
rect 23477 29591 23535 29597
rect 16868 29464 17264 29492
rect 17770 29452 17776 29504
rect 17828 29492 17834 29504
rect 18233 29495 18291 29501
rect 18233 29492 18245 29495
rect 17828 29464 18245 29492
rect 17828 29452 17834 29464
rect 18233 29461 18245 29464
rect 18279 29461 18291 29495
rect 18233 29455 18291 29461
rect 20162 29452 20168 29504
rect 20220 29492 20226 29504
rect 20625 29495 20683 29501
rect 20625 29492 20637 29495
rect 20220 29464 20637 29492
rect 20220 29452 20226 29464
rect 20625 29461 20637 29464
rect 20671 29461 20683 29495
rect 22572 29492 22600 29588
rect 22649 29563 22707 29569
rect 22649 29529 22661 29563
rect 22695 29560 22707 29563
rect 23492 29560 23520 29591
rect 23566 29588 23572 29640
rect 23624 29628 23630 29640
rect 23624 29600 23669 29628
rect 23624 29588 23630 29600
rect 24026 29588 24032 29640
rect 24084 29628 24090 29640
rect 25777 29631 25835 29637
rect 25777 29628 25789 29631
rect 24084 29600 25789 29628
rect 24084 29588 24090 29600
rect 25777 29597 25789 29600
rect 25823 29597 25835 29631
rect 25777 29591 25835 29597
rect 26329 29631 26387 29637
rect 26329 29597 26341 29631
rect 26375 29597 26387 29631
rect 26329 29591 26387 29597
rect 22695 29532 23520 29560
rect 23845 29563 23903 29569
rect 22695 29529 22707 29532
rect 22649 29523 22707 29529
rect 23845 29529 23857 29563
rect 23891 29560 23903 29563
rect 25510 29563 25568 29569
rect 25510 29560 25522 29563
rect 23891 29532 25522 29560
rect 23891 29529 23903 29532
rect 23845 29523 23903 29529
rect 25510 29529 25522 29532
rect 25556 29529 25568 29563
rect 25510 29523 25568 29529
rect 25682 29520 25688 29572
rect 25740 29560 25746 29572
rect 26142 29560 26148 29572
rect 25740 29532 26148 29560
rect 25740 29520 25746 29532
rect 26142 29520 26148 29532
rect 26200 29560 26206 29572
rect 26344 29560 26372 29591
rect 26200 29532 26372 29560
rect 26200 29520 26206 29532
rect 24397 29495 24455 29501
rect 24397 29492 24409 29495
rect 22572 29464 24409 29492
rect 20625 29455 20683 29461
rect 24397 29461 24409 29464
rect 24443 29461 24455 29495
rect 24397 29455 24455 29461
rect 1104 29402 28888 29424
rect 1104 29350 10214 29402
rect 10266 29350 10278 29402
rect 10330 29350 10342 29402
rect 10394 29350 10406 29402
rect 10458 29350 10470 29402
rect 10522 29350 19478 29402
rect 19530 29350 19542 29402
rect 19594 29350 19606 29402
rect 19658 29350 19670 29402
rect 19722 29350 19734 29402
rect 19786 29350 28888 29402
rect 1104 29328 28888 29350
rect 19058 29248 19064 29300
rect 19116 29288 19122 29300
rect 27157 29291 27215 29297
rect 27157 29288 27169 29291
rect 19116 29260 27169 29288
rect 19116 29248 19122 29260
rect 27157 29257 27169 29260
rect 27203 29257 27215 29291
rect 27157 29251 27215 29257
rect 27338 29152 27344 29164
rect 27299 29124 27344 29152
rect 27338 29112 27344 29124
rect 27396 29112 27402 29164
rect 13354 28976 13360 29028
rect 13412 29016 13418 29028
rect 16574 29016 16580 29028
rect 13412 28988 16580 29016
rect 13412 28976 13418 28988
rect 16574 28976 16580 28988
rect 16632 28976 16638 29028
rect 27982 28948 27988 28960
rect 27943 28920 27988 28948
rect 27982 28908 27988 28920
rect 28040 28908 28046 28960
rect 1104 28858 28888 28880
rect 1104 28806 5582 28858
rect 5634 28806 5646 28858
rect 5698 28806 5710 28858
rect 5762 28806 5774 28858
rect 5826 28806 5838 28858
rect 5890 28806 14846 28858
rect 14898 28806 14910 28858
rect 14962 28806 14974 28858
rect 15026 28806 15038 28858
rect 15090 28806 15102 28858
rect 15154 28806 24110 28858
rect 24162 28806 24174 28858
rect 24226 28806 24238 28858
rect 24290 28806 24302 28858
rect 24354 28806 24366 28858
rect 24418 28806 28888 28858
rect 1104 28784 28888 28806
rect 21818 28744 21824 28756
rect 21779 28716 21824 28744
rect 21818 28704 21824 28716
rect 21876 28704 21882 28756
rect 23569 28747 23627 28753
rect 23569 28713 23581 28747
rect 23615 28744 23627 28747
rect 23658 28744 23664 28756
rect 23615 28716 23664 28744
rect 23615 28713 23627 28716
rect 23569 28707 23627 28713
rect 23658 28704 23664 28716
rect 23716 28704 23722 28756
rect 17681 28679 17739 28685
rect 17681 28645 17693 28679
rect 17727 28676 17739 28679
rect 17862 28676 17868 28688
rect 17727 28648 17868 28676
rect 17727 28645 17739 28648
rect 17681 28639 17739 28645
rect 17862 28636 17868 28648
rect 17920 28636 17926 28688
rect 27522 28608 27528 28620
rect 27483 28580 27528 28608
rect 27522 28568 27528 28580
rect 27580 28568 27586 28620
rect 27982 28568 27988 28620
rect 28040 28608 28046 28620
rect 28169 28611 28227 28617
rect 28169 28608 28181 28611
rect 28040 28580 28181 28608
rect 28040 28568 28046 28580
rect 28169 28577 28181 28580
rect 28215 28577 28227 28611
rect 28169 28571 28227 28577
rect 21450 28500 21456 28552
rect 21508 28540 21514 28552
rect 21729 28543 21787 28549
rect 21729 28540 21741 28543
rect 21508 28512 21741 28540
rect 21508 28500 21514 28512
rect 21729 28509 21741 28512
rect 21775 28509 21787 28543
rect 21729 28503 21787 28509
rect 22094 28500 22100 28552
rect 22152 28540 22158 28552
rect 22465 28543 22523 28549
rect 22465 28540 22477 28543
rect 22152 28512 22477 28540
rect 22152 28500 22158 28512
rect 22465 28509 22477 28512
rect 22511 28509 22523 28543
rect 22465 28503 22523 28509
rect 22649 28543 22707 28549
rect 22649 28509 22661 28543
rect 22695 28540 22707 28543
rect 22738 28540 22744 28552
rect 22695 28512 22744 28540
rect 22695 28509 22707 28512
rect 22649 28503 22707 28509
rect 22738 28500 22744 28512
rect 22796 28500 22802 28552
rect 23109 28543 23167 28549
rect 23109 28509 23121 28543
rect 23155 28540 23167 28543
rect 23290 28540 23296 28552
rect 23155 28512 23296 28540
rect 23155 28509 23167 28512
rect 23109 28503 23167 28509
rect 23290 28500 23296 28512
rect 23348 28500 23354 28552
rect 23385 28543 23443 28549
rect 23385 28509 23397 28543
rect 23431 28509 23443 28543
rect 23385 28503 23443 28509
rect 14182 28472 14188 28484
rect 14143 28444 14188 28472
rect 14182 28432 14188 28444
rect 14240 28432 14246 28484
rect 14366 28472 14372 28484
rect 14327 28444 14372 28472
rect 14366 28432 14372 28444
rect 14424 28432 14430 28484
rect 17313 28475 17371 28481
rect 17313 28441 17325 28475
rect 17359 28472 17371 28475
rect 17586 28472 17592 28484
rect 17359 28444 17592 28472
rect 17359 28441 17371 28444
rect 17313 28435 17371 28441
rect 17586 28432 17592 28444
rect 17644 28432 17650 28484
rect 23400 28472 23428 28503
rect 22664 28444 23428 28472
rect 22664 28416 22692 28444
rect 27338 28432 27344 28484
rect 27396 28472 27402 28484
rect 27985 28475 28043 28481
rect 27985 28472 27997 28475
rect 27396 28444 27997 28472
rect 27396 28432 27402 28444
rect 27985 28441 27997 28444
rect 28031 28441 28043 28475
rect 27985 28435 28043 28441
rect 13814 28364 13820 28416
rect 13872 28404 13878 28416
rect 14553 28407 14611 28413
rect 14553 28404 14565 28407
rect 13872 28376 14565 28404
rect 13872 28364 13878 28376
rect 14553 28373 14565 28376
rect 14599 28373 14611 28407
rect 14553 28367 14611 28373
rect 17773 28407 17831 28413
rect 17773 28373 17785 28407
rect 17819 28404 17831 28407
rect 18506 28404 18512 28416
rect 17819 28376 18512 28404
rect 17819 28373 17831 28376
rect 17773 28367 17831 28373
rect 18506 28364 18512 28376
rect 18564 28364 18570 28416
rect 22554 28404 22560 28416
rect 22515 28376 22560 28404
rect 22554 28364 22560 28376
rect 22612 28364 22618 28416
rect 22646 28364 22652 28416
rect 22704 28364 22710 28416
rect 23201 28407 23259 28413
rect 23201 28373 23213 28407
rect 23247 28404 23259 28407
rect 23290 28404 23296 28416
rect 23247 28376 23296 28404
rect 23247 28373 23259 28376
rect 23201 28367 23259 28373
rect 23290 28364 23296 28376
rect 23348 28364 23354 28416
rect 1104 28314 28888 28336
rect 1104 28262 10214 28314
rect 10266 28262 10278 28314
rect 10330 28262 10342 28314
rect 10394 28262 10406 28314
rect 10458 28262 10470 28314
rect 10522 28262 19478 28314
rect 19530 28262 19542 28314
rect 19594 28262 19606 28314
rect 19658 28262 19670 28314
rect 19722 28262 19734 28314
rect 19786 28262 28888 28314
rect 1104 28240 28888 28262
rect 16117 28203 16175 28209
rect 16117 28169 16129 28203
rect 16163 28169 16175 28203
rect 20714 28200 20720 28212
rect 20675 28172 20720 28200
rect 16117 28163 16175 28169
rect 14642 28132 14648 28144
rect 12406 28104 14648 28132
rect 1394 28064 1400 28076
rect 1355 28036 1400 28064
rect 1394 28024 1400 28036
rect 1452 28024 1458 28076
rect 1581 27863 1639 27869
rect 1581 27829 1593 27863
rect 1627 27860 1639 27863
rect 12406 27860 12434 28104
rect 14642 28092 14648 28104
rect 14700 28092 14706 28144
rect 15746 28132 15752 28144
rect 15707 28104 15752 28132
rect 15746 28092 15752 28104
rect 15804 28092 15810 28144
rect 15949 28135 16007 28141
rect 15949 28132 15961 28135
rect 15948 28101 15961 28132
rect 15995 28101 16007 28135
rect 15948 28095 16007 28101
rect 13630 28073 13636 28076
rect 13624 28027 13636 28073
rect 13688 28064 13694 28076
rect 13688 28036 13724 28064
rect 13630 28024 13636 28027
rect 13688 28024 13694 28036
rect 13357 27999 13415 28005
rect 13357 27965 13369 27999
rect 13403 27965 13415 27999
rect 15948 27996 15976 28095
rect 16132 28064 16160 28163
rect 20714 28160 20720 28172
rect 20772 28160 20778 28212
rect 22094 28160 22100 28212
rect 22152 28200 22158 28212
rect 25501 28203 25559 28209
rect 25501 28200 25513 28203
rect 22152 28172 22197 28200
rect 22388 28172 25513 28200
rect 22152 28160 22158 28172
rect 21818 28132 21824 28144
rect 19444 28104 21824 28132
rect 16853 28067 16911 28073
rect 16853 28064 16865 28067
rect 16132 28036 16865 28064
rect 16853 28033 16865 28036
rect 16899 28033 16911 28067
rect 16853 28027 16911 28033
rect 18046 28024 18052 28076
rect 18104 28064 18110 28076
rect 18325 28067 18383 28073
rect 18325 28064 18337 28067
rect 18104 28036 18337 28064
rect 18104 28024 18110 28036
rect 18325 28033 18337 28036
rect 18371 28033 18383 28067
rect 18506 28064 18512 28076
rect 18467 28036 18512 28064
rect 18325 28027 18383 28033
rect 18506 28024 18512 28036
rect 18564 28024 18570 28076
rect 18598 28024 18604 28076
rect 18656 28064 18662 28076
rect 19444 28073 19472 28104
rect 21818 28092 21824 28104
rect 21876 28092 21882 28144
rect 22388 28076 22416 28172
rect 25501 28169 25513 28172
rect 25547 28169 25559 28203
rect 27338 28200 27344 28212
rect 27299 28172 27344 28200
rect 25501 28163 25559 28169
rect 27338 28160 27344 28172
rect 27396 28160 27402 28212
rect 22554 28092 22560 28144
rect 22612 28132 22618 28144
rect 23661 28135 23719 28141
rect 22612 28104 23336 28132
rect 22612 28092 22618 28104
rect 19429 28067 19487 28073
rect 18656 28036 18701 28064
rect 18656 28024 18662 28036
rect 19429 28033 19441 28067
rect 19475 28033 19487 28067
rect 19429 28027 19487 28033
rect 19705 28067 19763 28073
rect 19705 28033 19717 28067
rect 19751 28064 19763 28067
rect 20162 28064 20168 28076
rect 19751 28036 20168 28064
rect 19751 28033 19763 28036
rect 19705 28027 19763 28033
rect 20162 28024 20168 28036
rect 20220 28024 20226 28076
rect 20530 28064 20536 28076
rect 20491 28036 20536 28064
rect 20530 28024 20536 28036
rect 20588 28024 20594 28076
rect 20625 28067 20683 28073
rect 20625 28033 20637 28067
rect 20671 28064 20683 28067
rect 20806 28064 20812 28076
rect 20671 28036 20812 28064
rect 20671 28033 20683 28036
rect 20625 28027 20683 28033
rect 16758 27996 16764 28008
rect 15948 27968 16764 27996
rect 13357 27959 13415 27965
rect 1627 27832 12434 27860
rect 13372 27860 13400 27959
rect 16758 27956 16764 27968
rect 16816 27956 16822 28008
rect 17405 27999 17463 28005
rect 17405 27965 17417 27999
rect 17451 27996 17463 27999
rect 17770 27996 17776 28008
rect 17451 27968 17776 27996
rect 17451 27965 17463 27968
rect 17405 27959 17463 27965
rect 17770 27956 17776 27968
rect 17828 27956 17834 28008
rect 19613 27999 19671 28005
rect 19613 27965 19625 27999
rect 19659 27996 19671 27999
rect 20640 27996 20668 28027
rect 20806 28024 20812 28036
rect 20864 28024 20870 28076
rect 22370 28064 22376 28076
rect 22331 28036 22376 28064
rect 22370 28024 22376 28036
rect 22428 28024 22434 28076
rect 23014 28064 23020 28076
rect 22975 28036 23020 28064
rect 23014 28024 23020 28036
rect 23072 28024 23078 28076
rect 23198 28064 23204 28076
rect 23159 28036 23204 28064
rect 23198 28024 23204 28036
rect 23256 28024 23262 28076
rect 23308 28073 23336 28104
rect 23661 28101 23673 28135
rect 23707 28132 23719 28135
rect 24366 28135 24424 28141
rect 24366 28132 24378 28135
rect 23707 28104 24378 28132
rect 23707 28101 23719 28104
rect 23661 28095 23719 28101
rect 24366 28101 24378 28104
rect 24412 28101 24424 28135
rect 24366 28095 24424 28101
rect 23293 28067 23351 28073
rect 23293 28033 23305 28067
rect 23339 28033 23351 28067
rect 23293 28027 23351 28033
rect 23385 28067 23443 28073
rect 23385 28033 23397 28067
rect 23431 28064 23443 28067
rect 23566 28064 23572 28076
rect 23431 28036 23572 28064
rect 23431 28033 23443 28036
rect 23385 28027 23443 28033
rect 23566 28024 23572 28036
rect 23624 28024 23630 28076
rect 27246 28064 27252 28076
rect 27207 28036 27252 28064
rect 27246 28024 27252 28036
rect 27304 28024 27310 28076
rect 19659 27968 20668 27996
rect 19659 27965 19671 27968
rect 19613 27959 19671 27965
rect 21818 27956 21824 28008
rect 21876 27996 21882 28008
rect 22097 27999 22155 28005
rect 22097 27996 22109 27999
rect 21876 27968 22109 27996
rect 21876 27956 21882 27968
rect 22097 27965 22109 27968
rect 22143 27965 22155 27999
rect 22097 27959 22155 27965
rect 24026 27956 24032 28008
rect 24084 27996 24090 28008
rect 24121 27999 24179 28005
rect 24121 27996 24133 27999
rect 24084 27968 24133 27996
rect 24084 27956 24090 27968
rect 24121 27965 24133 27968
rect 24167 27965 24179 27999
rect 24121 27959 24179 27965
rect 17678 27928 17684 27940
rect 17639 27900 17684 27928
rect 17678 27888 17684 27900
rect 17736 27888 17742 27940
rect 13998 27860 14004 27872
rect 13372 27832 14004 27860
rect 1627 27829 1639 27832
rect 1581 27823 1639 27829
rect 13998 27820 14004 27832
rect 14056 27820 14062 27872
rect 14734 27860 14740 27872
rect 14695 27832 14740 27860
rect 14734 27820 14740 27832
rect 14792 27820 14798 27872
rect 15930 27860 15936 27872
rect 15891 27832 15936 27860
rect 15930 27820 15936 27832
rect 15988 27820 15994 27872
rect 16666 27860 16672 27872
rect 16627 27832 16672 27860
rect 16666 27820 16672 27832
rect 16724 27820 16730 27872
rect 17865 27863 17923 27869
rect 17865 27829 17877 27863
rect 17911 27860 17923 27863
rect 18046 27860 18052 27872
rect 17911 27832 18052 27860
rect 17911 27829 17923 27832
rect 17865 27823 17923 27829
rect 18046 27820 18052 27832
rect 18104 27820 18110 27872
rect 18322 27860 18328 27872
rect 18283 27832 18328 27860
rect 18322 27820 18328 27832
rect 18380 27820 18386 27872
rect 18782 27860 18788 27872
rect 18743 27832 18788 27860
rect 18782 27820 18788 27832
rect 18840 27820 18846 27872
rect 19242 27860 19248 27872
rect 19203 27832 19248 27860
rect 19242 27820 19248 27832
rect 19300 27820 19306 27872
rect 22281 27863 22339 27869
rect 22281 27829 22293 27863
rect 22327 27860 22339 27863
rect 22554 27860 22560 27872
rect 22327 27832 22560 27860
rect 22327 27829 22339 27832
rect 22281 27823 22339 27829
rect 22554 27820 22560 27832
rect 22612 27820 22618 27872
rect 28077 27863 28135 27869
rect 28077 27829 28089 27863
rect 28123 27860 28135 27863
rect 28166 27860 28172 27872
rect 28123 27832 28172 27860
rect 28123 27829 28135 27832
rect 28077 27823 28135 27829
rect 28166 27820 28172 27832
rect 28224 27820 28230 27872
rect 1104 27770 28888 27792
rect 1104 27718 5582 27770
rect 5634 27718 5646 27770
rect 5698 27718 5710 27770
rect 5762 27718 5774 27770
rect 5826 27718 5838 27770
rect 5890 27718 14846 27770
rect 14898 27718 14910 27770
rect 14962 27718 14974 27770
rect 15026 27718 15038 27770
rect 15090 27718 15102 27770
rect 15154 27718 24110 27770
rect 24162 27718 24174 27770
rect 24226 27718 24238 27770
rect 24290 27718 24302 27770
rect 24354 27718 24366 27770
rect 24418 27718 28888 27770
rect 1104 27696 28888 27718
rect 13541 27659 13599 27665
rect 13541 27625 13553 27659
rect 13587 27656 13599 27659
rect 13630 27656 13636 27668
rect 13587 27628 13636 27656
rect 13587 27625 13599 27628
rect 13541 27619 13599 27625
rect 13630 27616 13636 27628
rect 13688 27616 13694 27668
rect 14182 27656 14188 27668
rect 14143 27628 14188 27656
rect 14182 27616 14188 27628
rect 14240 27616 14246 27668
rect 23017 27659 23075 27665
rect 23017 27625 23029 27659
rect 23063 27656 23075 27659
rect 23198 27656 23204 27668
rect 23063 27628 23204 27656
rect 23063 27625 23075 27628
rect 23017 27619 23075 27625
rect 23198 27616 23204 27628
rect 23256 27616 23262 27668
rect 13906 27548 13912 27600
rect 13964 27588 13970 27600
rect 14458 27588 14464 27600
rect 13964 27560 14464 27588
rect 13964 27548 13970 27560
rect 14458 27548 14464 27560
rect 14516 27588 14522 27600
rect 17037 27591 17095 27597
rect 14516 27560 14780 27588
rect 14516 27548 14522 27560
rect 14642 27520 14648 27532
rect 14603 27492 14648 27520
rect 14642 27480 14648 27492
rect 14700 27480 14706 27532
rect 14752 27529 14780 27560
rect 17037 27557 17049 27591
rect 17083 27588 17095 27591
rect 17310 27588 17316 27600
rect 17083 27560 17316 27588
rect 17083 27557 17095 27560
rect 17037 27551 17095 27557
rect 17310 27548 17316 27560
rect 17368 27588 17374 27600
rect 17368 27560 17540 27588
rect 17368 27548 17374 27560
rect 17512 27529 17540 27560
rect 20070 27548 20076 27600
rect 20128 27588 20134 27600
rect 21358 27588 21364 27600
rect 20128 27560 21364 27588
rect 20128 27548 20134 27560
rect 21358 27548 21364 27560
rect 21416 27548 21422 27600
rect 21634 27588 21640 27600
rect 21595 27560 21640 27588
rect 21634 27548 21640 27560
rect 21692 27548 21698 27600
rect 22373 27591 22431 27597
rect 22373 27557 22385 27591
rect 22419 27588 22431 27591
rect 23106 27588 23112 27600
rect 22419 27560 23112 27588
rect 22419 27557 22431 27560
rect 22373 27551 22431 27557
rect 23106 27548 23112 27560
rect 23164 27548 23170 27600
rect 14737 27523 14795 27529
rect 14737 27489 14749 27523
rect 14783 27489 14795 27523
rect 14737 27483 14795 27489
rect 17497 27523 17555 27529
rect 17497 27489 17509 27523
rect 17543 27489 17555 27523
rect 17497 27483 17555 27489
rect 17773 27523 17831 27529
rect 17773 27489 17785 27523
rect 17819 27520 17831 27523
rect 17862 27520 17868 27532
rect 17819 27492 17868 27520
rect 17819 27489 17831 27492
rect 17773 27483 17831 27489
rect 17862 27480 17868 27492
rect 17920 27480 17926 27532
rect 19705 27523 19763 27529
rect 19705 27489 19717 27523
rect 19751 27520 19763 27523
rect 20257 27523 20315 27529
rect 20257 27520 20269 27523
rect 19751 27492 20269 27520
rect 19751 27489 19763 27492
rect 19705 27483 19763 27489
rect 20257 27489 20269 27492
rect 20303 27520 20315 27523
rect 20530 27520 20536 27532
rect 20303 27492 20536 27520
rect 20303 27489 20315 27492
rect 20257 27483 20315 27489
rect 20530 27480 20536 27492
rect 20588 27520 20594 27532
rect 20588 27492 20668 27520
rect 20588 27480 20594 27492
rect 13357 27455 13415 27461
rect 13357 27421 13369 27455
rect 13403 27452 13415 27455
rect 13814 27452 13820 27464
rect 13403 27424 13820 27452
rect 13403 27421 13415 27424
rect 13357 27415 13415 27421
rect 13814 27412 13820 27424
rect 13872 27412 13878 27464
rect 13998 27412 14004 27464
rect 14056 27452 14062 27464
rect 15102 27452 15108 27464
rect 14056 27424 15108 27452
rect 14056 27412 14062 27424
rect 15102 27412 15108 27424
rect 15160 27452 15166 27464
rect 15657 27455 15715 27461
rect 15657 27452 15669 27455
rect 15160 27424 15669 27452
rect 15160 27412 15166 27424
rect 15657 27421 15669 27424
rect 15703 27421 15715 27455
rect 15657 27415 15715 27421
rect 15924 27455 15982 27461
rect 15924 27421 15936 27455
rect 15970 27452 15982 27455
rect 16666 27452 16672 27464
rect 15970 27424 16672 27452
rect 15970 27421 15982 27424
rect 15924 27415 15982 27421
rect 16666 27412 16672 27424
rect 16724 27412 16730 27464
rect 19797 27455 19855 27461
rect 19797 27421 19809 27455
rect 19843 27452 19855 27455
rect 20162 27452 20168 27464
rect 19843 27424 20168 27452
rect 19843 27421 19855 27424
rect 19797 27415 19855 27421
rect 20162 27412 20168 27424
rect 20220 27412 20226 27464
rect 20438 27452 20444 27464
rect 20399 27424 20444 27452
rect 20438 27412 20444 27424
rect 20496 27412 20502 27464
rect 20640 27452 20668 27492
rect 20714 27480 20720 27532
rect 20772 27520 20778 27532
rect 20809 27523 20867 27529
rect 20809 27520 20821 27523
rect 20772 27492 20821 27520
rect 20772 27480 20778 27492
rect 20809 27489 20821 27492
rect 20855 27489 20867 27523
rect 27522 27520 27528 27532
rect 27483 27492 27528 27520
rect 20809 27483 20867 27489
rect 27522 27480 27528 27492
rect 27580 27480 27586 27532
rect 28166 27520 28172 27532
rect 28127 27492 28172 27520
rect 28166 27480 28172 27492
rect 28224 27480 28230 27532
rect 22189 27455 22247 27461
rect 22189 27452 22201 27455
rect 20640 27424 22201 27452
rect 22189 27421 22201 27424
rect 22235 27421 22247 27455
rect 22189 27415 22247 27421
rect 22370 27412 22376 27464
rect 22428 27452 22434 27464
rect 22646 27452 22652 27464
rect 22428 27424 22652 27452
rect 22428 27412 22434 27424
rect 22646 27412 22652 27424
rect 22704 27452 22710 27464
rect 23201 27455 23259 27461
rect 23201 27452 23213 27455
rect 22704 27424 23213 27452
rect 22704 27412 22710 27424
rect 23201 27421 23213 27424
rect 23247 27421 23259 27455
rect 23201 27415 23259 27421
rect 23382 27412 23388 27464
rect 23440 27452 23446 27464
rect 23477 27455 23535 27461
rect 23477 27452 23489 27455
rect 23440 27424 23489 27452
rect 23440 27412 23446 27424
rect 23477 27421 23489 27424
rect 23523 27452 23535 27455
rect 23842 27452 23848 27464
rect 23523 27424 23848 27452
rect 23523 27421 23535 27424
rect 23477 27415 23535 27421
rect 23842 27412 23848 27424
rect 23900 27412 23906 27464
rect 14366 27344 14372 27396
rect 14424 27384 14430 27396
rect 20180 27384 20208 27412
rect 21269 27387 21327 27393
rect 21269 27384 21281 27387
rect 14424 27356 14872 27384
rect 20180 27356 21281 27384
rect 14424 27344 14430 27356
rect 14090 27276 14096 27328
rect 14148 27316 14154 27328
rect 14553 27319 14611 27325
rect 14553 27316 14565 27319
rect 14148 27288 14565 27316
rect 14148 27276 14154 27288
rect 14553 27285 14565 27288
rect 14599 27316 14611 27319
rect 14734 27316 14740 27328
rect 14599 27288 14740 27316
rect 14599 27285 14611 27288
rect 14553 27279 14611 27285
rect 14734 27276 14740 27288
rect 14792 27276 14798 27328
rect 14844 27316 14872 27356
rect 21269 27353 21281 27356
rect 21315 27353 21327 27387
rect 21269 27347 21327 27353
rect 21358 27344 21364 27396
rect 21416 27384 21422 27396
rect 21453 27387 21511 27393
rect 21453 27384 21465 27387
rect 21416 27356 21465 27384
rect 21416 27344 21422 27356
rect 21453 27353 21465 27356
rect 21499 27384 21511 27387
rect 21634 27384 21640 27396
rect 21499 27356 21640 27384
rect 21499 27353 21511 27356
rect 21453 27347 21511 27353
rect 21634 27344 21640 27356
rect 21692 27344 21698 27396
rect 27706 27344 27712 27396
rect 27764 27384 27770 27396
rect 27985 27387 28043 27393
rect 27985 27384 27997 27387
rect 27764 27356 27997 27384
rect 27764 27344 27770 27356
rect 27985 27353 27997 27356
rect 28031 27353 28043 27387
rect 27985 27347 28043 27353
rect 20346 27316 20352 27328
rect 14844 27288 20352 27316
rect 20346 27276 20352 27288
rect 20404 27276 20410 27328
rect 20717 27319 20775 27325
rect 20717 27285 20729 27319
rect 20763 27316 20775 27319
rect 21542 27316 21548 27328
rect 20763 27288 21548 27316
rect 20763 27285 20775 27288
rect 20717 27279 20775 27285
rect 21542 27276 21548 27288
rect 21600 27276 21606 27328
rect 23290 27276 23296 27328
rect 23348 27316 23354 27328
rect 23385 27319 23443 27325
rect 23385 27316 23397 27319
rect 23348 27288 23397 27316
rect 23348 27276 23354 27288
rect 23385 27285 23397 27288
rect 23431 27285 23443 27319
rect 23385 27279 23443 27285
rect 1104 27226 28888 27248
rect 1104 27174 10214 27226
rect 10266 27174 10278 27226
rect 10330 27174 10342 27226
rect 10394 27174 10406 27226
rect 10458 27174 10470 27226
rect 10522 27174 19478 27226
rect 19530 27174 19542 27226
rect 19594 27174 19606 27226
rect 19658 27174 19670 27226
rect 19722 27174 19734 27226
rect 19786 27174 28888 27226
rect 1104 27152 28888 27174
rect 15749 27115 15807 27121
rect 15749 27081 15761 27115
rect 15795 27112 15807 27115
rect 15930 27112 15936 27124
rect 15795 27084 15936 27112
rect 15795 27081 15807 27084
rect 15749 27075 15807 27081
rect 15930 27072 15936 27084
rect 15988 27072 15994 27124
rect 16758 27112 16764 27124
rect 16719 27084 16764 27112
rect 16758 27072 16764 27084
rect 16816 27072 16822 27124
rect 18690 27072 18696 27124
rect 18748 27112 18754 27124
rect 18748 27084 19380 27112
rect 18748 27072 18754 27084
rect 15102 27004 15108 27056
rect 15160 27044 15166 27056
rect 15160 27016 18920 27044
rect 15160 27004 15166 27016
rect 15930 26976 15936 26988
rect 15891 26948 15936 26976
rect 15930 26936 15936 26948
rect 15988 26936 15994 26988
rect 16117 26979 16175 26985
rect 16117 26945 16129 26979
rect 16163 26976 16175 26979
rect 16669 26979 16727 26985
rect 16669 26976 16681 26979
rect 16163 26948 16681 26976
rect 16163 26945 16175 26948
rect 16117 26939 16175 26945
rect 16669 26945 16681 26948
rect 16715 26945 16727 26979
rect 16669 26939 16727 26945
rect 16853 26979 16911 26985
rect 16853 26945 16865 26979
rect 16899 26945 16911 26979
rect 17310 26976 17316 26988
rect 17271 26948 17316 26976
rect 16853 26939 16911 26945
rect 15654 26868 15660 26920
rect 15712 26908 15718 26920
rect 16132 26908 16160 26939
rect 15712 26880 16160 26908
rect 16868 26908 16896 26939
rect 17310 26936 17316 26948
rect 17368 26936 17374 26988
rect 17862 26976 17868 26988
rect 17420 26948 17868 26976
rect 17420 26908 17448 26948
rect 17862 26936 17868 26948
rect 17920 26936 17926 26988
rect 18233 26979 18291 26985
rect 18233 26945 18245 26979
rect 18279 26976 18291 26979
rect 18322 26976 18328 26988
rect 18279 26948 18328 26976
rect 18279 26945 18291 26948
rect 18233 26939 18291 26945
rect 18322 26936 18328 26948
rect 18380 26936 18386 26988
rect 18417 26979 18475 26985
rect 18417 26945 18429 26979
rect 18463 26976 18475 26979
rect 18598 26976 18604 26988
rect 18463 26948 18604 26976
rect 18463 26945 18475 26948
rect 18417 26939 18475 26945
rect 16868 26880 17448 26908
rect 17773 26911 17831 26917
rect 15712 26868 15718 26880
rect 15930 26800 15936 26852
rect 15988 26840 15994 26852
rect 16868 26840 16896 26880
rect 17773 26877 17785 26911
rect 17819 26908 17831 26911
rect 18432 26908 18460 26939
rect 18598 26936 18604 26948
rect 18656 26936 18662 26988
rect 18892 26985 18920 27016
rect 19150 26985 19156 26988
rect 18877 26979 18935 26985
rect 18877 26945 18889 26979
rect 18923 26945 18935 26979
rect 18877 26939 18935 26945
rect 19144 26939 19156 26985
rect 19208 26976 19214 26988
rect 19352 26976 19380 27084
rect 20162 27072 20168 27124
rect 20220 27112 20226 27124
rect 20257 27115 20315 27121
rect 20257 27112 20269 27115
rect 20220 27084 20269 27112
rect 20220 27072 20226 27084
rect 20257 27081 20269 27084
rect 20303 27112 20315 27115
rect 27706 27112 27712 27124
rect 20303 27084 20852 27112
rect 20303 27081 20315 27084
rect 20257 27075 20315 27081
rect 20824 27053 20852 27084
rect 20916 27084 25912 27112
rect 27667 27084 27712 27112
rect 20809 27047 20867 27053
rect 20809 27013 20821 27047
rect 20855 27013 20867 27047
rect 20809 27007 20867 27013
rect 20916 26976 20944 27084
rect 20993 27047 21051 27053
rect 20993 27013 21005 27047
rect 21039 27044 21051 27047
rect 21450 27044 21456 27056
rect 21039 27016 21456 27044
rect 21039 27013 21051 27016
rect 20993 27007 21051 27013
rect 21450 27004 21456 27016
rect 21508 27004 21514 27056
rect 22830 27044 22836 27056
rect 22112 27016 22836 27044
rect 19208 26948 19244 26976
rect 19352 26948 20944 26976
rect 19150 26936 19156 26939
rect 19208 26936 19214 26948
rect 17819 26880 18460 26908
rect 21468 26908 21496 27004
rect 22112 26985 22140 27016
rect 22830 27004 22836 27016
rect 22888 27004 22894 27056
rect 25884 27044 25912 27084
rect 27706 27072 27712 27084
rect 27764 27072 27770 27124
rect 25884 27016 27660 27044
rect 22097 26979 22155 26985
rect 22097 26945 22109 26979
rect 22143 26945 22155 26979
rect 22097 26939 22155 26945
rect 22186 26936 22192 26988
rect 22244 26976 22250 26988
rect 22741 26979 22799 26985
rect 22741 26976 22753 26979
rect 22244 26948 22753 26976
rect 22244 26936 22250 26948
rect 22741 26945 22753 26948
rect 22787 26945 22799 26979
rect 22922 26976 22928 26988
rect 22883 26948 22928 26976
rect 22741 26939 22799 26945
rect 22922 26936 22928 26948
rect 22980 26936 22986 26988
rect 27632 26985 27660 27016
rect 27617 26979 27675 26985
rect 27617 26945 27629 26979
rect 27663 26976 27675 26979
rect 27890 26976 27896 26988
rect 27663 26948 27896 26976
rect 27663 26945 27675 26948
rect 27617 26939 27675 26945
rect 27890 26936 27896 26948
rect 27948 26936 27954 26988
rect 21821 26911 21879 26917
rect 21821 26908 21833 26911
rect 21468 26880 21833 26908
rect 17819 26877 17831 26880
rect 17773 26871 17831 26877
rect 21821 26877 21833 26880
rect 21867 26877 21879 26911
rect 21821 26871 21879 26877
rect 22005 26911 22063 26917
rect 22005 26877 22017 26911
rect 22051 26908 22063 26911
rect 22051 26880 22784 26908
rect 22051 26877 22063 26880
rect 22005 26871 22063 26877
rect 22756 26852 22784 26880
rect 17586 26840 17592 26852
rect 15988 26812 16896 26840
rect 17547 26812 17592 26840
rect 15988 26800 15994 26812
rect 17586 26800 17592 26812
rect 17644 26800 17650 26852
rect 22738 26800 22744 26852
rect 22796 26800 22802 26852
rect 18138 26732 18144 26784
rect 18196 26772 18202 26784
rect 18233 26775 18291 26781
rect 18233 26772 18245 26775
rect 18196 26744 18245 26772
rect 18196 26732 18202 26744
rect 18233 26741 18245 26744
rect 18279 26741 18291 26775
rect 21910 26772 21916 26784
rect 21871 26744 21916 26772
rect 18233 26735 18291 26741
rect 21910 26732 21916 26744
rect 21968 26732 21974 26784
rect 22925 26775 22983 26781
rect 22925 26741 22937 26775
rect 22971 26772 22983 26775
rect 23382 26772 23388 26784
rect 22971 26744 23388 26772
rect 22971 26741 22983 26744
rect 22925 26735 22983 26741
rect 23382 26732 23388 26744
rect 23440 26732 23446 26784
rect 1104 26682 28888 26704
rect 1104 26630 5582 26682
rect 5634 26630 5646 26682
rect 5698 26630 5710 26682
rect 5762 26630 5774 26682
rect 5826 26630 5838 26682
rect 5890 26630 14846 26682
rect 14898 26630 14910 26682
rect 14962 26630 14974 26682
rect 15026 26630 15038 26682
rect 15090 26630 15102 26682
rect 15154 26630 24110 26682
rect 24162 26630 24174 26682
rect 24226 26630 24238 26682
rect 24290 26630 24302 26682
rect 24354 26630 24366 26682
rect 24418 26630 28888 26682
rect 1104 26608 28888 26630
rect 17957 26571 18015 26577
rect 17957 26537 17969 26571
rect 18003 26568 18015 26571
rect 18322 26568 18328 26580
rect 18003 26540 18328 26568
rect 18003 26537 18015 26540
rect 17957 26531 18015 26537
rect 18322 26528 18328 26540
rect 18380 26528 18386 26580
rect 21542 26528 21548 26580
rect 21600 26568 21606 26580
rect 23198 26568 23204 26580
rect 21600 26540 23204 26568
rect 21600 26528 21606 26540
rect 23198 26528 23204 26540
rect 23256 26568 23262 26580
rect 23842 26568 23848 26580
rect 23256 26540 23848 26568
rect 23256 26528 23262 26540
rect 23842 26528 23848 26540
rect 23900 26528 23906 26580
rect 17770 26500 17776 26512
rect 17731 26472 17776 26500
rect 17770 26460 17776 26472
rect 17828 26460 17834 26512
rect 19058 26460 19064 26512
rect 19116 26500 19122 26512
rect 19245 26503 19303 26509
rect 19245 26500 19257 26503
rect 19116 26472 19257 26500
rect 19116 26460 19122 26472
rect 19245 26469 19257 26472
rect 19291 26469 19303 26503
rect 19245 26463 19303 26469
rect 21821 26503 21879 26509
rect 21821 26469 21833 26503
rect 21867 26500 21879 26503
rect 23750 26500 23756 26512
rect 21867 26472 23756 26500
rect 21867 26469 21879 26472
rect 21821 26463 21879 26469
rect 23750 26460 23756 26472
rect 23808 26460 23814 26512
rect 16482 26432 16488 26444
rect 15580 26404 16488 26432
rect 15580 26376 15608 26404
rect 16482 26392 16488 26404
rect 16540 26432 16546 26444
rect 17497 26435 17555 26441
rect 17497 26432 17509 26435
rect 16540 26404 17509 26432
rect 16540 26392 16546 26404
rect 17497 26401 17509 26404
rect 17543 26432 17555 26435
rect 17678 26432 17684 26444
rect 17543 26404 17684 26432
rect 17543 26401 17555 26404
rect 17497 26395 17555 26401
rect 17678 26392 17684 26404
rect 17736 26392 17742 26444
rect 21542 26432 21548 26444
rect 17788 26404 19472 26432
rect 21503 26404 21548 26432
rect 14734 26364 14740 26376
rect 14695 26336 14740 26364
rect 14734 26324 14740 26336
rect 14792 26324 14798 26376
rect 15562 26364 15568 26376
rect 15475 26336 15568 26364
rect 15562 26324 15568 26336
rect 15620 26324 15626 26376
rect 15654 26324 15660 26376
rect 15712 26364 15718 26376
rect 15841 26367 15899 26373
rect 15841 26364 15853 26367
rect 15712 26336 15853 26364
rect 15712 26324 15718 26336
rect 15841 26333 15853 26336
rect 15887 26333 15899 26367
rect 15841 26327 15899 26333
rect 16574 26324 16580 26376
rect 16632 26364 16638 26376
rect 17788 26364 17816 26404
rect 19242 26364 19248 26376
rect 16632 26336 17816 26364
rect 19203 26336 19248 26364
rect 16632 26324 16638 26336
rect 19242 26324 19248 26336
rect 19300 26324 19306 26376
rect 19444 26373 19472 26404
rect 21542 26392 21548 26404
rect 21600 26392 21606 26444
rect 21910 26392 21916 26444
rect 21968 26432 21974 26444
rect 21968 26404 22508 26432
rect 21968 26392 21974 26404
rect 19429 26367 19487 26373
rect 19429 26333 19441 26367
rect 19475 26333 19487 26367
rect 19429 26327 19487 26333
rect 19521 26367 19579 26373
rect 19521 26333 19533 26367
rect 19567 26333 19579 26367
rect 19521 26327 19579 26333
rect 15749 26299 15807 26305
rect 15749 26265 15761 26299
rect 15795 26296 15807 26299
rect 15930 26296 15936 26308
rect 15795 26268 15936 26296
rect 15795 26265 15807 26268
rect 15749 26259 15807 26265
rect 15930 26256 15936 26268
rect 15988 26256 15994 26308
rect 18506 26256 18512 26308
rect 18564 26296 18570 26308
rect 19536 26296 19564 26327
rect 19886 26324 19892 26376
rect 19944 26364 19950 26376
rect 19981 26367 20039 26373
rect 19981 26364 19993 26367
rect 19944 26336 19993 26364
rect 19944 26324 19950 26336
rect 19981 26333 19993 26336
rect 20027 26333 20039 26367
rect 19981 26327 20039 26333
rect 20346 26324 20352 26376
rect 20404 26364 20410 26376
rect 21358 26364 21364 26376
rect 20404 26336 21364 26364
rect 20404 26324 20410 26336
rect 21358 26324 21364 26336
rect 21416 26324 21422 26376
rect 22480 26373 22508 26404
rect 21453 26367 21511 26373
rect 21453 26333 21465 26367
rect 21499 26333 21511 26367
rect 21453 26327 21511 26333
rect 21637 26367 21695 26373
rect 21637 26333 21649 26367
rect 21683 26364 21695 26367
rect 22281 26367 22339 26373
rect 22281 26364 22293 26367
rect 21683 26336 22293 26364
rect 21683 26333 21695 26336
rect 21637 26327 21695 26333
rect 22281 26333 22293 26336
rect 22327 26333 22339 26367
rect 22281 26327 22339 26333
rect 22465 26367 22523 26373
rect 22465 26333 22477 26367
rect 22511 26333 22523 26367
rect 22738 26364 22744 26376
rect 22699 26336 22744 26364
rect 22465 26327 22523 26333
rect 18564 26268 19564 26296
rect 20073 26299 20131 26305
rect 18564 26256 18570 26268
rect 20073 26265 20085 26299
rect 20119 26296 20131 26299
rect 20438 26296 20444 26308
rect 20119 26268 20444 26296
rect 20119 26265 20131 26268
rect 20073 26259 20131 26265
rect 20438 26256 20444 26268
rect 20496 26256 20502 26308
rect 21468 26296 21496 26327
rect 22738 26324 22744 26336
rect 22796 26324 22802 26376
rect 23198 26364 23204 26376
rect 23159 26336 23204 26364
rect 23198 26324 23204 26336
rect 23256 26324 23262 26376
rect 23290 26324 23296 26376
rect 23348 26364 23354 26376
rect 23474 26364 23480 26376
rect 23348 26336 23393 26364
rect 23435 26336 23480 26364
rect 23348 26324 23354 26336
rect 23474 26324 23480 26336
rect 23532 26324 23538 26376
rect 24026 26324 24032 26376
rect 24084 26364 24090 26376
rect 24397 26367 24455 26373
rect 24397 26364 24409 26367
rect 24084 26336 24409 26364
rect 24084 26324 24090 26336
rect 24397 26333 24409 26336
rect 24443 26333 24455 26367
rect 24397 26327 24455 26333
rect 26418 26324 26424 26376
rect 26476 26364 26482 26376
rect 27249 26367 27307 26373
rect 27249 26364 27261 26367
rect 26476 26336 27261 26364
rect 26476 26324 26482 26336
rect 27249 26333 27261 26336
rect 27295 26333 27307 26367
rect 27249 26327 27307 26333
rect 28077 26367 28135 26373
rect 28077 26333 28089 26367
rect 28123 26364 28135 26367
rect 28166 26364 28172 26376
rect 28123 26336 28172 26364
rect 28123 26333 28135 26336
rect 28077 26327 28135 26333
rect 28166 26324 28172 26336
rect 28224 26324 28230 26376
rect 22649 26299 22707 26305
rect 21468 26268 22094 26296
rect 22066 26240 22094 26268
rect 22649 26265 22661 26299
rect 22695 26296 22707 26299
rect 22830 26296 22836 26308
rect 22695 26268 22836 26296
rect 22695 26265 22707 26268
rect 22649 26259 22707 26265
rect 22830 26256 22836 26268
rect 22888 26296 22894 26308
rect 22888 26268 24440 26296
rect 22888 26256 22894 26268
rect 14550 26228 14556 26240
rect 14511 26200 14556 26228
rect 14550 26188 14556 26200
rect 14608 26188 14614 26240
rect 15378 26228 15384 26240
rect 15339 26200 15384 26228
rect 15378 26188 15384 26200
rect 15436 26188 15442 26240
rect 22002 26188 22008 26240
rect 22060 26228 22094 26240
rect 23290 26228 23296 26240
rect 22060 26200 23296 26228
rect 22060 26188 22066 26200
rect 23290 26188 23296 26200
rect 23348 26188 23354 26240
rect 23658 26228 23664 26240
rect 23619 26200 23664 26228
rect 23658 26188 23664 26200
rect 23716 26188 23722 26240
rect 24412 26228 24440 26268
rect 24486 26256 24492 26308
rect 24544 26296 24550 26308
rect 24642 26299 24700 26305
rect 24642 26296 24654 26299
rect 24544 26268 24654 26296
rect 24544 26256 24550 26268
rect 24642 26265 24654 26268
rect 24688 26265 24700 26299
rect 24642 26259 24700 26265
rect 25130 26228 25136 26240
rect 24412 26200 25136 26228
rect 25130 26188 25136 26200
rect 25188 26228 25194 26240
rect 25777 26231 25835 26237
rect 25777 26228 25789 26231
rect 25188 26200 25789 26228
rect 25188 26188 25194 26200
rect 25777 26197 25789 26200
rect 25823 26197 25835 26231
rect 25777 26191 25835 26197
rect 1104 26138 28888 26160
rect 1104 26086 10214 26138
rect 10266 26086 10278 26138
rect 10330 26086 10342 26138
rect 10394 26086 10406 26138
rect 10458 26086 10470 26138
rect 10522 26086 19478 26138
rect 19530 26086 19542 26138
rect 19594 26086 19606 26138
rect 19658 26086 19670 26138
rect 19722 26086 19734 26138
rect 19786 26086 28888 26138
rect 1104 26064 28888 26086
rect 15381 26027 15439 26033
rect 15381 25993 15393 26027
rect 15427 26024 15439 26027
rect 15562 26024 15568 26036
rect 15427 25996 15568 26024
rect 15427 25993 15439 25996
rect 15381 25987 15439 25993
rect 15562 25984 15568 25996
rect 15620 25984 15626 26036
rect 19150 26024 19156 26036
rect 19111 25996 19156 26024
rect 19150 25984 19156 25996
rect 19208 25984 19214 26036
rect 22649 26027 22707 26033
rect 22649 25993 22661 26027
rect 22695 26024 22707 26027
rect 22738 26024 22744 26036
rect 22695 25996 22744 26024
rect 22695 25993 22707 25996
rect 22649 25987 22707 25993
rect 22738 25984 22744 25996
rect 22796 25984 22802 26036
rect 14268 25959 14326 25965
rect 14268 25925 14280 25959
rect 14314 25956 14326 25959
rect 14550 25956 14556 25968
rect 14314 25928 14556 25956
rect 14314 25925 14326 25928
rect 14268 25919 14326 25925
rect 14550 25916 14556 25928
rect 14608 25916 14614 25968
rect 18782 25956 18788 25968
rect 17788 25928 18788 25956
rect 12526 25888 12532 25900
rect 12487 25860 12532 25888
rect 12526 25848 12532 25860
rect 12584 25848 12590 25900
rect 12710 25888 12716 25900
rect 12671 25860 12716 25888
rect 12710 25848 12716 25860
rect 12768 25848 12774 25900
rect 17788 25897 17816 25928
rect 18782 25916 18788 25928
rect 18840 25916 18846 25968
rect 18966 25916 18972 25968
rect 19024 25956 19030 25968
rect 23658 25956 23664 25968
rect 19024 25928 19288 25956
rect 19024 25916 19030 25928
rect 12897 25891 12955 25897
rect 12897 25857 12909 25891
rect 12943 25888 12955 25891
rect 13541 25891 13599 25897
rect 13541 25888 13553 25891
rect 12943 25860 13553 25888
rect 12943 25857 12955 25860
rect 12897 25851 12955 25857
rect 13541 25857 13553 25860
rect 13587 25857 13599 25891
rect 13541 25851 13599 25857
rect 17773 25891 17831 25897
rect 17773 25857 17785 25891
rect 17819 25857 17831 25891
rect 17773 25851 17831 25857
rect 17862 25848 17868 25900
rect 17920 25888 17926 25900
rect 18138 25888 18144 25900
rect 17920 25860 17965 25888
rect 18099 25860 18144 25888
rect 17920 25848 17926 25860
rect 18138 25848 18144 25860
rect 18196 25848 18202 25900
rect 19058 25888 19064 25900
rect 19019 25860 19064 25888
rect 19058 25848 19064 25860
rect 19116 25848 19122 25900
rect 19260 25897 19288 25928
rect 23308 25928 23664 25956
rect 19245 25891 19303 25897
rect 19245 25857 19257 25891
rect 19291 25888 19303 25891
rect 19334 25888 19340 25900
rect 19291 25860 19340 25888
rect 19291 25857 19303 25860
rect 19245 25851 19303 25857
rect 19334 25848 19340 25860
rect 19392 25848 19398 25900
rect 22465 25891 22523 25897
rect 22465 25857 22477 25891
rect 22511 25888 22523 25891
rect 22554 25888 22560 25900
rect 22511 25860 22560 25888
rect 22511 25857 22523 25860
rect 22465 25851 22523 25857
rect 22554 25848 22560 25860
rect 22612 25848 22618 25900
rect 23014 25848 23020 25900
rect 23072 25888 23078 25900
rect 23308 25897 23336 25928
rect 23658 25916 23664 25928
rect 23716 25916 23722 25968
rect 23750 25916 23756 25968
rect 23808 25956 23814 25968
rect 24489 25959 24547 25965
rect 24489 25956 24501 25959
rect 23808 25928 24501 25956
rect 23808 25916 23814 25928
rect 24489 25925 24501 25928
rect 24535 25925 24547 25959
rect 24489 25919 24547 25925
rect 24946 25916 24952 25968
rect 25004 25956 25010 25968
rect 26878 25956 26884 25968
rect 25004 25928 26884 25956
rect 25004 25916 25010 25928
rect 26878 25916 26884 25928
rect 26936 25956 26942 25968
rect 26936 25928 27568 25956
rect 26936 25916 26942 25928
rect 23109 25891 23167 25897
rect 23109 25888 23121 25891
rect 23072 25860 23121 25888
rect 23072 25848 23078 25860
rect 23109 25857 23121 25860
rect 23155 25857 23167 25891
rect 23109 25851 23167 25857
rect 23293 25891 23351 25897
rect 23293 25857 23305 25891
rect 23339 25857 23351 25891
rect 23293 25851 23351 25857
rect 23382 25848 23388 25900
rect 23440 25888 23446 25900
rect 23566 25897 23572 25900
rect 23523 25891 23572 25897
rect 23440 25860 23485 25888
rect 23440 25848 23446 25860
rect 23523 25857 23535 25891
rect 23569 25857 23572 25891
rect 23523 25851 23572 25857
rect 23566 25848 23572 25851
rect 23624 25888 23630 25900
rect 24213 25891 24271 25897
rect 24213 25888 24225 25891
rect 23624 25860 24225 25888
rect 23624 25848 23630 25860
rect 24213 25857 24225 25860
rect 24259 25857 24271 25891
rect 24213 25851 24271 25857
rect 24305 25891 24363 25897
rect 24305 25857 24317 25891
rect 24351 25857 24363 25891
rect 25130 25888 25136 25900
rect 25091 25860 25136 25888
rect 24305 25851 24363 25857
rect 13998 25820 14004 25832
rect 13959 25792 14004 25820
rect 13998 25780 14004 25792
rect 14056 25780 14062 25832
rect 18046 25820 18052 25832
rect 18007 25792 18052 25820
rect 18046 25780 18052 25792
rect 18104 25780 18110 25832
rect 22281 25823 22339 25829
rect 22281 25789 22293 25823
rect 22327 25820 22339 25823
rect 22646 25820 22652 25832
rect 22327 25792 22652 25820
rect 22327 25789 22339 25792
rect 22281 25783 22339 25789
rect 22646 25780 22652 25792
rect 22704 25820 22710 25832
rect 23198 25820 23204 25832
rect 22704 25792 23204 25820
rect 22704 25780 22710 25792
rect 23198 25780 23204 25792
rect 23256 25780 23262 25832
rect 24320 25820 24348 25851
rect 25130 25848 25136 25860
rect 25188 25848 25194 25900
rect 27540 25897 27568 25928
rect 27525 25891 27583 25897
rect 27525 25857 27537 25891
rect 27571 25857 27583 25891
rect 27525 25851 27583 25857
rect 24320 25792 24716 25820
rect 24688 25764 24716 25792
rect 24486 25752 24492 25764
rect 24447 25724 24492 25752
rect 24486 25712 24492 25724
rect 24544 25712 24550 25764
rect 24670 25712 24676 25764
rect 24728 25752 24734 25764
rect 25041 25755 25099 25761
rect 25041 25752 25053 25755
rect 24728 25724 25053 25752
rect 24728 25712 24734 25724
rect 25041 25721 25053 25724
rect 25087 25721 25099 25755
rect 25041 25715 25099 25721
rect 1394 25644 1400 25696
rect 1452 25684 1458 25696
rect 1489 25687 1547 25693
rect 1489 25684 1501 25687
rect 1452 25656 1501 25684
rect 1452 25644 1458 25656
rect 1489 25653 1501 25656
rect 1535 25653 1547 25687
rect 1489 25647 1547 25653
rect 13262 25644 13268 25696
rect 13320 25684 13326 25696
rect 13357 25687 13415 25693
rect 13357 25684 13369 25687
rect 13320 25656 13369 25684
rect 13320 25644 13326 25656
rect 13357 25653 13369 25656
rect 13403 25653 13415 25687
rect 13357 25647 13415 25653
rect 17589 25687 17647 25693
rect 17589 25653 17601 25687
rect 17635 25684 17647 25687
rect 17770 25684 17776 25696
rect 17635 25656 17776 25684
rect 17635 25653 17647 25656
rect 17589 25647 17647 25653
rect 17770 25644 17776 25656
rect 17828 25644 17834 25696
rect 23753 25687 23811 25693
rect 23753 25653 23765 25687
rect 23799 25684 23811 25687
rect 24946 25684 24952 25696
rect 23799 25656 24952 25684
rect 23799 25653 23811 25656
rect 23753 25647 23811 25653
rect 24946 25644 24952 25656
rect 25004 25644 25010 25696
rect 27617 25687 27675 25693
rect 27617 25653 27629 25687
rect 27663 25684 27675 25687
rect 27982 25684 27988 25696
rect 27663 25656 27988 25684
rect 27663 25653 27675 25656
rect 27617 25647 27675 25653
rect 27982 25644 27988 25656
rect 28040 25644 28046 25696
rect 1104 25594 28888 25616
rect 1104 25542 5582 25594
rect 5634 25542 5646 25594
rect 5698 25542 5710 25594
rect 5762 25542 5774 25594
rect 5826 25542 5838 25594
rect 5890 25542 14846 25594
rect 14898 25542 14910 25594
rect 14962 25542 14974 25594
rect 15026 25542 15038 25594
rect 15090 25542 15102 25594
rect 15154 25542 24110 25594
rect 24162 25542 24174 25594
rect 24226 25542 24238 25594
rect 24290 25542 24302 25594
rect 24354 25542 24366 25594
rect 24418 25542 28888 25594
rect 1104 25520 28888 25542
rect 14734 25440 14740 25492
rect 14792 25480 14798 25492
rect 14921 25483 14979 25489
rect 14921 25480 14933 25483
rect 14792 25452 14933 25480
rect 14792 25440 14798 25452
rect 14921 25449 14933 25452
rect 14967 25449 14979 25483
rect 14921 25443 14979 25449
rect 15105 25483 15163 25489
rect 15105 25449 15117 25483
rect 15151 25480 15163 25483
rect 15378 25480 15384 25492
rect 15151 25452 15384 25480
rect 15151 25449 15163 25452
rect 15105 25443 15163 25449
rect 15378 25440 15384 25452
rect 15436 25440 15442 25492
rect 22186 25480 22192 25492
rect 22147 25452 22192 25480
rect 22186 25440 22192 25452
rect 22244 25440 22250 25492
rect 22649 25483 22707 25489
rect 22649 25449 22661 25483
rect 22695 25480 22707 25483
rect 22922 25480 22928 25492
rect 22695 25452 22928 25480
rect 22695 25449 22707 25452
rect 22649 25443 22707 25449
rect 22922 25440 22928 25452
rect 22980 25440 22986 25492
rect 23566 25440 23572 25492
rect 23624 25480 23630 25492
rect 23753 25483 23811 25489
rect 23753 25480 23765 25483
rect 23624 25452 23765 25480
rect 23624 25440 23630 25452
rect 23753 25449 23765 25452
rect 23799 25449 23811 25483
rect 23753 25443 23811 25449
rect 16482 25412 16488 25424
rect 16443 25384 16488 25412
rect 16482 25372 16488 25384
rect 16540 25372 16546 25424
rect 1394 25344 1400 25356
rect 1355 25316 1400 25344
rect 1394 25304 1400 25316
rect 1452 25304 1458 25356
rect 2774 25344 2780 25356
rect 2735 25316 2780 25344
rect 2774 25304 2780 25316
rect 2832 25304 2838 25356
rect 13541 25347 13599 25353
rect 13541 25313 13553 25347
rect 13587 25344 13599 25347
rect 13998 25344 14004 25356
rect 13587 25316 14004 25344
rect 13587 25313 13599 25316
rect 13541 25307 13599 25313
rect 13998 25304 14004 25316
rect 14056 25304 14062 25356
rect 22738 25344 22744 25356
rect 21928 25316 22744 25344
rect 5534 25276 5540 25288
rect 5495 25248 5540 25276
rect 5534 25236 5540 25248
rect 5592 25236 5598 25288
rect 13262 25236 13268 25288
rect 13320 25285 13326 25288
rect 13320 25276 13332 25285
rect 13320 25248 13365 25276
rect 13320 25239 13332 25248
rect 13320 25236 13326 25239
rect 15930 25236 15936 25288
rect 15988 25276 15994 25288
rect 21928 25285 21956 25316
rect 22738 25304 22744 25316
rect 22796 25344 22802 25356
rect 22833 25347 22891 25353
rect 22833 25344 22845 25347
rect 22796 25316 22845 25344
rect 22796 25304 22802 25316
rect 22833 25313 22845 25316
rect 22879 25313 22891 25347
rect 22833 25307 22891 25313
rect 22922 25304 22928 25356
rect 22980 25344 22986 25356
rect 23106 25344 23112 25356
rect 22980 25316 23025 25344
rect 23067 25316 23112 25344
rect 22980 25304 22986 25316
rect 23106 25304 23112 25316
rect 23164 25304 23170 25356
rect 23290 25304 23296 25356
rect 23348 25344 23354 25356
rect 27522 25344 27528 25356
rect 23348 25316 23888 25344
rect 27483 25316 27528 25344
rect 23348 25304 23354 25316
rect 16301 25279 16359 25285
rect 16301 25276 16313 25279
rect 15988 25248 16313 25276
rect 15988 25236 15994 25248
rect 16301 25245 16313 25248
rect 16347 25245 16359 25279
rect 16301 25239 16359 25245
rect 21913 25279 21971 25285
rect 21913 25245 21925 25279
rect 21959 25245 21971 25279
rect 21913 25239 21971 25245
rect 22005 25279 22063 25285
rect 22005 25245 22017 25279
rect 22051 25276 22063 25279
rect 22940 25276 22968 25304
rect 22051 25248 22968 25276
rect 23017 25279 23075 25285
rect 22051 25245 22063 25248
rect 22005 25239 22063 25245
rect 23017 25245 23029 25279
rect 23063 25245 23075 25279
rect 23017 25239 23075 25245
rect 23661 25279 23719 25285
rect 23661 25245 23673 25279
rect 23707 25276 23719 25279
rect 23750 25276 23756 25288
rect 23707 25248 23756 25276
rect 23707 25245 23719 25248
rect 23661 25239 23719 25245
rect 1578 25208 1584 25220
rect 1539 25180 1584 25208
rect 1578 25168 1584 25180
rect 1636 25168 1642 25220
rect 4706 25168 4712 25220
rect 4764 25208 4770 25220
rect 4982 25208 4988 25220
rect 4764 25180 4988 25208
rect 4764 25168 4770 25180
rect 4982 25168 4988 25180
rect 5040 25168 5046 25220
rect 15289 25211 15347 25217
rect 15289 25177 15301 25211
rect 15335 25208 15347 25211
rect 15746 25208 15752 25220
rect 15335 25180 15752 25208
rect 15335 25177 15347 25180
rect 15289 25171 15347 25177
rect 15746 25168 15752 25180
rect 15804 25168 15810 25220
rect 16022 25168 16028 25220
rect 16080 25208 16086 25220
rect 16117 25211 16175 25217
rect 16117 25208 16129 25211
rect 16080 25180 16129 25208
rect 16080 25168 16086 25180
rect 16117 25177 16129 25180
rect 16163 25177 16175 25211
rect 16117 25171 16175 25177
rect 22189 25211 22247 25217
rect 22189 25177 22201 25211
rect 22235 25208 22247 25211
rect 23032 25208 23060 25239
rect 23750 25236 23756 25248
rect 23808 25236 23814 25288
rect 23860 25285 23888 25316
rect 27522 25304 27528 25316
rect 27580 25304 27586 25356
rect 27982 25344 27988 25356
rect 27943 25316 27988 25344
rect 27982 25304 27988 25316
rect 28040 25304 28046 25356
rect 28166 25344 28172 25356
rect 28127 25316 28172 25344
rect 28166 25304 28172 25316
rect 28224 25304 28230 25356
rect 23845 25279 23903 25285
rect 23845 25245 23857 25279
rect 23891 25245 23903 25279
rect 23845 25239 23903 25245
rect 24026 25236 24032 25288
rect 24084 25276 24090 25288
rect 25777 25279 25835 25285
rect 25777 25276 25789 25279
rect 24084 25248 25789 25276
rect 24084 25236 24090 25248
rect 25777 25245 25789 25248
rect 25823 25245 25835 25279
rect 25777 25239 25835 25245
rect 23474 25208 23480 25220
rect 22235 25180 23480 25208
rect 22235 25177 22247 25180
rect 22189 25171 22247 25177
rect 23474 25168 23480 25180
rect 23532 25208 23538 25220
rect 23532 25180 23980 25208
rect 23532 25168 23538 25180
rect 23952 25152 23980 25180
rect 24946 25168 24952 25220
rect 25004 25208 25010 25220
rect 25510 25211 25568 25217
rect 25510 25208 25522 25211
rect 25004 25180 25522 25208
rect 25004 25168 25010 25180
rect 25510 25177 25522 25180
rect 25556 25177 25568 25211
rect 25510 25171 25568 25177
rect 12158 25140 12164 25152
rect 12119 25112 12164 25140
rect 12158 25100 12164 25112
rect 12216 25100 12222 25152
rect 15089 25143 15147 25149
rect 15089 25109 15101 25143
rect 15135 25140 15147 25143
rect 15194 25140 15200 25152
rect 15135 25112 15200 25140
rect 15135 25109 15147 25112
rect 15089 25103 15147 25109
rect 15194 25100 15200 25112
rect 15252 25100 15258 25152
rect 15470 25100 15476 25152
rect 15528 25140 15534 25152
rect 15933 25143 15991 25149
rect 15933 25140 15945 25143
rect 15528 25112 15945 25140
rect 15528 25100 15534 25112
rect 15933 25109 15945 25112
rect 15979 25109 15991 25143
rect 16206 25140 16212 25152
rect 16167 25112 16212 25140
rect 15933 25103 15991 25109
rect 16206 25100 16212 25112
rect 16264 25100 16270 25152
rect 23934 25100 23940 25152
rect 23992 25140 23998 25152
rect 24397 25143 24455 25149
rect 24397 25140 24409 25143
rect 23992 25112 24409 25140
rect 23992 25100 23998 25112
rect 24397 25109 24409 25112
rect 24443 25109 24455 25143
rect 24397 25103 24455 25109
rect 1104 25050 28888 25072
rect 1104 24998 10214 25050
rect 10266 24998 10278 25050
rect 10330 24998 10342 25050
rect 10394 24998 10406 25050
rect 10458 24998 10470 25050
rect 10522 24998 19478 25050
rect 19530 24998 19542 25050
rect 19594 24998 19606 25050
rect 19658 24998 19670 25050
rect 19722 24998 19734 25050
rect 19786 24998 28888 25050
rect 1104 24976 28888 24998
rect 1578 24896 1584 24948
rect 1636 24936 1642 24948
rect 1765 24939 1823 24945
rect 1765 24936 1777 24939
rect 1636 24908 1777 24936
rect 1636 24896 1642 24908
rect 1765 24905 1777 24908
rect 1811 24905 1823 24939
rect 1765 24899 1823 24905
rect 12526 24896 12532 24948
rect 12584 24936 12590 24948
rect 12713 24939 12771 24945
rect 12713 24936 12725 24939
rect 12584 24908 12725 24936
rect 12584 24896 12590 24908
rect 12713 24905 12725 24908
rect 12759 24905 12771 24939
rect 12713 24899 12771 24905
rect 15194 24896 15200 24948
rect 15252 24936 15258 24948
rect 15289 24939 15347 24945
rect 15289 24936 15301 24939
rect 15252 24908 15301 24936
rect 15252 24896 15258 24908
rect 15289 24905 15301 24908
rect 15335 24905 15347 24939
rect 15289 24899 15347 24905
rect 17773 24939 17831 24945
rect 17773 24905 17785 24939
rect 17819 24936 17831 24939
rect 17862 24936 17868 24948
rect 17819 24908 17868 24936
rect 17819 24905 17831 24908
rect 17773 24899 17831 24905
rect 17862 24896 17868 24908
rect 17920 24896 17926 24948
rect 12158 24828 12164 24880
rect 12216 24868 12222 24880
rect 13081 24871 13139 24877
rect 13081 24868 13093 24871
rect 12216 24840 13093 24868
rect 12216 24828 12222 24840
rect 13081 24837 13093 24840
rect 13127 24868 13139 24871
rect 13127 24840 16712 24868
rect 13127 24837 13139 24840
rect 13081 24831 13139 24837
rect 16684 24812 16712 24840
rect 1762 24760 1768 24812
rect 1820 24800 1826 24812
rect 1857 24803 1915 24809
rect 1857 24800 1869 24803
rect 1820 24772 1869 24800
rect 1820 24760 1826 24772
rect 1857 24769 1869 24772
rect 1903 24769 1915 24803
rect 1857 24763 1915 24769
rect 4341 24803 4399 24809
rect 4341 24769 4353 24803
rect 4387 24800 4399 24803
rect 4985 24803 5043 24809
rect 4985 24800 4997 24803
rect 4387 24772 4997 24800
rect 4387 24769 4399 24772
rect 4341 24763 4399 24769
rect 4985 24769 4997 24772
rect 5031 24800 5043 24803
rect 5534 24800 5540 24812
rect 5031 24772 5540 24800
rect 5031 24769 5043 24772
rect 4985 24763 5043 24769
rect 5534 24760 5540 24772
rect 5592 24800 5598 24812
rect 5902 24800 5908 24812
rect 5592 24772 5908 24800
rect 5592 24760 5598 24772
rect 5902 24760 5908 24772
rect 5960 24800 5966 24812
rect 6365 24803 6423 24809
rect 6365 24800 6377 24803
rect 5960 24772 6377 24800
rect 5960 24760 5966 24772
rect 6365 24769 6377 24772
rect 6411 24769 6423 24803
rect 6365 24763 6423 24769
rect 15289 24803 15347 24809
rect 15289 24769 15301 24803
rect 15335 24769 15347 24803
rect 15470 24800 15476 24812
rect 15431 24772 15476 24800
rect 15289 24763 15347 24769
rect 2038 24692 2044 24744
rect 2096 24732 2102 24744
rect 4062 24732 4068 24744
rect 2096 24704 4068 24732
rect 2096 24692 2102 24704
rect 4062 24692 4068 24704
rect 4120 24692 4126 24744
rect 5169 24735 5227 24741
rect 5169 24701 5181 24735
rect 5215 24701 5227 24735
rect 5169 24695 5227 24701
rect 6549 24735 6607 24741
rect 6549 24701 6561 24735
rect 6595 24701 6607 24735
rect 13170 24732 13176 24744
rect 13131 24704 13176 24732
rect 6549 24695 6607 24701
rect 3142 24624 3148 24676
rect 3200 24664 3206 24676
rect 5184 24664 5212 24695
rect 3200 24636 5212 24664
rect 6564 24664 6592 24695
rect 13170 24692 13176 24704
rect 13228 24692 13234 24744
rect 13354 24732 13360 24744
rect 13315 24704 13360 24732
rect 13354 24692 13360 24704
rect 13412 24692 13418 24744
rect 15304 24732 15332 24763
rect 15470 24760 15476 24772
rect 15528 24760 15534 24812
rect 16666 24800 16672 24812
rect 16579 24772 16672 24800
rect 16666 24760 16672 24772
rect 16724 24760 16730 24812
rect 17402 24760 17408 24812
rect 17460 24800 17466 24812
rect 17589 24803 17647 24809
rect 17589 24800 17601 24803
rect 17460 24772 17601 24800
rect 17460 24760 17466 24772
rect 17589 24769 17601 24772
rect 17635 24769 17647 24803
rect 17589 24763 17647 24769
rect 17678 24760 17684 24812
rect 17736 24800 17742 24812
rect 17736 24772 17781 24800
rect 17736 24760 17742 24772
rect 17862 24760 17868 24812
rect 17920 24800 17926 24812
rect 18877 24803 18935 24809
rect 18877 24800 18889 24803
rect 17920 24772 18889 24800
rect 17920 24760 17926 24772
rect 18877 24769 18889 24772
rect 18923 24769 18935 24803
rect 18877 24763 18935 24769
rect 21269 24803 21327 24809
rect 21269 24769 21281 24803
rect 21315 24800 21327 24803
rect 25038 24800 25044 24812
rect 21315 24772 25044 24800
rect 21315 24769 21327 24772
rect 21269 24763 21327 24769
rect 25038 24760 25044 24772
rect 25096 24760 25102 24812
rect 26418 24760 26424 24812
rect 26476 24800 26482 24812
rect 26476 24772 26521 24800
rect 26476 24760 26482 24772
rect 26786 24760 26792 24812
rect 26844 24800 26850 24812
rect 26973 24803 27031 24809
rect 26973 24800 26985 24803
rect 26844 24772 26985 24800
rect 26844 24760 26850 24772
rect 26973 24769 26985 24772
rect 27019 24769 27031 24803
rect 26973 24763 27031 24769
rect 27709 24803 27767 24809
rect 27709 24769 27721 24803
rect 27755 24800 27767 24803
rect 27755 24772 27936 24800
rect 27755 24769 27767 24772
rect 27709 24763 27767 24769
rect 16574 24732 16580 24744
rect 15304 24704 16580 24732
rect 16574 24692 16580 24704
rect 16632 24732 16638 24744
rect 16942 24732 16948 24744
rect 16632 24704 16948 24732
rect 16632 24692 16638 24704
rect 16942 24692 16948 24704
rect 17000 24692 17006 24744
rect 17310 24692 17316 24744
rect 17368 24732 17374 24744
rect 18049 24735 18107 24741
rect 18049 24732 18061 24735
rect 17368 24704 18061 24732
rect 17368 24692 17374 24704
rect 18049 24701 18061 24704
rect 18095 24701 18107 24735
rect 21818 24732 21824 24744
rect 21779 24704 21824 24732
rect 18049 24695 18107 24701
rect 21818 24692 21824 24704
rect 21876 24692 21882 24744
rect 22094 24692 22100 24744
rect 22152 24732 22158 24744
rect 25958 24732 25964 24744
rect 22152 24704 22197 24732
rect 25919 24704 25964 24732
rect 22152 24692 22158 24704
rect 25958 24692 25964 24704
rect 26016 24692 26022 24744
rect 26237 24735 26295 24741
rect 26237 24701 26249 24735
rect 26283 24732 26295 24735
rect 27801 24735 27859 24741
rect 27801 24732 27813 24735
rect 26283 24704 27813 24732
rect 26283 24701 26295 24704
rect 26237 24695 26295 24701
rect 27801 24701 27813 24704
rect 27847 24701 27859 24735
rect 27801 24695 27859 24701
rect 27908 24664 27936 24772
rect 28258 24664 28264 24676
rect 6564 24636 28264 24664
rect 3200 24624 3206 24636
rect 1762 24556 1768 24608
rect 1820 24596 1826 24608
rect 6564 24596 6592 24636
rect 28258 24624 28264 24636
rect 28316 24624 28322 24676
rect 1820 24568 6592 24596
rect 1820 24556 1826 24568
rect 16574 24556 16580 24608
rect 16632 24596 16638 24608
rect 16761 24599 16819 24605
rect 16761 24596 16773 24599
rect 16632 24568 16773 24596
rect 16632 24556 16638 24568
rect 16761 24565 16773 24568
rect 16807 24565 16819 24599
rect 16761 24559 16819 24565
rect 17129 24599 17187 24605
rect 17129 24565 17141 24599
rect 17175 24596 17187 24599
rect 17310 24596 17316 24608
rect 17175 24568 17316 24596
rect 17175 24565 17187 24568
rect 17129 24559 17187 24565
rect 17310 24556 17316 24568
rect 17368 24556 17374 24608
rect 18874 24556 18880 24608
rect 18932 24596 18938 24608
rect 18969 24599 19027 24605
rect 18969 24596 18981 24599
rect 18932 24568 18981 24596
rect 18932 24556 18938 24568
rect 18969 24565 18981 24568
rect 19015 24565 19027 24599
rect 19978 24596 19984 24608
rect 19939 24568 19984 24596
rect 18969 24559 19027 24565
rect 19978 24556 19984 24568
rect 20036 24556 20042 24608
rect 27157 24599 27215 24605
rect 27157 24565 27169 24599
rect 27203 24596 27215 24599
rect 27430 24596 27436 24608
rect 27203 24568 27436 24596
rect 27203 24565 27215 24568
rect 27157 24559 27215 24565
rect 27430 24556 27436 24568
rect 27488 24556 27494 24608
rect 1104 24506 28888 24528
rect 1104 24454 5582 24506
rect 5634 24454 5646 24506
rect 5698 24454 5710 24506
rect 5762 24454 5774 24506
rect 5826 24454 5838 24506
rect 5890 24454 14846 24506
rect 14898 24454 14910 24506
rect 14962 24454 14974 24506
rect 15026 24454 15038 24506
rect 15090 24454 15102 24506
rect 15154 24454 24110 24506
rect 24162 24454 24174 24506
rect 24226 24454 24238 24506
rect 24290 24454 24302 24506
rect 24354 24454 24366 24506
rect 24418 24454 28888 24506
rect 1104 24432 28888 24454
rect 15933 24395 15991 24401
rect 15933 24361 15945 24395
rect 15979 24361 15991 24395
rect 16666 24392 16672 24404
rect 16627 24364 16672 24392
rect 15933 24355 15991 24361
rect 15948 24324 15976 24355
rect 16666 24352 16672 24364
rect 16724 24352 16730 24404
rect 19429 24395 19487 24401
rect 19429 24361 19441 24395
rect 19475 24392 19487 24395
rect 19886 24392 19892 24404
rect 19475 24364 19892 24392
rect 19475 24361 19487 24364
rect 19429 24355 19487 24361
rect 16206 24324 16212 24336
rect 15948 24296 16212 24324
rect 16206 24284 16212 24296
rect 16264 24324 16270 24336
rect 16264 24296 16620 24324
rect 16264 24284 16270 24296
rect 16592 24200 16620 24296
rect 18601 24259 18659 24265
rect 18601 24225 18613 24259
rect 18647 24256 18659 24259
rect 19444 24256 19472 24355
rect 19886 24352 19892 24364
rect 19944 24352 19950 24404
rect 22281 24395 22339 24401
rect 22281 24361 22293 24395
rect 22327 24392 22339 24395
rect 23014 24392 23020 24404
rect 22327 24364 23020 24392
rect 22327 24361 22339 24364
rect 22281 24355 22339 24361
rect 23014 24352 23020 24364
rect 23072 24352 23078 24404
rect 18647 24228 19472 24256
rect 20809 24259 20867 24265
rect 18647 24225 18659 24228
rect 18601 24219 18659 24225
rect 20809 24225 20821 24259
rect 20855 24256 20867 24259
rect 24026 24256 24032 24268
rect 20855 24228 24032 24256
rect 20855 24225 20867 24228
rect 20809 24219 20867 24225
rect 24026 24216 24032 24228
rect 24084 24216 24090 24268
rect 27522 24256 27528 24268
rect 27483 24228 27528 24256
rect 27522 24216 27528 24228
rect 27580 24216 27586 24268
rect 1394 24188 1400 24200
rect 1355 24160 1400 24188
rect 1394 24148 1400 24160
rect 1452 24148 1458 24200
rect 4985 24191 5043 24197
rect 4985 24157 4997 24191
rect 5031 24188 5043 24191
rect 5902 24188 5908 24200
rect 5031 24160 5908 24188
rect 5031 24157 5043 24160
rect 4985 24151 5043 24157
rect 5902 24148 5908 24160
rect 5960 24148 5966 24200
rect 12161 24191 12219 24197
rect 12161 24157 12173 24191
rect 12207 24188 12219 24191
rect 12894 24188 12900 24200
rect 12207 24160 12900 24188
rect 12207 24157 12219 24160
rect 12161 24151 12219 24157
rect 12894 24148 12900 24160
rect 12952 24148 12958 24200
rect 15286 24188 15292 24200
rect 15247 24160 15292 24188
rect 15286 24148 15292 24160
rect 15344 24148 15350 24200
rect 16574 24188 16580 24200
rect 16535 24160 16580 24188
rect 16574 24148 16580 24160
rect 16632 24148 16638 24200
rect 18325 24191 18383 24197
rect 18325 24157 18337 24191
rect 18371 24157 18383 24191
rect 18325 24151 18383 24157
rect 5442 24120 5448 24132
rect 5403 24092 5448 24120
rect 5442 24080 5448 24092
rect 5500 24080 5506 24132
rect 16117 24123 16175 24129
rect 16117 24089 16129 24123
rect 16163 24120 16175 24123
rect 16850 24120 16856 24132
rect 16163 24092 16856 24120
rect 16163 24089 16175 24092
rect 16117 24083 16175 24089
rect 16850 24080 16856 24092
rect 16908 24120 16914 24132
rect 18340 24120 18368 24151
rect 19058 24148 19064 24200
rect 19116 24188 19122 24200
rect 21269 24191 21327 24197
rect 21269 24188 21281 24191
rect 19116 24160 21281 24188
rect 19116 24148 19122 24160
rect 21269 24157 21281 24160
rect 21315 24188 21327 24191
rect 21818 24188 21824 24200
rect 21315 24160 21824 24188
rect 21315 24157 21327 24160
rect 21269 24151 21327 24157
rect 21818 24148 21824 24160
rect 21876 24148 21882 24200
rect 25869 24191 25927 24197
rect 25869 24157 25881 24191
rect 25915 24157 25927 24191
rect 25869 24151 25927 24157
rect 16908 24092 18368 24120
rect 16908 24080 16914 24092
rect 20254 24080 20260 24132
rect 20312 24120 20318 24132
rect 20542 24123 20600 24129
rect 20542 24120 20554 24123
rect 20312 24092 20554 24120
rect 20312 24080 20318 24092
rect 20542 24089 20554 24092
rect 20588 24089 20600 24123
rect 22370 24120 22376 24132
rect 22331 24092 22376 24120
rect 20542 24083 20600 24089
rect 22370 24080 22376 24092
rect 22428 24080 22434 24132
rect 25038 24120 25044 24132
rect 24999 24092 25044 24120
rect 25038 24080 25044 24092
rect 25096 24080 25102 24132
rect 25590 24080 25596 24132
rect 25648 24120 25654 24132
rect 25884 24120 25912 24151
rect 28166 24148 28172 24200
rect 28224 24188 28230 24200
rect 28224 24160 28269 24188
rect 28224 24148 28230 24160
rect 27430 24120 27436 24132
rect 25648 24092 27436 24120
rect 25648 24080 25654 24092
rect 27430 24080 27436 24092
rect 27488 24080 27494 24132
rect 27982 24120 27988 24132
rect 27943 24092 27988 24120
rect 27982 24080 27988 24092
rect 28040 24080 28046 24132
rect 1578 24052 1584 24064
rect 1539 24024 1584 24052
rect 1578 24012 1584 24024
rect 1636 24012 1642 24064
rect 12345 24055 12403 24061
rect 12345 24021 12357 24055
rect 12391 24052 12403 24055
rect 12434 24052 12440 24064
rect 12391 24024 12440 24052
rect 12391 24021 12403 24024
rect 12345 24015 12403 24021
rect 12434 24012 12440 24024
rect 12492 24012 12498 24064
rect 15102 24052 15108 24064
rect 15063 24024 15108 24052
rect 15102 24012 15108 24024
rect 15160 24012 15166 24064
rect 15654 24012 15660 24064
rect 15712 24052 15718 24064
rect 15749 24055 15807 24061
rect 15749 24052 15761 24055
rect 15712 24024 15761 24052
rect 15712 24012 15718 24024
rect 15749 24021 15761 24024
rect 15795 24021 15807 24055
rect 15749 24015 15807 24021
rect 15917 24055 15975 24061
rect 15917 24021 15929 24055
rect 15963 24052 15975 24055
rect 16022 24052 16028 24064
rect 15963 24024 16028 24052
rect 15963 24021 15975 24024
rect 15917 24015 15975 24021
rect 16022 24012 16028 24024
rect 16080 24052 16086 24064
rect 16758 24052 16764 24064
rect 16080 24024 16764 24052
rect 16080 24012 16086 24024
rect 16758 24012 16764 24024
rect 16816 24012 16822 24064
rect 17037 24055 17095 24061
rect 17037 24021 17049 24055
rect 17083 24052 17095 24055
rect 17402 24052 17408 24064
rect 17083 24024 17408 24052
rect 17083 24021 17095 24024
rect 17037 24015 17095 24021
rect 17402 24012 17408 24024
rect 17460 24012 17466 24064
rect 21450 24052 21456 24064
rect 21411 24024 21456 24052
rect 21450 24012 21456 24024
rect 21508 24012 21514 24064
rect 1104 23962 28888 23984
rect 1104 23910 10214 23962
rect 10266 23910 10278 23962
rect 10330 23910 10342 23962
rect 10394 23910 10406 23962
rect 10458 23910 10470 23962
rect 10522 23910 19478 23962
rect 19530 23910 19542 23962
rect 19594 23910 19606 23962
rect 19658 23910 19670 23962
rect 19722 23910 19734 23962
rect 19786 23910 28888 23962
rect 1104 23888 28888 23910
rect 1578 23808 1584 23860
rect 1636 23848 1642 23860
rect 13170 23848 13176 23860
rect 1636 23820 13176 23848
rect 1636 23808 1642 23820
rect 13170 23808 13176 23820
rect 13228 23808 13234 23860
rect 17589 23851 17647 23857
rect 17589 23817 17601 23851
rect 17635 23848 17647 23851
rect 17678 23848 17684 23860
rect 17635 23820 17684 23848
rect 17635 23817 17647 23820
rect 17589 23811 17647 23817
rect 17678 23808 17684 23820
rect 17736 23808 17742 23860
rect 17862 23808 17868 23860
rect 17920 23848 17926 23860
rect 18509 23851 18567 23857
rect 18509 23848 18521 23851
rect 17920 23820 18521 23848
rect 17920 23808 17926 23820
rect 18509 23817 18521 23820
rect 18555 23817 18567 23851
rect 18509 23811 18567 23817
rect 21358 23808 21364 23860
rect 21416 23848 21422 23860
rect 22370 23848 22376 23860
rect 21416 23820 22376 23848
rect 21416 23808 21422 23820
rect 22370 23808 22376 23820
rect 22428 23848 22434 23860
rect 22428 23820 22876 23848
rect 22428 23808 22434 23820
rect 2314 23740 2320 23792
rect 2372 23780 2378 23792
rect 4893 23783 4951 23789
rect 4893 23780 4905 23783
rect 2372 23752 4905 23780
rect 2372 23740 2378 23752
rect 4893 23749 4905 23752
rect 4939 23749 4951 23783
rect 4893 23743 4951 23749
rect 15004 23783 15062 23789
rect 15004 23749 15016 23783
rect 15050 23780 15062 23783
rect 15102 23780 15108 23792
rect 15050 23752 15108 23780
rect 15050 23749 15062 23752
rect 15004 23743 15062 23749
rect 15102 23740 15108 23752
rect 15160 23740 15166 23792
rect 4709 23715 4767 23721
rect 4709 23681 4721 23715
rect 4755 23712 4767 23715
rect 5902 23712 5908 23724
rect 4755 23684 5908 23712
rect 4755 23681 4767 23684
rect 4709 23675 4767 23681
rect 5902 23672 5908 23684
rect 5960 23672 5966 23724
rect 12621 23715 12679 23721
rect 12621 23681 12633 23715
rect 12667 23712 12679 23715
rect 13538 23712 13544 23724
rect 12667 23684 13544 23712
rect 12667 23681 12679 23684
rect 12621 23675 12679 23681
rect 13538 23672 13544 23684
rect 13596 23712 13602 23724
rect 13596 23684 16712 23712
rect 13596 23672 13602 23684
rect 9490 23604 9496 23656
rect 9548 23644 9554 23656
rect 12713 23647 12771 23653
rect 12713 23644 12725 23647
rect 9548 23616 12725 23644
rect 9548 23604 9554 23616
rect 12713 23613 12725 23616
rect 12759 23613 12771 23647
rect 12713 23607 12771 23613
rect 12802 23604 12808 23656
rect 12860 23644 12866 23656
rect 12897 23647 12955 23653
rect 12897 23644 12909 23647
rect 12860 23616 12909 23644
rect 12860 23604 12866 23616
rect 12897 23613 12909 23616
rect 12943 23644 12955 23647
rect 13354 23644 13360 23656
rect 12943 23616 13360 23644
rect 12943 23613 12955 23616
rect 12897 23607 12955 23613
rect 13354 23604 13360 23616
rect 13412 23604 13418 23656
rect 14734 23644 14740 23656
rect 14695 23616 14740 23644
rect 14734 23604 14740 23616
rect 14792 23604 14798 23656
rect 3142 23468 3148 23520
rect 3200 23508 3206 23520
rect 4154 23508 4160 23520
rect 3200 23480 4160 23508
rect 3200 23468 3206 23480
rect 4154 23468 4160 23480
rect 4212 23468 4218 23520
rect 12253 23511 12311 23517
rect 12253 23477 12265 23511
rect 12299 23508 12311 23511
rect 12526 23508 12532 23520
rect 12299 23480 12532 23508
rect 12299 23477 12311 23480
rect 12253 23471 12311 23477
rect 12526 23468 12532 23480
rect 12584 23468 12590 23520
rect 16117 23511 16175 23517
rect 16117 23477 16129 23511
rect 16163 23508 16175 23511
rect 16574 23508 16580 23520
rect 16163 23480 16580 23508
rect 16163 23477 16175 23480
rect 16117 23471 16175 23477
rect 16574 23468 16580 23480
rect 16632 23468 16638 23520
rect 16684 23508 16712 23684
rect 16758 23672 16764 23724
rect 16816 23712 16822 23724
rect 17126 23712 17132 23724
rect 16816 23684 17132 23712
rect 16816 23672 16822 23684
rect 17126 23672 17132 23684
rect 17184 23712 17190 23724
rect 17880 23712 17908 23808
rect 21726 23740 21732 23792
rect 21784 23780 21790 23792
rect 21821 23783 21879 23789
rect 21821 23780 21833 23783
rect 21784 23752 21833 23780
rect 21784 23740 21790 23752
rect 21821 23749 21833 23752
rect 21867 23749 21879 23783
rect 21821 23743 21879 23749
rect 21910 23740 21916 23792
rect 21968 23780 21974 23792
rect 22848 23789 22876 23820
rect 27614 23808 27620 23860
rect 27672 23848 27678 23860
rect 27709 23851 27767 23857
rect 27709 23848 27721 23851
rect 27672 23820 27721 23848
rect 27672 23808 27678 23820
rect 27709 23817 27721 23820
rect 27755 23817 27767 23851
rect 27709 23811 27767 23817
rect 22021 23783 22079 23789
rect 22021 23780 22033 23783
rect 21968 23752 22033 23780
rect 21968 23740 21974 23752
rect 22021 23749 22033 23752
rect 22067 23749 22079 23783
rect 22021 23743 22079 23749
rect 22833 23783 22891 23789
rect 22833 23749 22845 23783
rect 22879 23749 22891 23783
rect 27430 23780 27436 23792
rect 27391 23752 27436 23780
rect 22833 23743 22891 23749
rect 27430 23740 27436 23752
rect 27488 23740 27494 23792
rect 17184 23684 17908 23712
rect 19633 23715 19691 23721
rect 17184 23672 17190 23684
rect 19633 23681 19645 23715
rect 19679 23712 19691 23715
rect 19794 23712 19800 23724
rect 19679 23684 19800 23712
rect 19679 23681 19691 23684
rect 19633 23675 19691 23681
rect 19794 23672 19800 23684
rect 19852 23672 19858 23724
rect 20806 23712 20812 23724
rect 20767 23684 20812 23712
rect 20806 23672 20812 23684
rect 20864 23672 20870 23724
rect 21177 23715 21235 23721
rect 21177 23681 21189 23715
rect 21223 23712 21235 23715
rect 21450 23712 21456 23724
rect 21223 23684 21456 23712
rect 21223 23681 21235 23684
rect 21177 23675 21235 23681
rect 21450 23672 21456 23684
rect 21508 23712 21514 23724
rect 21928 23712 21956 23740
rect 25590 23712 25596 23724
rect 21508 23684 21956 23712
rect 25551 23684 25596 23712
rect 21508 23672 21514 23684
rect 25590 23672 25596 23684
rect 25648 23672 25654 23724
rect 19889 23647 19947 23653
rect 19889 23613 19901 23647
rect 19935 23644 19947 23647
rect 20714 23644 20720 23656
rect 19935 23616 20720 23644
rect 19935 23613 19947 23616
rect 19889 23607 19947 23613
rect 20714 23604 20720 23616
rect 20772 23604 20778 23656
rect 22002 23604 22008 23656
rect 22060 23644 22066 23656
rect 22060 23616 22140 23644
rect 22060 23604 22066 23616
rect 20530 23536 20536 23588
rect 20588 23576 20594 23588
rect 21818 23576 21824 23588
rect 20588 23548 21824 23576
rect 20588 23536 20594 23548
rect 21818 23536 21824 23548
rect 21876 23576 21882 23588
rect 22112 23576 22140 23616
rect 25406 23604 25412 23656
rect 25464 23644 25470 23656
rect 26145 23647 26203 23653
rect 26145 23644 26157 23647
rect 25464 23616 26157 23644
rect 25464 23604 25470 23616
rect 26145 23613 26157 23616
rect 26191 23644 26203 23647
rect 27062 23644 27068 23656
rect 26191 23616 27068 23644
rect 26191 23613 26203 23616
rect 26145 23607 26203 23613
rect 27062 23604 27068 23616
rect 27120 23604 27126 23656
rect 22649 23579 22707 23585
rect 22649 23576 22661 23579
rect 21876 23548 22661 23576
rect 21876 23536 21882 23548
rect 22649 23545 22661 23548
rect 22695 23545 22707 23579
rect 22649 23539 22707 23545
rect 17221 23511 17279 23517
rect 17221 23508 17233 23511
rect 16684 23480 17233 23508
rect 17221 23477 17233 23480
rect 17267 23508 17279 23511
rect 18138 23508 18144 23520
rect 17267 23480 18144 23508
rect 17267 23477 17279 23480
rect 17221 23471 17279 23477
rect 18138 23468 18144 23480
rect 18196 23468 18202 23520
rect 20070 23468 20076 23520
rect 20128 23508 20134 23520
rect 20625 23511 20683 23517
rect 20625 23508 20637 23511
rect 20128 23480 20637 23508
rect 20128 23468 20134 23480
rect 20625 23477 20637 23480
rect 20671 23477 20683 23511
rect 20625 23471 20683 23477
rect 21085 23511 21143 23517
rect 21085 23477 21097 23511
rect 21131 23508 21143 23511
rect 21542 23508 21548 23520
rect 21131 23480 21548 23508
rect 21131 23477 21143 23480
rect 21085 23471 21143 23477
rect 21542 23468 21548 23480
rect 21600 23468 21606 23520
rect 21634 23468 21640 23520
rect 21692 23508 21698 23520
rect 22005 23511 22063 23517
rect 22005 23508 22017 23511
rect 21692 23480 22017 23508
rect 21692 23468 21698 23480
rect 22005 23477 22017 23480
rect 22051 23477 22063 23511
rect 22005 23471 22063 23477
rect 22094 23468 22100 23520
rect 22152 23508 22158 23520
rect 22189 23511 22247 23517
rect 22189 23508 22201 23511
rect 22152 23480 22201 23508
rect 22152 23468 22158 23480
rect 22189 23477 22201 23480
rect 22235 23477 22247 23511
rect 22189 23471 22247 23477
rect 1104 23418 28888 23440
rect 1104 23366 5582 23418
rect 5634 23366 5646 23418
rect 5698 23366 5710 23418
rect 5762 23366 5774 23418
rect 5826 23366 5838 23418
rect 5890 23366 14846 23418
rect 14898 23366 14910 23418
rect 14962 23366 14974 23418
rect 15026 23366 15038 23418
rect 15090 23366 15102 23418
rect 15154 23366 24110 23418
rect 24162 23366 24174 23418
rect 24226 23366 24238 23418
rect 24290 23366 24302 23418
rect 24354 23366 24366 23418
rect 24418 23366 28888 23418
rect 1104 23344 28888 23366
rect 13538 23304 13544 23316
rect 13499 23276 13544 23304
rect 13538 23264 13544 23276
rect 13596 23264 13602 23316
rect 15286 23264 15292 23316
rect 15344 23304 15350 23316
rect 15381 23307 15439 23313
rect 15381 23304 15393 23307
rect 15344 23276 15393 23304
rect 15344 23264 15350 23276
rect 15381 23273 15393 23276
rect 15427 23273 15439 23307
rect 15381 23267 15439 23273
rect 15565 23307 15623 23313
rect 15565 23273 15577 23307
rect 15611 23304 15623 23307
rect 16666 23304 16672 23316
rect 15611 23276 16672 23304
rect 15611 23273 15623 23276
rect 15565 23267 15623 23273
rect 16666 23264 16672 23276
rect 16724 23264 16730 23316
rect 17497 23307 17555 23313
rect 17497 23273 17509 23307
rect 17543 23304 17555 23307
rect 17678 23304 17684 23316
rect 17543 23276 17684 23304
rect 17543 23273 17555 23276
rect 17497 23267 17555 23273
rect 17678 23264 17684 23276
rect 17736 23264 17742 23316
rect 19794 23264 19800 23316
rect 19852 23304 19858 23316
rect 19889 23307 19947 23313
rect 19889 23304 19901 23307
rect 19852 23276 19901 23304
rect 19852 23264 19858 23276
rect 19889 23273 19901 23276
rect 19935 23273 19947 23307
rect 19889 23267 19947 23273
rect 20809 23307 20867 23313
rect 20809 23273 20821 23307
rect 20855 23304 20867 23307
rect 21082 23304 21088 23316
rect 20855 23276 21088 23304
rect 20855 23273 20867 23276
rect 20809 23267 20867 23273
rect 21082 23264 21088 23276
rect 21140 23264 21146 23316
rect 21266 23264 21272 23316
rect 21324 23304 21330 23316
rect 21637 23307 21695 23313
rect 21637 23304 21649 23307
rect 21324 23276 21649 23304
rect 21324 23264 21330 23276
rect 21637 23273 21649 23276
rect 21683 23273 21695 23307
rect 26970 23304 26976 23316
rect 21637 23267 21695 23273
rect 22066 23276 26976 23304
rect 15654 23196 15660 23248
rect 15712 23236 15718 23248
rect 15933 23239 15991 23245
rect 15933 23236 15945 23239
rect 15712 23208 15945 23236
rect 15712 23196 15718 23208
rect 15933 23205 15945 23208
rect 15979 23205 15991 23239
rect 18414 23236 18420 23248
rect 18375 23208 18420 23236
rect 15933 23199 15991 23205
rect 18414 23196 18420 23208
rect 18472 23196 18478 23248
rect 22066 23236 22094 23276
rect 26970 23264 26976 23276
rect 27028 23264 27034 23316
rect 27982 23304 27988 23316
rect 27943 23276 27988 23304
rect 27982 23264 27988 23276
rect 28040 23264 28046 23316
rect 18524 23208 22094 23236
rect 23109 23239 23167 23245
rect 18524 23168 18552 23208
rect 23109 23205 23121 23239
rect 23155 23205 23167 23239
rect 23109 23199 23167 23205
rect 24857 23239 24915 23245
rect 24857 23205 24869 23239
rect 24903 23236 24915 23239
rect 25222 23236 25228 23248
rect 24903 23208 25228 23236
rect 24903 23205 24915 23208
rect 24857 23199 24915 23205
rect 20530 23168 20536 23180
rect 14844 23140 18552 23168
rect 19444 23140 20536 23168
rect 12158 23100 12164 23112
rect 12119 23072 12164 23100
rect 12158 23060 12164 23072
rect 12216 23060 12222 23112
rect 12434 23109 12440 23112
rect 12428 23063 12440 23109
rect 12492 23100 12498 23112
rect 12492 23072 12528 23100
rect 12434 23060 12440 23063
rect 12492 23060 12498 23072
rect 12176 23032 12204 23060
rect 14734 23032 14740 23044
rect 12176 23004 14740 23032
rect 14734 22992 14740 23004
rect 14792 22992 14798 23044
rect 12618 22924 12624 22976
rect 12676 22964 12682 22976
rect 14844 22964 14872 23140
rect 16574 23100 16580 23112
rect 16535 23072 16580 23100
rect 16574 23060 16580 23072
rect 16632 23060 16638 23112
rect 16853 23103 16911 23109
rect 16853 23069 16865 23103
rect 16899 23100 16911 23103
rect 17126 23100 17132 23112
rect 16899 23072 17132 23100
rect 16899 23069 16911 23072
rect 16853 23063 16911 23069
rect 17126 23060 17132 23072
rect 17184 23060 17190 23112
rect 18138 23100 18144 23112
rect 18099 23072 18144 23100
rect 18138 23060 18144 23072
rect 18196 23060 18202 23112
rect 18233 23103 18291 23109
rect 18233 23069 18245 23103
rect 18279 23100 18291 23103
rect 18279 23072 18920 23100
rect 18279 23069 18291 23072
rect 18233 23063 18291 23069
rect 18892 23044 18920 23072
rect 18966 23060 18972 23112
rect 19024 23100 19030 23112
rect 19444 23109 19472 23140
rect 20530 23128 20536 23140
rect 20588 23128 20594 23180
rect 20806 23168 20812 23180
rect 20640 23140 20812 23168
rect 19245 23103 19303 23109
rect 19245 23100 19257 23103
rect 19024 23072 19257 23100
rect 19024 23060 19030 23072
rect 19245 23069 19257 23072
rect 19291 23069 19303 23103
rect 19245 23063 19303 23069
rect 19429 23103 19487 23109
rect 19429 23069 19441 23103
rect 19475 23069 19487 23103
rect 19429 23063 19487 23069
rect 19521 23103 19579 23109
rect 19521 23069 19533 23103
rect 19567 23069 19579 23103
rect 19521 23063 19579 23069
rect 19613 23103 19671 23109
rect 19613 23069 19625 23103
rect 19659 23100 19671 23103
rect 20438 23100 20444 23112
rect 19659 23072 20444 23100
rect 19659 23069 19671 23072
rect 19613 23063 19671 23069
rect 16758 23032 16764 23044
rect 16671 23004 16764 23032
rect 16758 22992 16764 23004
rect 16816 23032 16822 23044
rect 16942 23032 16948 23044
rect 16816 23004 16948 23032
rect 16816 22992 16822 23004
rect 16942 22992 16948 23004
rect 17000 22992 17006 23044
rect 17310 23032 17316 23044
rect 17271 23004 17316 23032
rect 17310 22992 17316 23004
rect 17368 22992 17374 23044
rect 17402 22992 17408 23044
rect 17460 23032 17466 23044
rect 17513 23035 17571 23041
rect 17513 23032 17525 23035
rect 17460 23004 17525 23032
rect 17460 22992 17466 23004
rect 17513 23001 17525 23004
rect 17559 23001 17571 23035
rect 17513 22995 17571 23001
rect 18417 23035 18475 23041
rect 18417 23001 18429 23035
rect 18463 23032 18475 23035
rect 18782 23032 18788 23044
rect 18463 23004 18788 23032
rect 18463 23001 18475 23004
rect 18417 22995 18475 23001
rect 18782 22992 18788 23004
rect 18840 22992 18846 23044
rect 18874 22992 18880 23044
rect 18932 23032 18938 23044
rect 19536 23032 19564 23063
rect 20438 23060 20444 23072
rect 20496 23060 20502 23112
rect 20640 23041 20668 23140
rect 20806 23128 20812 23140
rect 20864 23168 20870 23180
rect 21450 23168 21456 23180
rect 20864 23140 21456 23168
rect 20864 23128 20870 23140
rect 21450 23128 21456 23140
rect 21508 23128 21514 23180
rect 21818 23128 21824 23180
rect 21876 23168 21882 23180
rect 22281 23171 22339 23177
rect 22281 23168 22293 23171
rect 21876 23140 22293 23168
rect 21876 23128 21882 23140
rect 22281 23137 22293 23140
rect 22327 23137 22339 23171
rect 22281 23131 22339 23137
rect 22465 23103 22523 23109
rect 21376 23072 21680 23100
rect 18932 23004 19564 23032
rect 20625 23035 20683 23041
rect 18932 22992 18938 23004
rect 20625 23001 20637 23035
rect 20671 23001 20683 23035
rect 20625 22995 20683 23001
rect 20841 23035 20899 23041
rect 20841 23001 20853 23035
rect 20887 23032 20899 23035
rect 21376 23032 21404 23072
rect 20887 23004 21404 23032
rect 20887 23001 20899 23004
rect 20841 22995 20899 23001
rect 21450 22992 21456 23044
rect 21508 23032 21514 23044
rect 21652 23041 21680 23072
rect 22465 23069 22477 23103
rect 22511 23100 22523 23103
rect 23124 23100 23152 23199
rect 25222 23196 25228 23208
rect 25280 23196 25286 23248
rect 27706 23196 27712 23248
rect 27764 23236 27770 23248
rect 28442 23236 28448 23248
rect 27764 23208 28448 23236
rect 27764 23196 27770 23208
rect 28442 23196 28448 23208
rect 28500 23196 28506 23248
rect 23658 23168 23664 23180
rect 23619 23140 23664 23168
rect 23658 23128 23664 23140
rect 23716 23168 23722 23180
rect 23716 23140 24624 23168
rect 23716 23128 23722 23140
rect 22511 23072 23152 23100
rect 22511 23069 22523 23072
rect 22465 23063 22523 23069
rect 23382 23060 23388 23112
rect 23440 23100 23446 23112
rect 24596 23109 24624 23140
rect 25866 23128 25872 23180
rect 25924 23168 25930 23180
rect 25924 23140 27936 23168
rect 25924 23128 25930 23140
rect 24581 23103 24639 23109
rect 23440 23072 23704 23100
rect 23440 23060 23446 23072
rect 21652 23035 21727 23041
rect 21508 23004 21553 23032
rect 21652 23004 21681 23035
rect 21508 22992 21514 23004
rect 21669 23001 21681 23004
rect 21715 23032 21727 23035
rect 21910 23032 21916 23044
rect 21715 23004 21916 23032
rect 21715 23001 21727 23004
rect 21669 22995 21727 23001
rect 21910 22992 21916 23004
rect 21968 22992 21974 23044
rect 22554 22992 22560 23044
rect 22612 23032 22618 23044
rect 23569 23035 23627 23041
rect 23569 23032 23581 23035
rect 22612 23004 23581 23032
rect 22612 22992 22618 23004
rect 23569 23001 23581 23004
rect 23615 23001 23627 23035
rect 23676 23032 23704 23072
rect 24581 23069 24593 23103
rect 24627 23069 24639 23103
rect 24581 23063 24639 23069
rect 24670 23060 24676 23112
rect 24728 23100 24734 23112
rect 24854 23100 24860 23112
rect 24728 23072 24773 23100
rect 24815 23072 24860 23100
rect 24728 23060 24734 23072
rect 24854 23060 24860 23072
rect 24912 23060 24918 23112
rect 25590 23100 25596 23112
rect 25551 23072 25596 23100
rect 25590 23060 25596 23072
rect 25648 23100 25654 23112
rect 26053 23103 26111 23109
rect 26053 23100 26065 23103
rect 25648 23072 26065 23100
rect 25648 23060 25654 23072
rect 26053 23069 26065 23072
rect 26099 23069 26111 23103
rect 26053 23063 26111 23069
rect 26881 23103 26939 23109
rect 26881 23069 26893 23103
rect 26927 23100 26939 23103
rect 26970 23100 26976 23112
rect 26927 23072 26976 23100
rect 26927 23069 26939 23072
rect 26881 23063 26939 23069
rect 26970 23060 26976 23072
rect 27028 23100 27034 23112
rect 27338 23100 27344 23112
rect 27028 23072 27344 23100
rect 27028 23060 27034 23072
rect 27338 23060 27344 23072
rect 27396 23060 27402 23112
rect 27908 23109 27936 23140
rect 27893 23103 27951 23109
rect 27893 23069 27905 23103
rect 27939 23100 27951 23103
rect 28350 23100 28356 23112
rect 27939 23072 28356 23100
rect 27939 23069 27951 23072
rect 27893 23063 27951 23069
rect 28350 23060 28356 23072
rect 28408 23060 28414 23112
rect 27706 23032 27712 23044
rect 23676 23004 27712 23032
rect 23569 22995 23627 23001
rect 27706 22992 27712 23004
rect 27764 22992 27770 23044
rect 12676 22936 14872 22964
rect 15565 22967 15623 22973
rect 12676 22924 12682 22936
rect 15565 22933 15577 22967
rect 15611 22964 15623 22967
rect 16393 22967 16451 22973
rect 16393 22964 16405 22967
rect 15611 22936 16405 22964
rect 15611 22933 15623 22936
rect 15565 22927 15623 22933
rect 16393 22933 16405 22936
rect 16439 22933 16451 22967
rect 17678 22964 17684 22976
rect 17639 22936 17684 22964
rect 16393 22927 16451 22933
rect 17678 22924 17684 22936
rect 17736 22924 17742 22976
rect 20993 22967 21051 22973
rect 20993 22933 21005 22967
rect 21039 22964 21051 22967
rect 21082 22964 21088 22976
rect 21039 22936 21088 22964
rect 21039 22933 21051 22936
rect 20993 22927 21051 22933
rect 21082 22924 21088 22936
rect 21140 22924 21146 22976
rect 21818 22964 21824 22976
rect 21779 22936 21824 22964
rect 21818 22924 21824 22936
rect 21876 22924 21882 22976
rect 22649 22967 22707 22973
rect 22649 22933 22661 22967
rect 22695 22964 22707 22967
rect 22738 22964 22744 22976
rect 22695 22936 22744 22964
rect 22695 22933 22707 22936
rect 22649 22927 22707 22933
rect 22738 22924 22744 22936
rect 22796 22924 22802 22976
rect 23474 22964 23480 22976
rect 23435 22936 23480 22964
rect 23474 22924 23480 22936
rect 23532 22924 23538 22976
rect 25130 22924 25136 22976
rect 25188 22964 25194 22976
rect 25409 22967 25467 22973
rect 25409 22964 25421 22967
rect 25188 22936 25421 22964
rect 25188 22924 25194 22936
rect 25409 22933 25421 22936
rect 25455 22933 25467 22967
rect 25409 22927 25467 22933
rect 1104 22874 28888 22896
rect 1104 22822 10214 22874
rect 10266 22822 10278 22874
rect 10330 22822 10342 22874
rect 10394 22822 10406 22874
rect 10458 22822 10470 22874
rect 10522 22822 19478 22874
rect 19530 22822 19542 22874
rect 19594 22822 19606 22874
rect 19658 22822 19670 22874
rect 19722 22822 19734 22874
rect 19786 22822 28888 22874
rect 1104 22800 28888 22822
rect 2682 22720 2688 22772
rect 2740 22760 2746 22772
rect 12618 22760 12624 22772
rect 2740 22732 12624 22760
rect 2740 22720 2746 22732
rect 12618 22720 12624 22732
rect 12676 22720 12682 22772
rect 12894 22760 12900 22772
rect 12855 22732 12900 22760
rect 12894 22720 12900 22732
rect 12952 22720 12958 22772
rect 18966 22760 18972 22772
rect 18927 22732 18972 22760
rect 18966 22720 18972 22732
rect 19024 22720 19030 22772
rect 20254 22760 20260 22772
rect 20215 22732 20260 22760
rect 20254 22720 20260 22732
rect 20312 22720 20318 22772
rect 23382 22760 23388 22772
rect 20364 22732 23388 22760
rect 4706 22652 4712 22704
rect 4764 22692 4770 22704
rect 12526 22692 12532 22704
rect 4764 22664 6914 22692
rect 12487 22664 12532 22692
rect 4764 22652 4770 22664
rect 6886 22488 6914 22664
rect 12526 22652 12532 22664
rect 12584 22652 12590 22704
rect 12710 22692 12716 22704
rect 12671 22664 12716 22692
rect 12710 22652 12716 22664
rect 12768 22652 12774 22704
rect 20364 22692 20392 22732
rect 23382 22720 23388 22732
rect 23440 22720 23446 22772
rect 23474 22720 23480 22772
rect 23532 22760 23538 22772
rect 24213 22763 24271 22769
rect 24213 22760 24225 22763
rect 23532 22732 24225 22760
rect 23532 22720 23538 22732
rect 24213 22729 24225 22732
rect 24259 22760 24271 22763
rect 24670 22760 24676 22772
rect 24259 22732 24676 22760
rect 24259 22729 24271 22732
rect 24213 22723 24271 22729
rect 24670 22720 24676 22732
rect 24728 22720 24734 22772
rect 25130 22720 25136 22772
rect 25188 22720 25194 22772
rect 13740 22664 20392 22692
rect 13740 22488 13768 22664
rect 21450 22652 21456 22704
rect 21508 22692 21514 22704
rect 21821 22695 21879 22701
rect 21821 22692 21833 22695
rect 21508 22664 21833 22692
rect 21508 22652 21514 22664
rect 21821 22661 21833 22664
rect 21867 22661 21879 22695
rect 21821 22655 21879 22661
rect 21910 22652 21916 22704
rect 21968 22692 21974 22704
rect 22021 22695 22079 22701
rect 22021 22692 22033 22695
rect 21968 22664 22033 22692
rect 21968 22652 21974 22664
rect 22021 22661 22033 22664
rect 22067 22661 22079 22695
rect 25148 22692 25176 22720
rect 22021 22655 22079 22661
rect 22848 22664 24992 22692
rect 25148 22664 27200 22692
rect 14458 22624 14464 22636
rect 14516 22633 14522 22636
rect 14428 22596 14464 22624
rect 14458 22584 14464 22596
rect 14516 22587 14528 22633
rect 14734 22624 14740 22636
rect 14695 22596 14740 22624
rect 14516 22584 14522 22587
rect 14734 22584 14740 22596
rect 14792 22584 14798 22636
rect 18874 22624 18880 22636
rect 18835 22596 18880 22624
rect 18874 22584 18880 22596
rect 18932 22584 18938 22636
rect 18966 22584 18972 22636
rect 19024 22624 19030 22636
rect 19061 22627 19119 22633
rect 19061 22624 19073 22627
rect 19024 22596 19073 22624
rect 19024 22584 19030 22596
rect 19061 22593 19073 22596
rect 19107 22593 19119 22627
rect 20070 22624 20076 22636
rect 20031 22596 20076 22624
rect 19061 22587 19119 22593
rect 20070 22584 20076 22596
rect 20128 22584 20134 22636
rect 22848 22633 22876 22664
rect 22833 22627 22891 22633
rect 22833 22624 22845 22627
rect 22066 22596 22845 22624
rect 20714 22516 20720 22568
rect 20772 22556 20778 22568
rect 22066 22556 22094 22596
rect 22833 22593 22845 22596
rect 22879 22593 22891 22627
rect 22833 22587 22891 22593
rect 22922 22584 22928 22636
rect 22980 22624 22986 22636
rect 24964 22633 24992 22664
rect 23089 22627 23147 22633
rect 23089 22624 23101 22627
rect 22980 22596 23101 22624
rect 22980 22584 22986 22596
rect 23089 22593 23101 22596
rect 23135 22593 23147 22627
rect 23089 22587 23147 22593
rect 24949 22627 25007 22633
rect 24949 22593 24961 22627
rect 24995 22593 25007 22627
rect 24949 22587 25007 22593
rect 25038 22584 25044 22636
rect 25096 22624 25102 22636
rect 27172 22633 27200 22664
rect 25205 22627 25263 22633
rect 25205 22624 25217 22627
rect 25096 22596 25217 22624
rect 25096 22584 25102 22596
rect 25205 22593 25217 22596
rect 25251 22593 25263 22627
rect 25205 22587 25263 22593
rect 27157 22627 27215 22633
rect 27157 22593 27169 22627
rect 27203 22593 27215 22627
rect 27706 22624 27712 22636
rect 27667 22596 27712 22624
rect 27157 22587 27215 22593
rect 27706 22584 27712 22596
rect 27764 22584 27770 22636
rect 20772 22528 22094 22556
rect 20772 22516 20778 22528
rect 6886 22460 13768 22488
rect 25958 22448 25964 22500
rect 26016 22488 26022 22500
rect 27801 22491 27859 22497
rect 27801 22488 27813 22491
rect 26016 22460 27813 22488
rect 26016 22448 26022 22460
rect 27801 22457 27813 22460
rect 27847 22457 27859 22491
rect 27801 22451 27859 22457
rect 13354 22420 13360 22432
rect 13315 22392 13360 22420
rect 13354 22380 13360 22392
rect 13412 22380 13418 22432
rect 22002 22420 22008 22432
rect 21963 22392 22008 22420
rect 22002 22380 22008 22392
rect 22060 22380 22066 22432
rect 22186 22420 22192 22432
rect 22147 22392 22192 22420
rect 22186 22380 22192 22392
rect 22244 22380 22250 22432
rect 26234 22380 26240 22432
rect 26292 22420 26298 22432
rect 26329 22423 26387 22429
rect 26329 22420 26341 22423
rect 26292 22392 26341 22420
rect 26292 22380 26298 22392
rect 26329 22389 26341 22392
rect 26375 22389 26387 22423
rect 26329 22383 26387 22389
rect 26510 22380 26516 22432
rect 26568 22420 26574 22432
rect 27065 22423 27123 22429
rect 27065 22420 27077 22423
rect 26568 22392 27077 22420
rect 26568 22380 26574 22392
rect 27065 22389 27077 22392
rect 27111 22389 27123 22423
rect 27065 22383 27123 22389
rect 1104 22330 28888 22352
rect 1104 22278 5582 22330
rect 5634 22278 5646 22330
rect 5698 22278 5710 22330
rect 5762 22278 5774 22330
rect 5826 22278 5838 22330
rect 5890 22278 14846 22330
rect 14898 22278 14910 22330
rect 14962 22278 14974 22330
rect 15026 22278 15038 22330
rect 15090 22278 15102 22330
rect 15154 22278 24110 22330
rect 24162 22278 24174 22330
rect 24226 22278 24238 22330
rect 24290 22278 24302 22330
rect 24354 22278 24366 22330
rect 24418 22278 28888 22330
rect 1104 22256 28888 22278
rect 14277 22219 14335 22225
rect 14277 22185 14289 22219
rect 14323 22216 14335 22219
rect 14458 22216 14464 22228
rect 14323 22188 14464 22216
rect 14323 22185 14335 22188
rect 14277 22179 14335 22185
rect 14458 22176 14464 22188
rect 14516 22176 14522 22228
rect 22922 22216 22928 22228
rect 22883 22188 22928 22216
rect 22922 22176 22928 22188
rect 22980 22176 22986 22228
rect 25038 22216 25044 22228
rect 24999 22188 25044 22216
rect 25038 22176 25044 22188
rect 25096 22176 25102 22228
rect 23845 22151 23903 22157
rect 23845 22117 23857 22151
rect 23891 22148 23903 22151
rect 25498 22148 25504 22160
rect 23891 22120 25504 22148
rect 23891 22117 23903 22120
rect 23845 22111 23903 22117
rect 25498 22108 25504 22120
rect 25556 22108 25562 22160
rect 26234 22148 26240 22160
rect 26068 22120 26240 22148
rect 12710 22040 12716 22092
rect 12768 22080 12774 22092
rect 17218 22080 17224 22092
rect 12768 22052 17224 22080
rect 12768 22040 12774 22052
rect 17218 22040 17224 22052
rect 17276 22040 17282 22092
rect 23658 22040 23664 22092
rect 23716 22080 23722 22092
rect 25409 22083 25467 22089
rect 23716 22052 25360 22080
rect 23716 22040 23722 22052
rect 25332 22024 25360 22052
rect 25409 22049 25421 22083
rect 25455 22080 25467 22083
rect 26068 22080 26096 22120
rect 26234 22108 26240 22120
rect 26292 22108 26298 22160
rect 26510 22080 26516 22092
rect 25455 22052 26096 22080
rect 26471 22052 26516 22080
rect 25455 22049 25467 22052
rect 25409 22043 25467 22049
rect 26510 22040 26516 22052
rect 26568 22040 26574 22092
rect 28169 22083 28227 22089
rect 28169 22049 28181 22083
rect 28215 22080 28227 22083
rect 28626 22080 28632 22092
rect 28215 22052 28632 22080
rect 28215 22049 28227 22052
rect 28169 22043 28227 22049
rect 28626 22040 28632 22052
rect 28684 22040 28690 22092
rect 1578 22012 1584 22024
rect 1539 21984 1584 22012
rect 1578 21972 1584 21984
rect 1636 21972 1642 22024
rect 14090 22012 14096 22024
rect 14051 21984 14096 22012
rect 14090 21972 14096 21984
rect 14148 21972 14154 22024
rect 19981 22015 20039 22021
rect 19981 21981 19993 22015
rect 20027 22012 20039 22015
rect 20162 22012 20168 22024
rect 20027 21984 20168 22012
rect 20027 21981 20039 21984
rect 19981 21975 20039 21981
rect 20162 21972 20168 21984
rect 20220 21972 20226 22024
rect 20898 21972 20904 22024
rect 20956 22012 20962 22024
rect 20993 22015 21051 22021
rect 20993 22012 21005 22015
rect 20956 21984 21005 22012
rect 20956 21972 20962 21984
rect 20993 21981 21005 21984
rect 21039 22012 21051 22015
rect 21634 22012 21640 22024
rect 21039 21984 21640 22012
rect 21039 21981 21051 21984
rect 20993 21975 21051 21981
rect 21634 21972 21640 21984
rect 21692 21972 21698 22024
rect 22738 22012 22744 22024
rect 22699 21984 22744 22012
rect 22738 21972 22744 21984
rect 22796 21972 22802 22024
rect 24578 22012 24584 22024
rect 24539 21984 24584 22012
rect 24578 21972 24584 21984
rect 24636 21972 24642 22024
rect 25222 22012 25228 22024
rect 25183 21984 25228 22012
rect 25222 21972 25228 21984
rect 25280 21972 25286 22024
rect 25314 21972 25320 22024
rect 25372 22012 25378 22024
rect 25501 22015 25559 22021
rect 25501 22012 25513 22015
rect 25372 21984 25513 22012
rect 25372 21972 25378 21984
rect 25501 21981 25513 21984
rect 25547 21981 25559 22015
rect 25501 21975 25559 21981
rect 26329 22015 26387 22021
rect 26329 21981 26341 22015
rect 26375 21981 26387 22015
rect 26329 21975 26387 21981
rect 21358 21944 21364 21956
rect 19812 21916 21364 21944
rect 19812 21885 19840 21916
rect 21358 21904 21364 21916
rect 21416 21904 21422 21956
rect 24489 21947 24547 21953
rect 24489 21913 24501 21947
rect 24535 21944 24547 21947
rect 26344 21944 26372 21975
rect 24535 21916 26372 21944
rect 24535 21913 24547 21916
rect 24489 21907 24547 21913
rect 19797 21879 19855 21885
rect 19797 21845 19809 21879
rect 19843 21845 19855 21879
rect 20806 21876 20812 21888
rect 20767 21848 20812 21876
rect 19797 21839 19855 21845
rect 20806 21836 20812 21848
rect 20864 21836 20870 21888
rect 1104 21786 28888 21808
rect 1104 21734 10214 21786
rect 10266 21734 10278 21786
rect 10330 21734 10342 21786
rect 10394 21734 10406 21786
rect 10458 21734 10470 21786
rect 10522 21734 19478 21786
rect 19530 21734 19542 21786
rect 19594 21734 19606 21786
rect 19658 21734 19670 21786
rect 19722 21734 19734 21786
rect 19786 21734 28888 21786
rect 1104 21712 28888 21734
rect 17218 21672 17224 21684
rect 17179 21644 17224 21672
rect 17218 21632 17224 21644
rect 17276 21632 17282 21684
rect 18049 21675 18107 21681
rect 18049 21641 18061 21675
rect 18095 21672 18107 21675
rect 18138 21672 18144 21684
rect 18095 21644 18144 21672
rect 18095 21641 18107 21644
rect 18049 21635 18107 21641
rect 18138 21632 18144 21644
rect 18196 21632 18202 21684
rect 18233 21675 18291 21681
rect 18233 21641 18245 21675
rect 18279 21672 18291 21675
rect 18414 21672 18420 21684
rect 18279 21644 18420 21672
rect 18279 21641 18291 21644
rect 18233 21635 18291 21641
rect 18414 21632 18420 21644
rect 18472 21632 18478 21684
rect 19334 21632 19340 21684
rect 19392 21672 19398 21684
rect 19705 21675 19763 21681
rect 19705 21672 19717 21675
rect 19392 21644 19717 21672
rect 19392 21632 19398 21644
rect 19705 21641 19717 21644
rect 19751 21641 19763 21675
rect 21358 21672 21364 21684
rect 19705 21635 19763 21641
rect 20364 21644 21364 21672
rect 15473 21607 15531 21613
rect 15473 21573 15485 21607
rect 15519 21604 15531 21607
rect 16758 21604 16764 21616
rect 15519 21576 16764 21604
rect 15519 21573 15531 21576
rect 15473 21567 15531 21573
rect 16758 21564 16764 21576
rect 16816 21564 16822 21616
rect 17678 21564 17684 21616
rect 17736 21604 17742 21616
rect 17865 21607 17923 21613
rect 17865 21604 17877 21607
rect 17736 21576 17877 21604
rect 17736 21564 17742 21576
rect 17865 21573 17877 21576
rect 17911 21573 17923 21607
rect 19058 21604 19064 21616
rect 19019 21576 19064 21604
rect 17865 21567 17923 21573
rect 19058 21564 19064 21576
rect 19116 21564 19122 21616
rect 2133 21539 2191 21545
rect 2133 21505 2145 21539
rect 2179 21536 2191 21539
rect 4706 21536 4712 21548
rect 2179 21508 4712 21536
rect 2179 21505 2191 21508
rect 2133 21499 2191 21505
rect 4706 21496 4712 21508
rect 4764 21496 4770 21548
rect 13354 21496 13360 21548
rect 13412 21536 13418 21548
rect 15289 21539 15347 21545
rect 15289 21536 15301 21539
rect 13412 21508 15301 21536
rect 13412 21496 13418 21508
rect 15289 21505 15301 21508
rect 15335 21536 15347 21539
rect 15378 21536 15384 21548
rect 15335 21508 15384 21536
rect 15335 21505 15347 21508
rect 15289 21499 15347 21505
rect 15378 21496 15384 21508
rect 15436 21496 15442 21548
rect 15562 21536 15568 21548
rect 15523 21508 15568 21536
rect 15562 21496 15568 21508
rect 15620 21496 15626 21548
rect 17310 21536 17316 21548
rect 17271 21508 17316 21536
rect 17310 21496 17316 21508
rect 17368 21496 17374 21548
rect 18046 21496 18052 21548
rect 18104 21536 18110 21548
rect 18141 21539 18199 21545
rect 18141 21536 18153 21539
rect 18104 21508 18153 21536
rect 18104 21496 18110 21508
rect 18141 21505 18153 21508
rect 18187 21505 18199 21539
rect 18141 21499 18199 21505
rect 2038 21332 2044 21344
rect 1999 21304 2044 21332
rect 2038 21292 2044 21304
rect 2096 21292 2102 21344
rect 14734 21292 14740 21344
rect 14792 21332 14798 21344
rect 15105 21335 15163 21341
rect 15105 21332 15117 21335
rect 14792 21304 15117 21332
rect 14792 21292 14798 21304
rect 15105 21301 15117 21304
rect 15151 21301 15163 21335
rect 15105 21295 15163 21301
rect 18417 21335 18475 21341
rect 18417 21301 18429 21335
rect 18463 21332 18475 21335
rect 18506 21332 18512 21344
rect 18463 21304 18512 21332
rect 18463 21301 18475 21304
rect 18417 21295 18475 21301
rect 18506 21292 18512 21304
rect 18564 21292 18570 21344
rect 18966 21332 18972 21344
rect 18927 21304 18972 21332
rect 18966 21292 18972 21304
rect 19024 21292 19030 21344
rect 19720 21332 19748 21635
rect 19889 21539 19947 21545
rect 19889 21505 19901 21539
rect 19935 21536 19947 21539
rect 20162 21536 20168 21548
rect 19935 21508 20168 21536
rect 19935 21505 19947 21508
rect 19889 21499 19947 21505
rect 20162 21496 20168 21508
rect 20220 21496 20226 21548
rect 20364 21545 20392 21644
rect 21358 21632 21364 21644
rect 21416 21672 21422 21684
rect 23658 21672 23664 21684
rect 21416 21644 23664 21672
rect 21416 21632 21422 21644
rect 23658 21632 23664 21644
rect 23716 21632 23722 21684
rect 20625 21607 20683 21613
rect 20625 21573 20637 21607
rect 20671 21604 20683 21607
rect 20806 21604 20812 21616
rect 20671 21576 20812 21604
rect 20671 21573 20683 21576
rect 20625 21567 20683 21573
rect 20806 21564 20812 21576
rect 20864 21564 20870 21616
rect 24765 21607 24823 21613
rect 24765 21573 24777 21607
rect 24811 21604 24823 21607
rect 25958 21604 25964 21616
rect 24811 21576 25964 21604
rect 24811 21573 24823 21576
rect 24765 21567 24823 21573
rect 25958 21564 25964 21576
rect 26016 21564 26022 21616
rect 20349 21539 20407 21545
rect 20349 21505 20361 21539
rect 20395 21505 20407 21539
rect 20349 21499 20407 21505
rect 20438 21496 20444 21548
rect 20496 21536 20502 21548
rect 21085 21539 21143 21545
rect 20496 21508 20541 21536
rect 20496 21496 20502 21508
rect 21085 21505 21097 21539
rect 21131 21505 21143 21539
rect 21085 21499 21143 21505
rect 21269 21539 21327 21545
rect 21269 21505 21281 21539
rect 21315 21505 21327 21539
rect 22002 21536 22008 21548
rect 21963 21508 22008 21536
rect 21269 21499 21327 21505
rect 21100 21468 21128 21499
rect 20640 21440 21128 21468
rect 20640 21409 20668 21440
rect 20625 21403 20683 21409
rect 20625 21369 20637 21403
rect 20671 21369 20683 21403
rect 21284 21400 21312 21499
rect 22002 21496 22008 21508
rect 22060 21496 22066 21548
rect 22186 21536 22192 21548
rect 22147 21508 22192 21536
rect 22186 21496 22192 21508
rect 22244 21496 22250 21548
rect 27706 21536 27712 21548
rect 27667 21508 27712 21536
rect 27706 21496 27712 21508
rect 27764 21496 27770 21548
rect 22278 21468 22284 21480
rect 22239 21440 22284 21468
rect 22278 21428 22284 21440
rect 22336 21428 22342 21480
rect 24121 21471 24179 21477
rect 24121 21437 24133 21471
rect 24167 21468 24179 21471
rect 24581 21471 24639 21477
rect 24581 21468 24593 21471
rect 24167 21440 24593 21468
rect 24167 21437 24179 21440
rect 24121 21431 24179 21437
rect 24581 21437 24593 21440
rect 24627 21437 24639 21471
rect 26142 21468 26148 21480
rect 26103 21440 26148 21468
rect 24581 21431 24639 21437
rect 26142 21428 26148 21440
rect 26200 21428 26206 21480
rect 24854 21400 24860 21412
rect 20625 21363 20683 21369
rect 20732 21372 24860 21400
rect 20732 21332 20760 21372
rect 24854 21360 24860 21372
rect 24912 21360 24918 21412
rect 19720 21304 20760 21332
rect 20806 21292 20812 21344
rect 20864 21332 20870 21344
rect 21085 21335 21143 21341
rect 21085 21332 21097 21335
rect 20864 21304 21097 21332
rect 20864 21292 20870 21304
rect 21085 21301 21097 21304
rect 21131 21301 21143 21335
rect 21085 21295 21143 21301
rect 21726 21292 21732 21344
rect 21784 21332 21790 21344
rect 21821 21335 21879 21341
rect 21821 21332 21833 21335
rect 21784 21304 21833 21332
rect 21784 21292 21790 21304
rect 21821 21301 21833 21304
rect 21867 21301 21879 21335
rect 21821 21295 21879 21301
rect 26510 21292 26516 21344
rect 26568 21332 26574 21344
rect 27617 21335 27675 21341
rect 27617 21332 27629 21335
rect 26568 21304 27629 21332
rect 26568 21292 26574 21304
rect 27617 21301 27629 21304
rect 27663 21301 27675 21335
rect 27617 21295 27675 21301
rect 1104 21242 28888 21264
rect 1104 21190 5582 21242
rect 5634 21190 5646 21242
rect 5698 21190 5710 21242
rect 5762 21190 5774 21242
rect 5826 21190 5838 21242
rect 5890 21190 14846 21242
rect 14898 21190 14910 21242
rect 14962 21190 14974 21242
rect 15026 21190 15038 21242
rect 15090 21190 15102 21242
rect 15154 21190 24110 21242
rect 24162 21190 24174 21242
rect 24226 21190 24238 21242
rect 24290 21190 24302 21242
rect 24354 21190 24366 21242
rect 24418 21190 28888 21242
rect 1104 21168 28888 21190
rect 14734 21088 14740 21140
rect 14792 21128 14798 21140
rect 15013 21131 15071 21137
rect 15013 21128 15025 21131
rect 14792 21100 15025 21128
rect 14792 21088 14798 21100
rect 15013 21097 15025 21100
rect 15059 21097 15071 21131
rect 15013 21091 15071 21097
rect 16758 21088 16764 21140
rect 16816 21128 16822 21140
rect 17037 21131 17095 21137
rect 17037 21128 17049 21131
rect 16816 21100 17049 21128
rect 16816 21088 16822 21100
rect 17037 21097 17049 21100
rect 17083 21097 17095 21131
rect 17037 21091 17095 21097
rect 19058 21088 19064 21140
rect 19116 21128 19122 21140
rect 19245 21131 19303 21137
rect 19245 21128 19257 21131
rect 19116 21100 19257 21128
rect 19116 21088 19122 21100
rect 19245 21097 19257 21100
rect 19291 21097 19303 21131
rect 19245 21091 19303 21097
rect 14090 21020 14096 21072
rect 14148 21060 14154 21072
rect 14829 21063 14887 21069
rect 14829 21060 14841 21063
rect 14148 21032 14841 21060
rect 14148 21020 14154 21032
rect 14829 21029 14841 21032
rect 14875 21029 14887 21063
rect 14829 21023 14887 21029
rect 1397 20995 1455 21001
rect 1397 20961 1409 20995
rect 1443 20992 1455 20995
rect 1578 20992 1584 21004
rect 1443 20964 1584 20992
rect 1443 20961 1455 20964
rect 1397 20955 1455 20961
rect 1578 20952 1584 20964
rect 1636 20952 1642 21004
rect 16776 20992 16804 21088
rect 15672 20964 16804 20992
rect 12437 20927 12495 20933
rect 12437 20893 12449 20927
rect 12483 20924 12495 20927
rect 13081 20927 13139 20933
rect 13081 20924 13093 20927
rect 12483 20896 13093 20924
rect 12483 20893 12495 20896
rect 12437 20887 12495 20893
rect 13081 20893 13093 20896
rect 13127 20893 13139 20927
rect 14274 20924 14280 20936
rect 14235 20896 14280 20924
rect 13081 20887 13139 20893
rect 14274 20884 14280 20896
rect 14332 20884 14338 20936
rect 15672 20933 15700 20964
rect 18506 20952 18512 21004
rect 18564 20992 18570 21004
rect 18564 20964 19748 20992
rect 18564 20952 18570 20964
rect 15657 20927 15715 20933
rect 15657 20893 15669 20927
rect 15703 20893 15715 20927
rect 15657 20887 15715 20893
rect 15841 20927 15899 20933
rect 15841 20893 15853 20927
rect 15887 20924 15899 20927
rect 16022 20924 16028 20936
rect 15887 20896 16028 20924
rect 15887 20893 15899 20896
rect 15841 20887 15899 20893
rect 16022 20884 16028 20896
rect 16080 20884 16086 20936
rect 16850 20884 16856 20936
rect 16908 20924 16914 20936
rect 16945 20927 17003 20933
rect 16945 20924 16957 20927
rect 16908 20896 16957 20924
rect 16908 20884 16914 20896
rect 16945 20893 16957 20896
rect 16991 20893 17003 20927
rect 16945 20887 17003 20893
rect 17770 20884 17776 20936
rect 17828 20924 17834 20936
rect 17921 20927 17979 20933
rect 17921 20924 17933 20927
rect 17828 20896 17933 20924
rect 17828 20884 17834 20896
rect 17921 20893 17933 20896
rect 17967 20893 17979 20927
rect 18046 20924 18052 20936
rect 18007 20896 18052 20924
rect 17921 20887 17979 20893
rect 18046 20884 18052 20896
rect 18104 20884 18110 20936
rect 18138 20884 18144 20936
rect 18196 20924 18202 20936
rect 18196 20896 18241 20924
rect 18196 20884 18202 20896
rect 18782 20884 18788 20936
rect 18840 20924 18846 20936
rect 19720 20933 19748 20964
rect 23198 20952 23204 21004
rect 23256 20992 23262 21004
rect 25225 20995 25283 21001
rect 25225 20992 25237 20995
rect 23256 20964 25237 20992
rect 23256 20952 23262 20964
rect 25225 20961 25237 20964
rect 25271 20961 25283 20995
rect 25225 20955 25283 20961
rect 25314 20952 25320 21004
rect 25372 20992 25378 21004
rect 25372 20964 25417 20992
rect 25372 20952 25378 20964
rect 25498 20952 25504 21004
rect 25556 20992 25562 21004
rect 26329 20995 26387 21001
rect 26329 20992 26341 20995
rect 25556 20964 26341 20992
rect 25556 20952 25562 20964
rect 26329 20961 26341 20964
rect 26375 20961 26387 20995
rect 26510 20992 26516 21004
rect 26471 20964 26516 20992
rect 26329 20955 26387 20961
rect 26510 20952 26516 20964
rect 26568 20952 26574 21004
rect 28166 20992 28172 21004
rect 28127 20964 28172 20992
rect 28166 20952 28172 20964
rect 28224 20952 28230 21004
rect 19429 20927 19487 20933
rect 19429 20924 19441 20927
rect 18840 20896 19441 20924
rect 18840 20884 18846 20896
rect 19429 20893 19441 20896
rect 19475 20893 19487 20927
rect 19429 20887 19487 20893
rect 19521 20927 19579 20933
rect 19521 20893 19533 20927
rect 19567 20893 19579 20927
rect 19521 20887 19579 20893
rect 19705 20927 19763 20933
rect 19705 20893 19717 20927
rect 19751 20893 19763 20927
rect 19705 20887 19763 20893
rect 19797 20927 19855 20933
rect 19797 20893 19809 20927
rect 19843 20924 19855 20927
rect 20438 20924 20444 20936
rect 19843 20896 20444 20924
rect 19843 20893 19855 20896
rect 19797 20887 19855 20893
rect 1581 20859 1639 20865
rect 1581 20825 1593 20859
rect 1627 20856 1639 20859
rect 2038 20856 2044 20868
rect 1627 20828 2044 20856
rect 1627 20825 1639 20828
rect 1581 20819 1639 20825
rect 2038 20816 2044 20828
rect 2096 20816 2102 20868
rect 3237 20859 3295 20865
rect 3237 20825 3249 20859
rect 3283 20856 3295 20859
rect 3694 20856 3700 20868
rect 3283 20828 3700 20856
rect 3283 20825 3295 20828
rect 3237 20819 3295 20825
rect 3694 20816 3700 20828
rect 3752 20816 3758 20868
rect 12066 20856 12072 20868
rect 12027 20828 12072 20856
rect 12066 20816 12072 20828
rect 12124 20816 12130 20868
rect 12253 20859 12311 20865
rect 12253 20825 12265 20859
rect 12299 20856 12311 20859
rect 12710 20856 12716 20868
rect 12299 20828 12716 20856
rect 12299 20825 12311 20828
rect 12253 20819 12311 20825
rect 12710 20816 12716 20828
rect 12768 20816 12774 20868
rect 15197 20859 15255 20865
rect 15197 20825 15209 20859
rect 15243 20856 15255 20859
rect 15470 20856 15476 20868
rect 15243 20828 15476 20856
rect 15243 20825 15255 20828
rect 15197 20819 15255 20825
rect 15470 20816 15476 20828
rect 15528 20856 15534 20868
rect 15746 20856 15752 20868
rect 15528 20828 15752 20856
rect 15528 20816 15534 20828
rect 15746 20816 15752 20828
rect 15804 20816 15810 20868
rect 18325 20859 18383 20865
rect 18325 20825 18337 20859
rect 18371 20856 18383 20859
rect 18690 20856 18696 20868
rect 18371 20828 18696 20856
rect 18371 20825 18383 20828
rect 18325 20819 18383 20825
rect 18690 20816 18696 20828
rect 18748 20856 18754 20868
rect 19536 20856 19564 20887
rect 20438 20884 20444 20896
rect 20496 20884 20502 20936
rect 20993 20927 21051 20933
rect 20993 20893 21005 20927
rect 21039 20924 21051 20927
rect 21082 20924 21088 20936
rect 21039 20896 21088 20924
rect 21039 20893 21051 20896
rect 20993 20887 21051 20893
rect 21082 20884 21088 20896
rect 21140 20884 21146 20936
rect 21450 20924 21456 20936
rect 21411 20896 21456 20924
rect 21450 20884 21456 20896
rect 21508 20884 21514 20936
rect 21726 20933 21732 20936
rect 21720 20924 21732 20933
rect 21687 20896 21732 20924
rect 21720 20887 21732 20896
rect 21726 20884 21732 20887
rect 21784 20884 21790 20936
rect 23293 20927 23351 20933
rect 23293 20893 23305 20927
rect 23339 20924 23351 20927
rect 23566 20924 23572 20936
rect 23339 20896 23572 20924
rect 23339 20893 23351 20896
rect 23293 20887 23351 20893
rect 23566 20884 23572 20896
rect 23624 20884 23630 20936
rect 18748 20828 19564 20856
rect 18748 20816 18754 20828
rect 12618 20748 12624 20800
rect 12676 20788 12682 20800
rect 12897 20791 12955 20797
rect 12897 20788 12909 20791
rect 12676 20760 12909 20788
rect 12676 20748 12682 20760
rect 12897 20757 12909 20760
rect 12943 20757 12955 20791
rect 14090 20788 14096 20800
rect 14051 20760 14096 20788
rect 12897 20751 12955 20757
rect 14090 20748 14096 20760
rect 14148 20748 14154 20800
rect 14734 20748 14740 20800
rect 14792 20788 14798 20800
rect 14987 20791 15045 20797
rect 14987 20788 14999 20791
rect 14792 20760 14999 20788
rect 14792 20748 14798 20760
rect 14987 20757 14999 20760
rect 15033 20757 15045 20791
rect 14987 20751 15045 20757
rect 15286 20748 15292 20800
rect 15344 20788 15350 20800
rect 15657 20791 15715 20797
rect 15657 20788 15669 20791
rect 15344 20760 15669 20788
rect 15344 20748 15350 20760
rect 15657 20757 15669 20760
rect 15703 20757 15715 20791
rect 15657 20751 15715 20757
rect 17310 20748 17316 20800
rect 17368 20788 17374 20800
rect 20162 20788 20168 20800
rect 17368 20760 20168 20788
rect 17368 20748 17374 20760
rect 20162 20748 20168 20760
rect 20220 20748 20226 20800
rect 20809 20791 20867 20797
rect 20809 20757 20821 20791
rect 20855 20788 20867 20791
rect 22462 20788 22468 20800
rect 20855 20760 22468 20788
rect 20855 20757 20867 20760
rect 20809 20751 20867 20757
rect 22462 20748 22468 20760
rect 22520 20748 22526 20800
rect 22830 20788 22836 20800
rect 22791 20760 22836 20788
rect 22830 20748 22836 20760
rect 22888 20748 22894 20800
rect 23477 20791 23535 20797
rect 23477 20757 23489 20791
rect 23523 20788 23535 20791
rect 23750 20788 23756 20800
rect 23523 20760 23756 20788
rect 23523 20757 23535 20760
rect 23477 20751 23535 20757
rect 23750 20748 23756 20760
rect 23808 20748 23814 20800
rect 24486 20748 24492 20800
rect 24544 20788 24550 20800
rect 24765 20791 24823 20797
rect 24765 20788 24777 20791
rect 24544 20760 24777 20788
rect 24544 20748 24550 20760
rect 24765 20757 24777 20760
rect 24811 20757 24823 20791
rect 25130 20788 25136 20800
rect 25091 20760 25136 20788
rect 24765 20751 24823 20757
rect 25130 20748 25136 20760
rect 25188 20748 25194 20800
rect 1104 20698 28888 20720
rect 1104 20646 10214 20698
rect 10266 20646 10278 20698
rect 10330 20646 10342 20698
rect 10394 20646 10406 20698
rect 10458 20646 10470 20698
rect 10522 20646 19478 20698
rect 19530 20646 19542 20698
rect 19594 20646 19606 20698
rect 19658 20646 19670 20698
rect 19722 20646 19734 20698
rect 19786 20646 28888 20698
rect 1104 20624 28888 20646
rect 18325 20587 18383 20593
rect 18325 20553 18337 20587
rect 18371 20584 18383 20587
rect 18414 20584 18420 20596
rect 18371 20556 18420 20584
rect 18371 20553 18383 20556
rect 18325 20547 18383 20553
rect 18414 20544 18420 20556
rect 18472 20544 18478 20596
rect 18690 20584 18696 20596
rect 18651 20556 18696 20584
rect 18690 20544 18696 20556
rect 18748 20544 18754 20596
rect 21082 20584 21088 20596
rect 21043 20556 21088 20584
rect 21082 20544 21088 20556
rect 21140 20544 21146 20596
rect 22557 20587 22615 20593
rect 22557 20553 22569 20587
rect 22603 20584 22615 20587
rect 22830 20584 22836 20596
rect 22603 20556 22836 20584
rect 22603 20553 22615 20556
rect 22557 20547 22615 20553
rect 22830 20544 22836 20556
rect 22888 20544 22894 20596
rect 25869 20587 25927 20593
rect 25869 20553 25881 20587
rect 25915 20584 25927 20587
rect 26142 20584 26148 20596
rect 25915 20556 26148 20584
rect 25915 20553 25927 20556
rect 25869 20547 25927 20553
rect 26142 20544 26148 20556
rect 26200 20544 26206 20596
rect 12158 20516 12164 20528
rect 11992 20488 12164 20516
rect 2314 20380 2320 20392
rect 2275 20352 2320 20380
rect 2314 20340 2320 20352
rect 2372 20340 2378 20392
rect 2501 20383 2559 20389
rect 2501 20349 2513 20383
rect 2547 20380 2559 20383
rect 2866 20380 2872 20392
rect 2547 20352 2872 20380
rect 2547 20349 2559 20352
rect 2501 20343 2559 20349
rect 2866 20340 2872 20352
rect 2924 20340 2930 20392
rect 2958 20340 2964 20392
rect 3016 20380 3022 20392
rect 3016 20352 3061 20380
rect 3016 20340 3022 20352
rect 11882 20340 11888 20392
rect 11940 20380 11946 20392
rect 11992 20389 12020 20488
rect 12158 20476 12164 20488
rect 12216 20516 12222 20528
rect 14090 20525 14096 20528
rect 14084 20516 14096 20525
rect 12216 20488 13860 20516
rect 14051 20488 14096 20516
rect 12216 20476 12222 20488
rect 12244 20451 12302 20457
rect 12244 20417 12256 20451
rect 12290 20448 12302 20451
rect 12618 20448 12624 20460
rect 12290 20420 12624 20448
rect 12290 20417 12302 20420
rect 12244 20411 12302 20417
rect 12618 20408 12624 20420
rect 12676 20408 12682 20460
rect 13832 20457 13860 20488
rect 14084 20479 14096 20488
rect 14090 20476 14096 20479
rect 14148 20476 14154 20528
rect 15657 20519 15715 20525
rect 15657 20516 15669 20519
rect 15212 20488 15669 20516
rect 13817 20451 13875 20457
rect 13817 20417 13829 20451
rect 13863 20417 13875 20451
rect 13817 20411 13875 20417
rect 11977 20383 12035 20389
rect 11977 20380 11989 20383
rect 11940 20352 11989 20380
rect 11940 20340 11946 20352
rect 11977 20349 11989 20352
rect 12023 20349 12035 20383
rect 11977 20343 12035 20349
rect 15212 20256 15240 20488
rect 15657 20485 15669 20488
rect 15703 20485 15715 20519
rect 15657 20479 15715 20485
rect 15887 20485 15945 20491
rect 15887 20482 15899 20485
rect 15562 20408 15568 20460
rect 15620 20448 15626 20460
rect 15872 20451 15899 20482
rect 15933 20460 15945 20485
rect 16850 20476 16856 20528
rect 16908 20516 16914 20528
rect 17221 20519 17279 20525
rect 17221 20516 17233 20519
rect 16908 20488 17233 20516
rect 16908 20476 16914 20488
rect 17221 20485 17233 20488
rect 17267 20485 17279 20519
rect 17221 20479 17279 20485
rect 19972 20519 20030 20525
rect 19972 20485 19984 20519
rect 20018 20516 20030 20519
rect 20806 20516 20812 20528
rect 20018 20488 20812 20516
rect 20018 20485 20030 20488
rect 19972 20479 20030 20485
rect 20806 20476 20812 20488
rect 20864 20476 20870 20528
rect 20990 20476 20996 20528
rect 21048 20516 21054 20528
rect 21450 20516 21456 20528
rect 21048 20488 21456 20516
rect 21048 20476 21054 20488
rect 21450 20476 21456 20488
rect 21508 20516 21514 20528
rect 23750 20525 23756 20528
rect 23744 20516 23756 20525
rect 21508 20488 23520 20516
rect 23711 20488 23756 20516
rect 21508 20476 21514 20488
rect 23492 20460 23520 20488
rect 23744 20479 23756 20488
rect 23750 20476 23756 20479
rect 23808 20476 23814 20528
rect 15933 20451 15936 20460
rect 15872 20448 15936 20451
rect 15620 20420 15936 20448
rect 15620 20408 15626 20420
rect 15930 20408 15936 20420
rect 15988 20408 15994 20460
rect 18506 20448 18512 20460
rect 18467 20420 18512 20448
rect 18506 20408 18512 20420
rect 18564 20408 18570 20460
rect 18782 20408 18788 20460
rect 18840 20448 18846 20460
rect 22649 20451 22707 20457
rect 18840 20420 18885 20448
rect 18840 20408 18846 20420
rect 22649 20417 22661 20451
rect 22695 20417 22707 20451
rect 23474 20448 23480 20460
rect 23387 20420 23480 20448
rect 22649 20411 22707 20417
rect 19705 20383 19763 20389
rect 19705 20349 19717 20383
rect 19751 20349 19763 20383
rect 22462 20380 22468 20392
rect 22423 20352 22468 20380
rect 19705 20343 19763 20349
rect 13357 20247 13415 20253
rect 13357 20213 13369 20247
rect 13403 20244 13415 20247
rect 14090 20244 14096 20256
rect 13403 20216 14096 20244
rect 13403 20213 13415 20216
rect 13357 20207 13415 20213
rect 14090 20204 14096 20216
rect 14148 20204 14154 20256
rect 15194 20244 15200 20256
rect 15155 20216 15200 20244
rect 15194 20204 15200 20216
rect 15252 20204 15258 20256
rect 15378 20204 15384 20256
rect 15436 20244 15442 20256
rect 15746 20244 15752 20256
rect 15436 20216 15752 20244
rect 15436 20204 15442 20216
rect 15746 20204 15752 20216
rect 15804 20244 15810 20256
rect 15841 20247 15899 20253
rect 15841 20244 15853 20247
rect 15804 20216 15853 20244
rect 15804 20204 15810 20216
rect 15841 20213 15853 20216
rect 15887 20213 15899 20247
rect 16022 20244 16028 20256
rect 15983 20216 16028 20244
rect 15841 20207 15899 20213
rect 16022 20204 16028 20216
rect 16080 20204 16086 20256
rect 17129 20247 17187 20253
rect 17129 20213 17141 20247
rect 17175 20244 17187 20247
rect 17678 20244 17684 20256
rect 17175 20216 17684 20244
rect 17175 20213 17187 20216
rect 17129 20207 17187 20213
rect 17678 20204 17684 20216
rect 17736 20204 17742 20256
rect 19720 20244 19748 20343
rect 22462 20340 22468 20352
rect 22520 20340 22526 20392
rect 22664 20312 22692 20411
rect 23474 20408 23480 20420
rect 23532 20408 23538 20460
rect 25777 20451 25835 20457
rect 25777 20448 25789 20451
rect 24872 20420 25789 20448
rect 22664 20284 23520 20312
rect 20714 20244 20720 20256
rect 19720 20216 20720 20244
rect 20714 20204 20720 20216
rect 20772 20244 20778 20256
rect 20990 20244 20996 20256
rect 20772 20216 20996 20244
rect 20772 20204 20778 20216
rect 20990 20204 20996 20216
rect 21048 20204 21054 20256
rect 23017 20247 23075 20253
rect 23017 20213 23029 20247
rect 23063 20244 23075 20247
rect 23382 20244 23388 20256
rect 23063 20216 23388 20244
rect 23063 20213 23075 20216
rect 23017 20207 23075 20213
rect 23382 20204 23388 20216
rect 23440 20204 23446 20256
rect 23492 20244 23520 20284
rect 24872 20253 24900 20420
rect 25777 20417 25789 20420
rect 25823 20417 25835 20451
rect 27338 20448 27344 20460
rect 27299 20420 27344 20448
rect 25777 20411 25835 20417
rect 27338 20408 27344 20420
rect 27396 20408 27402 20460
rect 28074 20448 28080 20460
rect 28035 20420 28080 20448
rect 28074 20408 28080 20420
rect 28132 20408 28138 20460
rect 24946 20340 24952 20392
rect 25004 20380 25010 20392
rect 25682 20380 25688 20392
rect 25004 20352 25688 20380
rect 25004 20340 25010 20352
rect 25682 20340 25688 20352
rect 25740 20380 25746 20392
rect 25961 20383 26019 20389
rect 25961 20380 25973 20383
rect 25740 20352 25973 20380
rect 25740 20340 25746 20352
rect 25961 20349 25973 20352
rect 26007 20349 26019 20383
rect 25961 20343 26019 20349
rect 24857 20247 24915 20253
rect 24857 20244 24869 20247
rect 23492 20216 24869 20244
rect 24857 20213 24869 20216
rect 24903 20213 24915 20247
rect 25406 20244 25412 20256
rect 25367 20216 25412 20244
rect 24857 20207 24915 20213
rect 25406 20204 25412 20216
rect 25464 20204 25470 20256
rect 26510 20204 26516 20256
rect 26568 20244 26574 20256
rect 27249 20247 27307 20253
rect 27249 20244 27261 20247
rect 26568 20216 27261 20244
rect 26568 20204 26574 20216
rect 27249 20213 27261 20216
rect 27295 20213 27307 20247
rect 27249 20207 27307 20213
rect 1104 20154 28888 20176
rect 1104 20102 5582 20154
rect 5634 20102 5646 20154
rect 5698 20102 5710 20154
rect 5762 20102 5774 20154
rect 5826 20102 5838 20154
rect 5890 20102 14846 20154
rect 14898 20102 14910 20154
rect 14962 20102 14974 20154
rect 15026 20102 15038 20154
rect 15090 20102 15102 20154
rect 15154 20102 24110 20154
rect 24162 20102 24174 20154
rect 24226 20102 24238 20154
rect 24290 20102 24302 20154
rect 24354 20102 24366 20154
rect 24418 20102 28888 20154
rect 1104 20080 28888 20102
rect 2314 20040 2320 20052
rect 2275 20012 2320 20040
rect 2314 20000 2320 20012
rect 2372 20000 2378 20052
rect 2866 20040 2872 20052
rect 2827 20012 2872 20040
rect 2866 20000 2872 20012
rect 2924 20000 2930 20052
rect 12066 20000 12072 20052
rect 12124 20040 12130 20052
rect 12253 20043 12311 20049
rect 12253 20040 12265 20043
rect 12124 20012 12265 20040
rect 12124 20000 12130 20012
rect 12253 20009 12265 20012
rect 12299 20009 12311 20043
rect 12253 20003 12311 20009
rect 14274 20000 14280 20052
rect 14332 20040 14338 20052
rect 14829 20043 14887 20049
rect 14829 20040 14841 20043
rect 14332 20012 14841 20040
rect 14332 20000 14338 20012
rect 14829 20009 14841 20012
rect 14875 20009 14887 20043
rect 14829 20003 14887 20009
rect 15013 20043 15071 20049
rect 15013 20009 15025 20043
rect 15059 20040 15071 20043
rect 15286 20040 15292 20052
rect 15059 20012 15292 20040
rect 15059 20009 15071 20012
rect 15013 20003 15071 20009
rect 15286 20000 15292 20012
rect 15344 20000 15350 20052
rect 18325 20043 18383 20049
rect 18325 20040 18337 20043
rect 15856 20012 18337 20040
rect 15856 19916 15884 20012
rect 18325 20009 18337 20012
rect 18371 20009 18383 20043
rect 21358 20040 21364 20052
rect 21319 20012 21364 20040
rect 18325 20003 18383 20009
rect 21358 20000 21364 20012
rect 21416 20000 21422 20052
rect 22278 20040 22284 20052
rect 22239 20012 22284 20040
rect 22278 20000 22284 20012
rect 22336 20000 22342 20052
rect 23566 20040 23572 20052
rect 23527 20012 23572 20040
rect 23566 20000 23572 20012
rect 23624 20000 23630 20052
rect 25130 20000 25136 20052
rect 25188 20040 25194 20052
rect 25869 20043 25927 20049
rect 25869 20040 25881 20043
rect 25188 20012 25881 20040
rect 25188 20000 25194 20012
rect 25869 20009 25881 20012
rect 25915 20009 25927 20043
rect 25869 20003 25927 20009
rect 16666 19932 16672 19984
rect 16724 19972 16730 19984
rect 16761 19975 16819 19981
rect 16761 19972 16773 19975
rect 16724 19944 16773 19972
rect 16724 19932 16730 19944
rect 16761 19941 16773 19944
rect 16807 19941 16819 19975
rect 16761 19935 16819 19941
rect 18966 19932 18972 19984
rect 19024 19972 19030 19984
rect 22186 19972 22192 19984
rect 19024 19944 22192 19972
rect 19024 19932 19030 19944
rect 22186 19932 22192 19944
rect 22244 19932 22250 19984
rect 12802 19904 12808 19916
rect 12763 19876 12808 19904
rect 12802 19864 12808 19876
rect 12860 19864 12866 19916
rect 15470 19904 15476 19916
rect 15304 19876 15476 19904
rect 1394 19796 1400 19848
rect 1452 19836 1458 19848
rect 1489 19839 1547 19845
rect 1489 19836 1501 19839
rect 1452 19808 1501 19836
rect 1452 19796 1458 19808
rect 1489 19805 1501 19808
rect 1535 19805 1547 19839
rect 1489 19799 1547 19805
rect 2961 19839 3019 19845
rect 2961 19805 2973 19839
rect 3007 19836 3019 19839
rect 4154 19836 4160 19848
rect 3007 19808 4160 19836
rect 3007 19805 3019 19808
rect 2961 19799 3019 19805
rect 2976 19712 3004 19799
rect 4154 19796 4160 19808
rect 4212 19796 4218 19848
rect 14182 19836 14188 19848
rect 14143 19808 14188 19836
rect 14182 19796 14188 19808
rect 14240 19796 14246 19848
rect 14369 19839 14427 19845
rect 14369 19805 14381 19839
rect 14415 19836 14427 19839
rect 14734 19836 14740 19848
rect 14415 19808 14740 19836
rect 14415 19805 14427 19808
rect 14369 19799 14427 19805
rect 14734 19796 14740 19808
rect 14792 19836 14798 19848
rect 14792 19808 15148 19836
rect 14792 19796 14798 19808
rect 12621 19771 12679 19777
rect 12621 19737 12633 19771
rect 12667 19768 12679 19771
rect 14090 19768 14096 19780
rect 12667 19740 14096 19768
rect 12667 19737 12679 19740
rect 12621 19731 12679 19737
rect 14090 19728 14096 19740
rect 14148 19728 14154 19780
rect 14277 19771 14335 19777
rect 14277 19737 14289 19771
rect 14323 19768 14335 19771
rect 14981 19771 15039 19777
rect 14981 19768 14993 19771
rect 14323 19740 14993 19768
rect 14323 19737 14335 19740
rect 14277 19731 14335 19737
rect 14981 19737 14993 19740
rect 15027 19737 15039 19771
rect 14981 19731 15039 19737
rect 2958 19660 2964 19712
rect 3016 19660 3022 19712
rect 12710 19660 12716 19712
rect 12768 19700 12774 19712
rect 15120 19700 15148 19808
rect 15197 19771 15255 19777
rect 15197 19737 15209 19771
rect 15243 19768 15255 19771
rect 15304 19768 15332 19876
rect 15470 19864 15476 19876
rect 15528 19904 15534 19916
rect 15838 19904 15844 19916
rect 15528 19876 15844 19904
rect 15528 19864 15534 19876
rect 15838 19864 15844 19876
rect 15896 19864 15902 19916
rect 20625 19907 20683 19913
rect 17696 19876 18460 19904
rect 15657 19839 15715 19845
rect 15657 19805 15669 19839
rect 15703 19805 15715 19839
rect 15657 19799 15715 19805
rect 15243 19740 15332 19768
rect 15243 19737 15255 19740
rect 15197 19731 15255 19737
rect 15378 19728 15384 19780
rect 15436 19768 15442 19780
rect 15672 19768 15700 19799
rect 15746 19796 15752 19848
rect 15804 19836 15810 19848
rect 15930 19836 15936 19848
rect 15804 19808 15849 19836
rect 15891 19808 15936 19836
rect 15804 19796 15810 19808
rect 15930 19796 15936 19808
rect 15988 19796 15994 19848
rect 16945 19839 17003 19845
rect 16945 19805 16957 19839
rect 16991 19836 17003 19839
rect 17402 19836 17408 19848
rect 16991 19808 17408 19836
rect 16991 19805 17003 19808
rect 16945 19799 17003 19805
rect 17402 19796 17408 19808
rect 17460 19836 17466 19848
rect 17569 19839 17627 19845
rect 17569 19836 17581 19839
rect 17460 19808 17581 19836
rect 17460 19796 17466 19808
rect 17569 19805 17581 19808
rect 17615 19836 17627 19839
rect 17696 19836 17724 19876
rect 17615 19808 17724 19836
rect 17773 19839 17831 19845
rect 17615 19805 17627 19808
rect 17569 19799 17627 19805
rect 17773 19805 17785 19839
rect 17819 19836 17831 19839
rect 18322 19836 18328 19848
rect 17819 19808 18328 19836
rect 17819 19805 17831 19808
rect 17773 19799 17831 19805
rect 18322 19796 18328 19808
rect 18380 19796 18386 19848
rect 18432 19845 18460 19876
rect 20625 19873 20637 19907
rect 20671 19904 20683 19907
rect 22465 19907 22523 19913
rect 20671 19876 22048 19904
rect 20671 19873 20683 19876
rect 20625 19867 20683 19873
rect 18417 19839 18475 19845
rect 18417 19805 18429 19839
rect 18463 19805 18475 19839
rect 18417 19799 18475 19805
rect 20257 19839 20315 19845
rect 20257 19805 20269 19839
rect 20303 19836 20315 19839
rect 20898 19836 20904 19848
rect 20303 19808 20904 19836
rect 20303 19805 20315 19808
rect 20257 19799 20315 19805
rect 20898 19796 20904 19808
rect 20956 19796 20962 19848
rect 21082 19796 21088 19848
rect 21140 19836 21146 19848
rect 22020 19845 22048 19876
rect 22465 19873 22477 19907
rect 22511 19904 22523 19907
rect 22830 19904 22836 19916
rect 22511 19876 22836 19904
rect 22511 19873 22523 19876
rect 22465 19867 22523 19873
rect 22830 19864 22836 19876
rect 22888 19864 22894 19916
rect 23474 19864 23480 19916
rect 23532 19904 23538 19916
rect 24489 19907 24547 19913
rect 24489 19904 24501 19907
rect 23532 19876 24501 19904
rect 23532 19864 23538 19876
rect 24489 19873 24501 19876
rect 24535 19873 24547 19907
rect 26510 19904 26516 19916
rect 26471 19876 26516 19904
rect 24489 19867 24547 19873
rect 26510 19864 26516 19876
rect 26568 19864 26574 19916
rect 28166 19904 28172 19916
rect 28127 19876 28172 19904
rect 28166 19864 28172 19876
rect 28224 19864 28230 19916
rect 21269 19839 21327 19845
rect 21269 19836 21281 19839
rect 21140 19808 21281 19836
rect 21140 19796 21146 19808
rect 21269 19805 21281 19808
rect 21315 19805 21327 19839
rect 21269 19799 21327 19805
rect 22005 19839 22063 19845
rect 22005 19805 22017 19839
rect 22051 19836 22063 19839
rect 22738 19836 22744 19848
rect 22051 19808 22744 19836
rect 22051 19805 22063 19808
rect 22005 19799 22063 19805
rect 22738 19796 22744 19808
rect 22796 19796 22802 19848
rect 23201 19839 23259 19845
rect 23201 19805 23213 19839
rect 23247 19805 23259 19839
rect 23382 19836 23388 19848
rect 23343 19808 23388 19836
rect 23201 19799 23259 19805
rect 15436 19740 15792 19768
rect 15436 19728 15442 19740
rect 15657 19703 15715 19709
rect 15657 19700 15669 19703
rect 12768 19672 12813 19700
rect 15120 19672 15669 19700
rect 12768 19660 12774 19672
rect 15657 19669 15669 19672
rect 15703 19669 15715 19703
rect 15764 19700 15792 19740
rect 17310 19728 17316 19780
rect 17368 19768 17374 19780
rect 17487 19771 17545 19777
rect 17487 19768 17499 19771
rect 17368 19740 17499 19768
rect 17368 19728 17374 19740
rect 17487 19737 17499 19740
rect 17533 19737 17545 19771
rect 17487 19731 17545 19737
rect 17678 19728 17684 19780
rect 17736 19768 17742 19780
rect 20441 19771 20499 19777
rect 20441 19768 20453 19771
rect 17736 19740 20453 19768
rect 17736 19728 17742 19740
rect 20441 19737 20453 19740
rect 20487 19737 20499 19771
rect 20441 19731 20499 19737
rect 22097 19771 22155 19777
rect 22097 19737 22109 19771
rect 22143 19768 22155 19771
rect 22186 19768 22192 19780
rect 22143 19740 22192 19768
rect 22143 19737 22155 19740
rect 22097 19731 22155 19737
rect 22186 19728 22192 19740
rect 22244 19768 22250 19780
rect 22830 19768 22836 19780
rect 22244 19740 22836 19768
rect 22244 19728 22250 19740
rect 22830 19728 22836 19740
rect 22888 19728 22894 19780
rect 23216 19768 23244 19799
rect 23382 19796 23388 19808
rect 23440 19796 23446 19848
rect 26326 19836 26332 19848
rect 26287 19808 26332 19836
rect 26326 19796 26332 19808
rect 26384 19796 26390 19848
rect 24026 19768 24032 19780
rect 23216 19740 24032 19768
rect 24026 19728 24032 19740
rect 24084 19728 24090 19780
rect 24756 19771 24814 19777
rect 24756 19737 24768 19771
rect 24802 19768 24814 19771
rect 25130 19768 25136 19780
rect 24802 19740 25136 19768
rect 24802 19737 24814 19740
rect 24756 19731 24814 19737
rect 25130 19728 25136 19740
rect 25188 19728 25194 19780
rect 17696 19700 17724 19728
rect 15764 19672 17724 19700
rect 15657 19663 15715 19669
rect 22462 19660 22468 19712
rect 22520 19700 22526 19712
rect 23658 19700 23664 19712
rect 22520 19672 23664 19700
rect 22520 19660 22526 19672
rect 23658 19660 23664 19672
rect 23716 19660 23722 19712
rect 1104 19610 28888 19632
rect 1104 19558 10214 19610
rect 10266 19558 10278 19610
rect 10330 19558 10342 19610
rect 10394 19558 10406 19610
rect 10458 19558 10470 19610
rect 10522 19558 19478 19610
rect 19530 19558 19542 19610
rect 19594 19558 19606 19610
rect 19658 19558 19670 19610
rect 19722 19558 19734 19610
rect 19786 19558 28888 19610
rect 1104 19536 28888 19558
rect 25130 19496 25136 19508
rect 25091 19468 25136 19496
rect 25130 19456 25136 19468
rect 25188 19456 25194 19508
rect 16850 19388 16856 19440
rect 16908 19428 16914 19440
rect 16945 19431 17003 19437
rect 16945 19428 16957 19431
rect 16908 19400 16957 19428
rect 16908 19388 16914 19400
rect 16945 19397 16957 19400
rect 16991 19397 17003 19431
rect 16945 19391 17003 19397
rect 17161 19431 17219 19437
rect 17161 19397 17173 19431
rect 17207 19428 17219 19431
rect 17402 19428 17408 19440
rect 17207 19400 17408 19428
rect 17207 19397 17219 19400
rect 17161 19391 17219 19397
rect 17402 19388 17408 19400
rect 17460 19388 17466 19440
rect 17957 19431 18015 19437
rect 17957 19397 17969 19431
rect 18003 19428 18015 19431
rect 19978 19428 19984 19440
rect 18003 19400 19984 19428
rect 18003 19397 18015 19400
rect 17957 19391 18015 19397
rect 19978 19388 19984 19400
rect 20036 19428 20042 19440
rect 20625 19431 20683 19437
rect 20625 19428 20637 19431
rect 20036 19400 20637 19428
rect 20036 19388 20042 19400
rect 20625 19397 20637 19400
rect 20671 19397 20683 19431
rect 20625 19391 20683 19397
rect 1394 19360 1400 19372
rect 1355 19332 1400 19360
rect 1394 19320 1400 19332
rect 1452 19320 1458 19372
rect 14274 19320 14280 19372
rect 14332 19360 14338 19372
rect 14829 19363 14887 19369
rect 14829 19360 14841 19363
rect 14332 19332 14841 19360
rect 14332 19320 14338 19332
rect 14829 19329 14841 19332
rect 14875 19329 14887 19363
rect 14829 19323 14887 19329
rect 14921 19363 14979 19369
rect 14921 19329 14933 19363
rect 14967 19360 14979 19363
rect 15194 19360 15200 19372
rect 14967 19332 15200 19360
rect 14967 19329 14979 19332
rect 14921 19323 14979 19329
rect 15194 19320 15200 19332
rect 15252 19320 15258 19372
rect 24486 19360 24492 19372
rect 24447 19332 24492 19360
rect 24486 19320 24492 19332
rect 24544 19320 24550 19372
rect 24673 19363 24731 19369
rect 24673 19329 24685 19363
rect 24719 19360 24731 19363
rect 25317 19363 25375 19369
rect 25317 19360 25329 19363
rect 24719 19332 25329 19360
rect 24719 19329 24731 19332
rect 24673 19323 24731 19329
rect 25317 19329 25329 19332
rect 25363 19329 25375 19363
rect 25317 19323 25375 19329
rect 26326 19320 26332 19372
rect 26384 19360 26390 19372
rect 26421 19363 26479 19369
rect 26421 19360 26433 19363
rect 26384 19332 26433 19360
rect 26384 19320 26390 19332
rect 26421 19329 26433 19332
rect 26467 19329 26479 19363
rect 26421 19323 26479 19329
rect 1578 19292 1584 19304
rect 1539 19264 1584 19292
rect 1578 19252 1584 19264
rect 1636 19252 1642 19304
rect 1854 19292 1860 19304
rect 1815 19264 1860 19292
rect 1854 19252 1860 19264
rect 1912 19252 1918 19304
rect 24026 19252 24032 19304
rect 24084 19292 24090 19304
rect 24305 19295 24363 19301
rect 24305 19292 24317 19295
rect 24084 19264 24317 19292
rect 24084 19252 24090 19264
rect 24305 19261 24317 19264
rect 24351 19261 24363 19295
rect 24305 19255 24363 19261
rect 19334 19224 19340 19236
rect 17144 19196 19340 19224
rect 16482 19116 16488 19168
rect 16540 19156 16546 19168
rect 17144 19165 17172 19196
rect 19334 19184 19340 19196
rect 19392 19184 19398 19236
rect 17129 19159 17187 19165
rect 17129 19156 17141 19159
rect 16540 19128 17141 19156
rect 16540 19116 16546 19128
rect 17129 19125 17141 19128
rect 17175 19125 17187 19159
rect 17310 19156 17316 19168
rect 17271 19128 17316 19156
rect 17129 19119 17187 19125
rect 17310 19116 17316 19128
rect 17368 19116 17374 19168
rect 17862 19156 17868 19168
rect 17823 19128 17868 19156
rect 17862 19116 17868 19128
rect 17920 19116 17926 19168
rect 20533 19159 20591 19165
rect 20533 19125 20545 19159
rect 20579 19156 20591 19159
rect 20990 19156 20996 19168
rect 20579 19128 20996 19156
rect 20579 19125 20591 19128
rect 20533 19119 20591 19125
rect 20990 19116 20996 19128
rect 21048 19116 21054 19168
rect 27430 19156 27436 19168
rect 27391 19128 27436 19156
rect 27430 19116 27436 19128
rect 27488 19116 27494 19168
rect 28077 19159 28135 19165
rect 28077 19125 28089 19159
rect 28123 19156 28135 19159
rect 28166 19156 28172 19168
rect 28123 19128 28172 19156
rect 28123 19125 28135 19128
rect 28077 19119 28135 19125
rect 28166 19116 28172 19128
rect 28224 19116 28230 19168
rect 1104 19066 28888 19088
rect 1104 19014 5582 19066
rect 5634 19014 5646 19066
rect 5698 19014 5710 19066
rect 5762 19014 5774 19066
rect 5826 19014 5838 19066
rect 5890 19014 14846 19066
rect 14898 19014 14910 19066
rect 14962 19014 14974 19066
rect 15026 19014 15038 19066
rect 15090 19014 15102 19066
rect 15154 19014 24110 19066
rect 24162 19014 24174 19066
rect 24226 19014 24238 19066
rect 24290 19014 24302 19066
rect 24354 19014 24366 19066
rect 24418 19014 28888 19066
rect 1104 18992 28888 19014
rect 1578 18912 1584 18964
rect 1636 18952 1642 18964
rect 1857 18955 1915 18961
rect 1857 18952 1869 18955
rect 1636 18924 1869 18952
rect 1636 18912 1642 18924
rect 1857 18921 1869 18924
rect 1903 18921 1915 18955
rect 17494 18952 17500 18964
rect 17455 18924 17500 18952
rect 1857 18915 1915 18921
rect 17494 18912 17500 18924
rect 17552 18912 17558 18964
rect 21818 18912 21824 18964
rect 21876 18952 21882 18964
rect 22005 18955 22063 18961
rect 22005 18952 22017 18955
rect 21876 18924 22017 18952
rect 21876 18912 21882 18924
rect 22005 18921 22017 18924
rect 22051 18921 22063 18955
rect 22005 18915 22063 18921
rect 24854 18884 24860 18896
rect 6886 18856 24860 18884
rect 6886 18816 6914 18856
rect 24854 18844 24860 18856
rect 24912 18844 24918 18896
rect 2240 18788 6914 18816
rect 17129 18819 17187 18825
rect 2240 18760 2268 18788
rect 17129 18785 17141 18819
rect 17175 18816 17187 18819
rect 17310 18816 17316 18828
rect 17175 18788 17316 18816
rect 17175 18785 17187 18788
rect 17129 18779 17187 18785
rect 17310 18776 17316 18788
rect 17368 18816 17374 18828
rect 17770 18816 17776 18828
rect 17368 18788 17776 18816
rect 17368 18776 17374 18788
rect 17770 18776 17776 18788
rect 17828 18776 17834 18828
rect 21361 18819 21419 18825
rect 21361 18785 21373 18819
rect 21407 18816 21419 18819
rect 27338 18816 27344 18828
rect 21407 18788 22048 18816
rect 27299 18788 27344 18816
rect 21407 18785 21419 18788
rect 21361 18779 21419 18785
rect 22020 18760 22048 18788
rect 27338 18776 27344 18788
rect 27396 18776 27402 18828
rect 27430 18776 27436 18828
rect 27488 18816 27494 18828
rect 28169 18819 28227 18825
rect 28169 18816 28181 18819
rect 27488 18788 28181 18816
rect 27488 18776 27494 18788
rect 28169 18785 28181 18788
rect 28215 18785 28227 18819
rect 28169 18779 28227 18785
rect 1949 18751 2007 18757
rect 1949 18717 1961 18751
rect 1995 18748 2007 18751
rect 2222 18748 2228 18760
rect 1995 18720 2228 18748
rect 1995 18717 2007 18720
rect 1949 18711 2007 18717
rect 2222 18708 2228 18720
rect 2280 18708 2286 18760
rect 2406 18748 2412 18760
rect 2367 18720 2412 18748
rect 2406 18708 2412 18720
rect 2464 18708 2470 18760
rect 16482 18748 16488 18760
rect 16443 18720 16488 18748
rect 16482 18708 16488 18720
rect 16540 18708 16546 18760
rect 18141 18751 18199 18757
rect 18141 18748 18153 18751
rect 17696 18720 18153 18748
rect 16298 18680 16304 18692
rect 16259 18652 16304 18680
rect 16298 18640 16304 18652
rect 16356 18640 16362 18692
rect 2593 18615 2651 18621
rect 2593 18581 2605 18615
rect 2639 18612 2651 18615
rect 12710 18612 12716 18624
rect 2639 18584 12716 18612
rect 2639 18581 2651 18584
rect 2593 18575 2651 18581
rect 12710 18572 12716 18584
rect 12768 18572 12774 18624
rect 17696 18621 17724 18720
rect 18141 18717 18153 18720
rect 18187 18717 18199 18751
rect 18141 18711 18199 18717
rect 21177 18751 21235 18757
rect 21177 18717 21189 18751
rect 21223 18748 21235 18751
rect 21266 18748 21272 18760
rect 21223 18720 21272 18748
rect 21223 18717 21235 18720
rect 21177 18711 21235 18717
rect 21266 18708 21272 18720
rect 21324 18708 21330 18760
rect 21910 18748 21916 18760
rect 21871 18720 21916 18748
rect 21910 18708 21916 18720
rect 21968 18708 21974 18760
rect 22002 18708 22008 18760
rect 22060 18748 22066 18760
rect 22189 18751 22247 18757
rect 22189 18748 22201 18751
rect 22060 18720 22201 18748
rect 22060 18708 22066 18720
rect 22189 18717 22201 18720
rect 22235 18717 22247 18751
rect 22189 18711 22247 18717
rect 27798 18640 27804 18692
rect 27856 18680 27862 18692
rect 27985 18683 28043 18689
rect 27985 18680 27997 18683
rect 27856 18652 27997 18680
rect 27856 18640 27862 18652
rect 27985 18649 27997 18652
rect 28031 18649 28043 18683
rect 27985 18643 28043 18649
rect 16669 18615 16727 18621
rect 16669 18581 16681 18615
rect 16715 18612 16727 18615
rect 17497 18615 17555 18621
rect 17497 18612 17509 18615
rect 16715 18584 17509 18612
rect 16715 18581 16727 18584
rect 16669 18575 16727 18581
rect 17497 18581 17509 18584
rect 17543 18581 17555 18615
rect 17497 18575 17555 18581
rect 17681 18615 17739 18621
rect 17681 18581 17693 18615
rect 17727 18581 17739 18615
rect 18322 18612 18328 18624
rect 18283 18584 18328 18612
rect 17681 18575 17739 18581
rect 18322 18572 18328 18584
rect 18380 18572 18386 18624
rect 22370 18612 22376 18624
rect 22331 18584 22376 18612
rect 22370 18572 22376 18584
rect 22428 18572 22434 18624
rect 1104 18522 28888 18544
rect 1104 18470 10214 18522
rect 10266 18470 10278 18522
rect 10330 18470 10342 18522
rect 10394 18470 10406 18522
rect 10458 18470 10470 18522
rect 10522 18470 19478 18522
rect 19530 18470 19542 18522
rect 19594 18470 19606 18522
rect 19658 18470 19670 18522
rect 19722 18470 19734 18522
rect 19786 18470 28888 18522
rect 1104 18448 28888 18470
rect 16298 18368 16304 18420
rect 16356 18408 16362 18420
rect 16669 18411 16727 18417
rect 16669 18408 16681 18411
rect 16356 18380 16681 18408
rect 16356 18368 16362 18380
rect 16669 18377 16681 18380
rect 16715 18377 16727 18411
rect 20806 18408 20812 18420
rect 16669 18371 16727 18377
rect 18156 18380 20812 18408
rect 18156 18340 18184 18380
rect 20806 18368 20812 18380
rect 20864 18368 20870 18420
rect 21910 18368 21916 18420
rect 21968 18408 21974 18420
rect 22925 18411 22983 18417
rect 22925 18408 22937 18411
rect 21968 18380 22937 18408
rect 21968 18368 21974 18380
rect 22925 18377 22937 18380
rect 22971 18377 22983 18411
rect 22925 18371 22983 18377
rect 25222 18368 25228 18420
rect 25280 18408 25286 18420
rect 25317 18411 25375 18417
rect 25317 18408 25329 18411
rect 25280 18380 25329 18408
rect 25280 18368 25286 18380
rect 25317 18377 25329 18380
rect 25363 18377 25375 18411
rect 27798 18408 27804 18420
rect 27759 18380 27804 18408
rect 25317 18371 25375 18377
rect 27798 18368 27804 18380
rect 27856 18368 27862 18420
rect 18322 18349 18328 18352
rect 18316 18340 18328 18349
rect 12452 18312 18184 18340
rect 18283 18312 18328 18340
rect 12452 18284 12480 18312
rect 18316 18303 18328 18312
rect 18322 18300 18328 18303
rect 18380 18300 18386 18352
rect 20824 18312 22048 18340
rect 12342 18272 12348 18284
rect 12303 18244 12348 18272
rect 12342 18232 12348 18244
rect 12400 18232 12406 18284
rect 12434 18232 12440 18284
rect 12492 18272 12498 18284
rect 13265 18275 13323 18281
rect 12492 18244 12537 18272
rect 12492 18232 12498 18244
rect 13265 18241 13277 18275
rect 13311 18272 13323 18275
rect 13354 18272 13360 18284
rect 13311 18244 13360 18272
rect 13311 18241 13323 18244
rect 13265 18235 13323 18241
rect 13354 18232 13360 18244
rect 13412 18232 13418 18284
rect 14366 18272 14372 18284
rect 14327 18244 14372 18272
rect 14366 18232 14372 18244
rect 14424 18232 14430 18284
rect 14550 18232 14556 18284
rect 14608 18272 14614 18284
rect 14645 18275 14703 18281
rect 14645 18272 14657 18275
rect 14608 18244 14657 18272
rect 14608 18232 14614 18244
rect 14645 18241 14657 18244
rect 14691 18241 14703 18275
rect 14826 18272 14832 18284
rect 14787 18244 14832 18272
rect 14645 18235 14703 18241
rect 14826 18232 14832 18244
rect 14884 18232 14890 18284
rect 16853 18275 16911 18281
rect 16853 18241 16865 18275
rect 16899 18241 16911 18275
rect 16853 18235 16911 18241
rect 14461 18207 14519 18213
rect 14461 18173 14473 18207
rect 14507 18204 14519 18207
rect 14734 18204 14740 18216
rect 14507 18176 14740 18204
rect 14507 18173 14519 18176
rect 14461 18167 14519 18173
rect 14734 18164 14740 18176
rect 14792 18164 14798 18216
rect 16868 18204 16896 18235
rect 16942 18232 16948 18284
rect 17000 18272 17006 18284
rect 17000 18244 17045 18272
rect 17000 18232 17006 18244
rect 17862 18232 17868 18284
rect 17920 18272 17926 18284
rect 20824 18281 20852 18312
rect 22020 18284 22048 18312
rect 22094 18300 22100 18352
rect 22152 18340 22158 18352
rect 22830 18340 22836 18352
rect 22152 18312 22232 18340
rect 22791 18312 22836 18340
rect 22152 18300 22158 18312
rect 18049 18275 18107 18281
rect 18049 18272 18061 18275
rect 17920 18244 18061 18272
rect 17920 18232 17926 18244
rect 18049 18241 18061 18244
rect 18095 18241 18107 18275
rect 18049 18235 18107 18241
rect 20809 18275 20867 18281
rect 20809 18241 20821 18275
rect 20855 18241 20867 18275
rect 20809 18235 20867 18241
rect 20993 18275 21051 18281
rect 20993 18241 21005 18275
rect 21039 18272 21051 18275
rect 21174 18272 21180 18284
rect 21039 18244 21180 18272
rect 21039 18241 21051 18244
rect 20993 18235 21051 18241
rect 21174 18232 21180 18244
rect 21232 18232 21238 18284
rect 22002 18272 22008 18284
rect 21963 18244 22008 18272
rect 22002 18232 22008 18244
rect 22060 18232 22066 18284
rect 22204 18281 22232 18312
rect 22830 18300 22836 18312
rect 22888 18300 22894 18352
rect 22189 18275 22247 18281
rect 22189 18241 22201 18275
rect 22235 18241 22247 18275
rect 22738 18272 22744 18284
rect 22699 18244 22744 18272
rect 22189 18235 22247 18241
rect 22738 18232 22744 18244
rect 22796 18232 22802 18284
rect 23842 18272 23848 18284
rect 23803 18244 23848 18272
rect 23842 18232 23848 18244
rect 23900 18232 23906 18284
rect 25409 18275 25467 18281
rect 25409 18241 25421 18275
rect 25455 18272 25467 18275
rect 25590 18272 25596 18284
rect 25455 18244 25596 18272
rect 25455 18241 25467 18244
rect 25409 18235 25467 18241
rect 25590 18232 25596 18244
rect 25648 18232 25654 18284
rect 27157 18275 27215 18281
rect 27157 18241 27169 18275
rect 27203 18272 27215 18275
rect 27246 18272 27252 18284
rect 27203 18244 27252 18272
rect 27203 18241 27215 18244
rect 27157 18235 27215 18241
rect 27246 18232 27252 18244
rect 27304 18272 27310 18284
rect 27614 18272 27620 18284
rect 27304 18244 27620 18272
rect 27304 18232 27310 18244
rect 27614 18232 27620 18244
rect 27672 18232 27678 18284
rect 27709 18275 27767 18281
rect 27709 18241 27721 18275
rect 27755 18272 27767 18275
rect 28442 18272 28448 18284
rect 27755 18244 28448 18272
rect 27755 18241 27767 18244
rect 27709 18235 27767 18241
rect 28442 18232 28448 18244
rect 28500 18272 28506 18284
rect 28718 18272 28724 18284
rect 28500 18244 28724 18272
rect 28500 18232 28506 18244
rect 28718 18232 28724 18244
rect 28776 18232 28782 18284
rect 17402 18204 17408 18216
rect 16868 18176 17408 18204
rect 17402 18164 17408 18176
rect 17460 18164 17466 18216
rect 21082 18204 21088 18216
rect 21043 18176 21088 18204
rect 21082 18164 21088 18176
rect 21140 18164 21146 18216
rect 22094 18164 22100 18216
rect 22152 18204 22158 18216
rect 22281 18207 22339 18213
rect 22281 18204 22293 18207
rect 22152 18176 22293 18204
rect 22152 18164 22158 18176
rect 22281 18173 22293 18176
rect 22327 18173 22339 18207
rect 23198 18204 23204 18216
rect 23159 18176 23204 18204
rect 22281 18167 22339 18173
rect 23198 18164 23204 18176
rect 23256 18164 23262 18216
rect 23474 18164 23480 18216
rect 23532 18204 23538 18216
rect 24026 18204 24032 18216
rect 23532 18176 24032 18204
rect 23532 18164 23538 18176
rect 24026 18164 24032 18176
rect 24084 18164 24090 18216
rect 24946 18164 24952 18216
rect 25004 18204 25010 18216
rect 25133 18207 25191 18213
rect 25133 18204 25145 18207
rect 25004 18176 25145 18204
rect 25004 18164 25010 18176
rect 25133 18173 25145 18176
rect 25179 18173 25191 18207
rect 25133 18167 25191 18173
rect 14550 18096 14556 18148
rect 14608 18136 14614 18148
rect 14608 18108 14653 18136
rect 14608 18096 14614 18108
rect 1394 18068 1400 18080
rect 1355 18040 1400 18068
rect 1394 18028 1400 18040
rect 1452 18028 1458 18080
rect 11238 18028 11244 18080
rect 11296 18068 11302 18080
rect 12161 18071 12219 18077
rect 12161 18068 12173 18071
rect 11296 18040 12173 18068
rect 11296 18028 11302 18040
rect 12161 18037 12173 18040
rect 12207 18037 12219 18071
rect 12161 18031 12219 18037
rect 13262 18028 13268 18080
rect 13320 18068 13326 18080
rect 13357 18071 13415 18077
rect 13357 18068 13369 18071
rect 13320 18040 13369 18068
rect 13320 18028 13326 18040
rect 13357 18037 13369 18040
rect 13403 18037 13415 18071
rect 13357 18031 13415 18037
rect 13725 18071 13783 18077
rect 13725 18037 13737 18071
rect 13771 18068 13783 18071
rect 14090 18068 14096 18080
rect 13771 18040 14096 18068
rect 13771 18037 13783 18040
rect 13725 18031 13783 18037
rect 14090 18028 14096 18040
rect 14148 18028 14154 18080
rect 14185 18071 14243 18077
rect 14185 18037 14197 18071
rect 14231 18068 14243 18071
rect 18322 18068 18328 18080
rect 14231 18040 18328 18068
rect 14231 18037 14243 18040
rect 14185 18031 14243 18037
rect 18322 18028 18328 18040
rect 18380 18028 18386 18080
rect 19334 18028 19340 18080
rect 19392 18068 19398 18080
rect 19429 18071 19487 18077
rect 19429 18068 19441 18071
rect 19392 18040 19441 18068
rect 19392 18028 19398 18040
rect 19429 18037 19441 18040
rect 19475 18037 19487 18071
rect 20622 18068 20628 18080
rect 20583 18040 20628 18068
rect 19429 18031 19487 18037
rect 20622 18028 20628 18040
rect 20680 18028 20686 18080
rect 21266 18028 21272 18080
rect 21324 18068 21330 18080
rect 21821 18071 21879 18077
rect 21821 18068 21833 18071
rect 21324 18040 21833 18068
rect 21324 18028 21330 18040
rect 21821 18037 21833 18040
rect 21867 18037 21879 18071
rect 21821 18031 21879 18037
rect 23566 18028 23572 18080
rect 23624 18068 23630 18080
rect 23661 18071 23719 18077
rect 23661 18068 23673 18071
rect 23624 18040 23673 18068
rect 23624 18028 23630 18040
rect 23661 18037 23673 18040
rect 23707 18037 23719 18071
rect 23661 18031 23719 18037
rect 25498 18028 25504 18080
rect 25556 18068 25562 18080
rect 25777 18071 25835 18077
rect 25777 18068 25789 18071
rect 25556 18040 25789 18068
rect 25556 18028 25562 18040
rect 25777 18037 25789 18040
rect 25823 18037 25835 18071
rect 25777 18031 25835 18037
rect 26510 18028 26516 18080
rect 26568 18068 26574 18080
rect 27065 18071 27123 18077
rect 27065 18068 27077 18071
rect 26568 18040 27077 18068
rect 26568 18028 26574 18040
rect 27065 18037 27077 18040
rect 27111 18037 27123 18071
rect 27065 18031 27123 18037
rect 1104 17978 28888 18000
rect 1104 17926 5582 17978
rect 5634 17926 5646 17978
rect 5698 17926 5710 17978
rect 5762 17926 5774 17978
rect 5826 17926 5838 17978
rect 5890 17926 14846 17978
rect 14898 17926 14910 17978
rect 14962 17926 14974 17978
rect 15026 17926 15038 17978
rect 15090 17926 15102 17978
rect 15154 17926 24110 17978
rect 24162 17926 24174 17978
rect 24226 17926 24238 17978
rect 24290 17926 24302 17978
rect 24354 17926 24366 17978
rect 24418 17926 28888 17978
rect 1104 17904 28888 17926
rect 16117 17867 16175 17873
rect 16117 17833 16129 17867
rect 16163 17864 16175 17867
rect 16666 17864 16672 17876
rect 16163 17836 16672 17864
rect 16163 17833 16175 17836
rect 16117 17827 16175 17833
rect 16666 17824 16672 17836
rect 16724 17824 16730 17876
rect 18601 17867 18659 17873
rect 18601 17833 18613 17867
rect 18647 17864 18659 17867
rect 18782 17864 18788 17876
rect 18647 17836 18788 17864
rect 18647 17833 18659 17836
rect 18601 17827 18659 17833
rect 18782 17824 18788 17836
rect 18840 17824 18846 17876
rect 23198 17824 23204 17876
rect 23256 17864 23262 17876
rect 23385 17867 23443 17873
rect 23385 17864 23397 17867
rect 23256 17836 23397 17864
rect 23256 17824 23262 17836
rect 23385 17833 23397 17836
rect 23431 17833 23443 17867
rect 23385 17827 23443 17833
rect 16298 17756 16304 17808
rect 16356 17796 16362 17808
rect 16485 17799 16543 17805
rect 16485 17796 16497 17799
rect 16356 17768 16497 17796
rect 16356 17756 16362 17768
rect 16485 17765 16497 17768
rect 16531 17765 16543 17799
rect 16485 17759 16543 17765
rect 26050 17756 26056 17808
rect 26108 17796 26114 17808
rect 26108 17768 26832 17796
rect 26108 17756 26114 17768
rect 1394 17728 1400 17740
rect 1355 17700 1400 17728
rect 1394 17688 1400 17700
rect 1452 17688 1458 17740
rect 2774 17728 2780 17740
rect 2735 17700 2780 17728
rect 2774 17688 2780 17700
rect 2832 17688 2838 17740
rect 14461 17731 14519 17737
rect 14461 17697 14473 17731
rect 14507 17728 14519 17731
rect 14734 17728 14740 17740
rect 14507 17700 14740 17728
rect 14507 17697 14519 17700
rect 14461 17691 14519 17697
rect 14734 17688 14740 17700
rect 14792 17688 14798 17740
rect 22005 17731 22063 17737
rect 22005 17728 22017 17731
rect 21008 17700 22017 17728
rect 21008 17672 21036 17700
rect 22005 17697 22017 17700
rect 22051 17728 22063 17731
rect 26510 17728 26516 17740
rect 22051 17700 22140 17728
rect 26471 17700 26516 17728
rect 22051 17697 22063 17700
rect 22005 17691 22063 17697
rect 11238 17660 11244 17672
rect 11199 17632 11244 17660
rect 11238 17620 11244 17632
rect 11296 17620 11302 17672
rect 11882 17660 11888 17672
rect 11843 17632 11888 17660
rect 11882 17620 11888 17632
rect 11940 17620 11946 17672
rect 14093 17663 14151 17669
rect 14093 17629 14105 17663
rect 14139 17660 14151 17663
rect 14182 17660 14188 17672
rect 14139 17632 14188 17660
rect 14139 17629 14151 17632
rect 14093 17623 14151 17629
rect 14182 17620 14188 17632
rect 14240 17620 14246 17672
rect 14366 17620 14372 17672
rect 14424 17660 14430 17672
rect 14553 17663 14611 17669
rect 14424 17632 14469 17660
rect 14424 17620 14430 17632
rect 14553 17629 14565 17663
rect 14599 17629 14611 17663
rect 14553 17623 14611 17629
rect 16945 17663 17003 17669
rect 16945 17629 16957 17663
rect 16991 17629 17003 17663
rect 18322 17660 18328 17672
rect 18283 17632 18328 17660
rect 16945 17623 17003 17629
rect 1581 17595 1639 17601
rect 1581 17561 1593 17595
rect 1627 17592 1639 17595
rect 1670 17592 1676 17604
rect 1627 17564 1676 17592
rect 1627 17561 1639 17564
rect 1581 17555 1639 17561
rect 1670 17552 1676 17564
rect 1728 17552 1734 17604
rect 12130 17595 12188 17601
rect 12130 17592 12142 17595
rect 11440 17564 12142 17592
rect 11440 17533 11468 17564
rect 12130 17561 12142 17564
rect 12176 17561 12188 17595
rect 12130 17555 12188 17561
rect 13906 17552 13912 17604
rect 13964 17592 13970 17604
rect 14568 17592 14596 17623
rect 16960 17592 16988 17623
rect 18322 17620 18328 17632
rect 18380 17620 18386 17672
rect 19797 17663 19855 17669
rect 19797 17629 19809 17663
rect 19843 17660 19855 17663
rect 20990 17660 20996 17672
rect 19843 17632 20996 17660
rect 19843 17629 19855 17632
rect 19797 17623 19855 17629
rect 20990 17620 20996 17632
rect 21048 17620 21054 17672
rect 22112 17660 22140 17700
rect 26510 17688 26516 17700
rect 26568 17688 26574 17740
rect 26804 17737 26832 17768
rect 26789 17731 26847 17737
rect 26789 17697 26801 17731
rect 26835 17697 26847 17731
rect 26789 17691 26847 17697
rect 24397 17663 24455 17669
rect 24397 17660 24409 17663
rect 22112 17632 24409 17660
rect 24397 17629 24409 17632
rect 24443 17629 24455 17663
rect 26326 17660 26332 17672
rect 26287 17632 26332 17660
rect 24397 17623 24455 17629
rect 26326 17620 26332 17632
rect 26384 17620 26390 17672
rect 13964 17564 14596 17592
rect 15948 17564 16988 17592
rect 18601 17595 18659 17601
rect 13964 17552 13970 17564
rect 11425 17527 11483 17533
rect 11425 17493 11437 17527
rect 11471 17493 11483 17527
rect 13262 17524 13268 17536
rect 13223 17496 13268 17524
rect 11425 17487 11483 17493
rect 13262 17484 13268 17496
rect 13320 17484 13326 17536
rect 14185 17527 14243 17533
rect 14185 17493 14197 17527
rect 14231 17524 14243 17527
rect 14274 17524 14280 17536
rect 14231 17496 14280 17524
rect 14231 17493 14243 17496
rect 14185 17487 14243 17493
rect 14274 17484 14280 17496
rect 14332 17484 14338 17536
rect 14642 17484 14648 17536
rect 14700 17524 14706 17536
rect 15948 17533 15976 17564
rect 18601 17561 18613 17595
rect 18647 17592 18659 17595
rect 19886 17592 19892 17604
rect 18647 17564 19892 17592
rect 18647 17561 18659 17564
rect 18601 17555 18659 17561
rect 19886 17552 19892 17564
rect 19944 17552 19950 17604
rect 20064 17595 20122 17601
rect 20064 17561 20076 17595
rect 20110 17592 20122 17595
rect 20622 17592 20628 17604
rect 20110 17564 20628 17592
rect 20110 17561 20122 17564
rect 20064 17555 20122 17561
rect 20622 17552 20628 17564
rect 20680 17552 20686 17604
rect 22272 17595 22330 17601
rect 22272 17561 22284 17595
rect 22318 17592 22330 17595
rect 22370 17592 22376 17604
rect 22318 17564 22376 17592
rect 22318 17561 22330 17564
rect 22272 17555 22330 17561
rect 22370 17552 22376 17564
rect 22428 17552 22434 17604
rect 23750 17552 23756 17604
rect 23808 17592 23814 17604
rect 24642 17595 24700 17601
rect 24642 17592 24654 17595
rect 23808 17564 24654 17592
rect 23808 17552 23814 17564
rect 24642 17561 24654 17564
rect 24688 17561 24700 17595
rect 24642 17555 24700 17561
rect 24854 17552 24860 17604
rect 24912 17592 24918 17604
rect 27522 17592 27528 17604
rect 24912 17564 27528 17592
rect 24912 17552 24918 17564
rect 27522 17552 27528 17564
rect 27580 17552 27586 17604
rect 14829 17527 14887 17533
rect 14829 17524 14841 17527
rect 14700 17496 14841 17524
rect 14700 17484 14706 17496
rect 14829 17493 14841 17496
rect 14875 17493 14887 17527
rect 14829 17487 14887 17493
rect 15933 17527 15991 17533
rect 15933 17493 15945 17527
rect 15979 17493 15991 17527
rect 16114 17524 16120 17536
rect 16075 17496 16120 17524
rect 15933 17487 15991 17493
rect 16114 17484 16120 17496
rect 16172 17484 16178 17536
rect 17129 17527 17187 17533
rect 17129 17493 17141 17527
rect 17175 17524 17187 17527
rect 17310 17524 17316 17536
rect 17175 17496 17316 17524
rect 17175 17493 17187 17496
rect 17129 17487 17187 17493
rect 17310 17484 17316 17496
rect 17368 17484 17374 17536
rect 18046 17484 18052 17536
rect 18104 17524 18110 17536
rect 18417 17527 18475 17533
rect 18417 17524 18429 17527
rect 18104 17496 18429 17524
rect 18104 17484 18110 17496
rect 18417 17493 18429 17496
rect 18463 17493 18475 17527
rect 18417 17487 18475 17493
rect 21177 17527 21235 17533
rect 21177 17493 21189 17527
rect 21223 17524 21235 17527
rect 21358 17524 21364 17536
rect 21223 17496 21364 17524
rect 21223 17493 21235 17496
rect 21177 17487 21235 17493
rect 21358 17484 21364 17496
rect 21416 17484 21422 17536
rect 25590 17484 25596 17536
rect 25648 17524 25654 17536
rect 25777 17527 25835 17533
rect 25777 17524 25789 17527
rect 25648 17496 25789 17524
rect 25648 17484 25654 17496
rect 25777 17493 25789 17496
rect 25823 17493 25835 17527
rect 25777 17487 25835 17493
rect 1104 17434 28888 17456
rect 1104 17382 10214 17434
rect 10266 17382 10278 17434
rect 10330 17382 10342 17434
rect 10394 17382 10406 17434
rect 10458 17382 10470 17434
rect 10522 17382 19478 17434
rect 19530 17382 19542 17434
rect 19594 17382 19606 17434
rect 19658 17382 19670 17434
rect 19722 17382 19734 17434
rect 19786 17382 28888 17434
rect 1104 17360 28888 17382
rect 1670 17320 1676 17332
rect 1631 17292 1676 17320
rect 1670 17280 1676 17292
rect 1728 17280 1734 17332
rect 12253 17323 12311 17329
rect 12253 17289 12265 17323
rect 12299 17320 12311 17323
rect 12342 17320 12348 17332
rect 12299 17292 12348 17320
rect 12299 17289 12311 17292
rect 12253 17283 12311 17289
rect 12342 17280 12348 17292
rect 12400 17280 12406 17332
rect 12621 17323 12679 17329
rect 12621 17289 12633 17323
rect 12667 17320 12679 17323
rect 13262 17320 13268 17332
rect 12667 17292 13268 17320
rect 12667 17289 12679 17292
rect 12621 17283 12679 17289
rect 13262 17280 13268 17292
rect 13320 17280 13326 17332
rect 13906 17320 13912 17332
rect 13867 17292 13912 17320
rect 13906 17280 13912 17292
rect 13964 17280 13970 17332
rect 14550 17280 14556 17332
rect 14608 17320 14614 17332
rect 14645 17323 14703 17329
rect 14645 17320 14657 17323
rect 14608 17292 14657 17320
rect 14608 17280 14614 17292
rect 14645 17289 14657 17292
rect 14691 17289 14703 17323
rect 14645 17283 14703 17289
rect 14734 17280 14740 17332
rect 14792 17320 14798 17332
rect 15473 17323 15531 17329
rect 15473 17320 15485 17323
rect 14792 17292 15485 17320
rect 14792 17280 14798 17292
rect 15473 17289 15485 17292
rect 15519 17289 15531 17323
rect 15473 17283 15531 17289
rect 20993 17323 21051 17329
rect 20993 17289 21005 17323
rect 21039 17320 21051 17323
rect 21082 17320 21088 17332
rect 21039 17292 21088 17320
rect 21039 17289 21051 17292
rect 20993 17283 21051 17289
rect 21082 17280 21088 17292
rect 21140 17280 21146 17332
rect 21913 17323 21971 17329
rect 21913 17289 21925 17323
rect 21959 17320 21971 17323
rect 22186 17320 22192 17332
rect 21959 17292 22192 17320
rect 21959 17289 21971 17292
rect 21913 17283 21971 17289
rect 22186 17280 22192 17292
rect 22244 17320 22250 17332
rect 22830 17320 22836 17332
rect 22244 17292 22836 17320
rect 22244 17280 22250 17292
rect 22830 17280 22836 17292
rect 22888 17280 22894 17332
rect 23477 17323 23535 17329
rect 23477 17289 23489 17323
rect 23523 17320 23535 17323
rect 23842 17320 23848 17332
rect 23523 17292 23848 17320
rect 23523 17289 23535 17292
rect 23477 17283 23535 17289
rect 23842 17280 23848 17292
rect 23900 17280 23906 17332
rect 26326 17280 26332 17332
rect 26384 17320 26390 17332
rect 27525 17323 27583 17329
rect 27525 17320 27537 17323
rect 26384 17292 27537 17320
rect 26384 17280 26390 17292
rect 27525 17289 27537 17292
rect 27571 17289 27583 17323
rect 27525 17283 27583 17289
rect 13354 17212 13360 17264
rect 13412 17252 13418 17264
rect 13449 17255 13507 17261
rect 13449 17252 13461 17255
rect 13412 17224 13461 17252
rect 13412 17212 13418 17224
rect 13449 17221 13461 17224
rect 13495 17221 13507 17255
rect 13449 17215 13507 17221
rect 14090 17212 14096 17264
rect 14148 17252 14154 17264
rect 14854 17255 14912 17261
rect 14854 17252 14866 17255
rect 14148 17224 14866 17252
rect 14148 17212 14154 17224
rect 14854 17221 14866 17224
rect 14900 17221 14912 17255
rect 17037 17255 17095 17261
rect 17037 17252 17049 17255
rect 14854 17215 14912 17221
rect 15488 17224 17049 17252
rect 1762 17184 1768 17196
rect 1723 17156 1768 17184
rect 1762 17144 1768 17156
rect 1820 17144 1826 17196
rect 14369 17187 14427 17193
rect 14369 17153 14381 17187
rect 14415 17184 14427 17187
rect 14642 17184 14648 17196
rect 14415 17156 14648 17184
rect 14415 17153 14427 17156
rect 14369 17147 14427 17153
rect 14642 17144 14648 17156
rect 14700 17144 14706 17196
rect 14737 17187 14795 17193
rect 14737 17153 14749 17187
rect 14783 17184 14795 17187
rect 15488 17184 15516 17224
rect 17037 17221 17049 17224
rect 17083 17221 17095 17255
rect 22738 17252 22744 17264
rect 17037 17215 17095 17221
rect 20824 17224 22744 17252
rect 14783 17156 15516 17184
rect 14783 17153 14795 17156
rect 14737 17147 14795 17153
rect 6546 17076 6552 17128
rect 6604 17116 6610 17128
rect 12713 17119 12771 17125
rect 12713 17116 12725 17119
rect 6604 17088 12725 17116
rect 6604 17076 6610 17088
rect 12713 17085 12725 17088
rect 12759 17085 12771 17119
rect 12894 17116 12900 17128
rect 12855 17088 12900 17116
rect 12713 17079 12771 17085
rect 12894 17076 12900 17088
rect 12952 17076 12958 17128
rect 14458 17076 14464 17128
rect 14516 17116 14522 17128
rect 14752 17116 14780 17147
rect 15562 17144 15568 17196
rect 15620 17184 15626 17196
rect 16669 17187 16727 17193
rect 16669 17184 16681 17187
rect 15620 17156 16681 17184
rect 15620 17144 15626 17156
rect 16669 17153 16681 17156
rect 16715 17153 16727 17187
rect 16850 17184 16856 17196
rect 16811 17156 16856 17184
rect 16669 17147 16727 17153
rect 16850 17144 16856 17156
rect 16908 17144 16914 17196
rect 20162 17184 20168 17196
rect 20075 17156 20168 17184
rect 20162 17144 20168 17156
rect 20220 17184 20226 17196
rect 20622 17184 20628 17196
rect 20220 17156 20628 17184
rect 20220 17144 20226 17156
rect 20622 17144 20628 17156
rect 20680 17144 20686 17196
rect 20824 17193 20852 17224
rect 21836 17193 21864 17224
rect 22738 17212 22744 17224
rect 22796 17212 22802 17264
rect 23198 17212 23204 17264
rect 23256 17252 23262 17264
rect 23937 17255 23995 17261
rect 23937 17252 23949 17255
rect 23256 17224 23949 17252
rect 23256 17212 23262 17224
rect 23937 17221 23949 17224
rect 23983 17221 23995 17255
rect 23937 17215 23995 17221
rect 26145 17255 26203 17261
rect 26145 17221 26157 17255
rect 26191 17252 26203 17255
rect 27154 17252 27160 17264
rect 26191 17224 27160 17252
rect 26191 17221 26203 17224
rect 26145 17215 26203 17221
rect 27154 17212 27160 17224
rect 27212 17212 27218 17264
rect 27430 17252 27436 17264
rect 27264 17224 27436 17252
rect 20809 17187 20867 17193
rect 20809 17153 20821 17187
rect 20855 17153 20867 17187
rect 20809 17147 20867 17153
rect 20901 17187 20959 17193
rect 20901 17153 20913 17187
rect 20947 17184 20959 17187
rect 21821 17187 21879 17193
rect 20947 17156 21496 17184
rect 20947 17153 20959 17156
rect 20901 17147 20959 17153
rect 14516 17088 14780 17116
rect 14516 17076 14522 17088
rect 15470 17076 15476 17128
rect 15528 17116 15534 17128
rect 15933 17119 15991 17125
rect 15933 17116 15945 17119
rect 15528 17088 15945 17116
rect 15528 17076 15534 17088
rect 15933 17085 15945 17088
rect 15979 17116 15991 17119
rect 18138 17116 18144 17128
rect 15979 17088 18144 17116
rect 15979 17085 15991 17088
rect 15933 17079 15991 17085
rect 18138 17076 18144 17088
rect 18196 17076 18202 17128
rect 21269 17119 21327 17125
rect 21269 17085 21281 17119
rect 21315 17116 21327 17119
rect 21358 17116 21364 17128
rect 21315 17088 21364 17116
rect 21315 17085 21327 17088
rect 21269 17079 21327 17085
rect 21358 17076 21364 17088
rect 21416 17076 21422 17128
rect 21468 17116 21496 17156
rect 21821 17153 21833 17187
rect 21867 17153 21879 17187
rect 21821 17147 21879 17153
rect 22094 17144 22100 17196
rect 22152 17184 22158 17196
rect 23845 17187 23903 17193
rect 22152 17156 22197 17184
rect 22152 17144 22158 17156
rect 23845 17153 23857 17187
rect 23891 17184 23903 17187
rect 25590 17184 25596 17196
rect 23891 17156 25596 17184
rect 23891 17153 23903 17156
rect 23845 17147 23903 17153
rect 25590 17144 25596 17156
rect 25648 17144 25654 17196
rect 25685 17187 25743 17193
rect 25685 17153 25697 17187
rect 25731 17153 25743 17187
rect 25685 17147 25743 17153
rect 25777 17187 25835 17193
rect 25777 17153 25789 17187
rect 25823 17153 25835 17187
rect 25777 17147 25835 17153
rect 22186 17116 22192 17128
rect 21468 17088 22192 17116
rect 22186 17076 22192 17088
rect 22244 17076 22250 17128
rect 22281 17119 22339 17125
rect 22281 17085 22293 17119
rect 22327 17116 22339 17119
rect 22830 17116 22836 17128
rect 22327 17088 22836 17116
rect 22327 17085 22339 17088
rect 22281 17079 22339 17085
rect 22830 17076 22836 17088
rect 22888 17076 22894 17128
rect 23658 17076 23664 17128
rect 23716 17116 23722 17128
rect 24029 17119 24087 17125
rect 24029 17116 24041 17119
rect 23716 17088 24041 17116
rect 23716 17076 23722 17088
rect 24029 17085 24041 17088
rect 24075 17085 24087 17119
rect 24029 17079 24087 17085
rect 13262 17008 13268 17060
rect 13320 17048 13326 17060
rect 13725 17051 13783 17057
rect 13725 17048 13737 17051
rect 13320 17020 13737 17048
rect 13320 17008 13326 17020
rect 13725 17017 13737 17020
rect 13771 17017 13783 17051
rect 13725 17011 13783 17017
rect 13998 17008 14004 17060
rect 14056 17048 14062 17060
rect 15562 17048 15568 17060
rect 14056 17020 15568 17048
rect 14056 17008 14062 17020
rect 15562 17008 15568 17020
rect 15620 17008 15626 17060
rect 15013 16983 15071 16989
rect 15013 16949 15025 16983
rect 15059 16980 15071 16983
rect 17954 16980 17960 16992
rect 15059 16952 17960 16980
rect 15059 16949 15071 16952
rect 15013 16943 15071 16949
rect 17954 16940 17960 16952
rect 18012 16940 18018 16992
rect 20254 16980 20260 16992
rect 20215 16952 20260 16980
rect 20254 16940 20260 16952
rect 20312 16940 20318 16992
rect 25700 16980 25728 17147
rect 25792 17048 25820 17147
rect 25866 17144 25872 17196
rect 25924 17184 25930 17196
rect 25961 17187 26019 17193
rect 25961 17184 25973 17187
rect 25924 17156 25973 17184
rect 25924 17144 25930 17156
rect 25961 17153 25973 17156
rect 26007 17153 26019 17187
rect 25961 17147 26019 17153
rect 26234 17144 26240 17196
rect 26292 17184 26298 17196
rect 26973 17187 27031 17193
rect 26973 17184 26985 17187
rect 26292 17156 26985 17184
rect 26292 17144 26298 17156
rect 26973 17153 26985 17156
rect 27019 17153 27031 17187
rect 26973 17147 27031 17153
rect 27062 17144 27068 17196
rect 27120 17184 27126 17196
rect 27264 17193 27292 17224
rect 27430 17212 27436 17224
rect 27488 17212 27494 17264
rect 27249 17187 27307 17193
rect 27120 17156 27165 17184
rect 27120 17144 27126 17156
rect 27249 17153 27261 17187
rect 27295 17153 27307 17187
rect 27249 17147 27307 17153
rect 27341 17187 27399 17193
rect 27341 17153 27353 17187
rect 27387 17153 27399 17187
rect 27341 17147 27399 17153
rect 26326 17076 26332 17128
rect 26384 17116 26390 17128
rect 27356 17116 27384 17147
rect 27614 17144 27620 17196
rect 27672 17184 27678 17196
rect 27985 17187 28043 17193
rect 27985 17184 27997 17187
rect 27672 17156 27997 17184
rect 27672 17144 27678 17156
rect 27985 17153 27997 17156
rect 28031 17153 28043 17187
rect 27985 17147 28043 17153
rect 26384 17088 27384 17116
rect 26384 17076 26390 17088
rect 27338 17048 27344 17060
rect 25792 17020 27344 17048
rect 27338 17008 27344 17020
rect 27396 17008 27402 17060
rect 26326 16980 26332 16992
rect 25700 16952 26332 16980
rect 26326 16940 26332 16952
rect 26384 16940 26390 16992
rect 27982 16940 27988 16992
rect 28040 16980 28046 16992
rect 28077 16983 28135 16989
rect 28077 16980 28089 16983
rect 28040 16952 28089 16980
rect 28040 16940 28046 16952
rect 28077 16949 28089 16952
rect 28123 16949 28135 16983
rect 28077 16943 28135 16949
rect 1104 16890 28888 16912
rect 1104 16838 5582 16890
rect 5634 16838 5646 16890
rect 5698 16838 5710 16890
rect 5762 16838 5774 16890
rect 5826 16838 5838 16890
rect 5890 16838 14846 16890
rect 14898 16838 14910 16890
rect 14962 16838 14974 16890
rect 15026 16838 15038 16890
rect 15090 16838 15102 16890
rect 15154 16838 24110 16890
rect 24162 16838 24174 16890
rect 24226 16838 24238 16890
rect 24290 16838 24302 16890
rect 24354 16838 24366 16890
rect 24418 16838 28888 16890
rect 1104 16816 28888 16838
rect 14182 16736 14188 16788
rect 14240 16776 14246 16788
rect 14240 16748 14504 16776
rect 14240 16736 14246 16748
rect 14182 16640 14188 16652
rect 14143 16612 14188 16640
rect 14182 16600 14188 16612
rect 14240 16600 14246 16652
rect 14274 16600 14280 16652
rect 14332 16640 14338 16652
rect 14332 16612 14412 16640
rect 14332 16600 14338 16612
rect 14090 16572 14096 16584
rect 14051 16544 14096 16572
rect 14090 16532 14096 16544
rect 14148 16532 14154 16584
rect 14384 16581 14412 16612
rect 14476 16581 14504 16748
rect 14550 16736 14556 16788
rect 14608 16776 14614 16788
rect 14645 16779 14703 16785
rect 14645 16776 14657 16779
rect 14608 16748 14657 16776
rect 14608 16736 14614 16748
rect 14645 16745 14657 16748
rect 14691 16745 14703 16779
rect 14645 16739 14703 16745
rect 15749 16779 15807 16785
rect 15749 16745 15761 16779
rect 15795 16776 15807 16779
rect 16114 16776 16120 16788
rect 15795 16748 16120 16776
rect 15795 16745 15807 16748
rect 15749 16739 15807 16745
rect 16114 16736 16120 16748
rect 16172 16736 16178 16788
rect 17402 16736 17408 16788
rect 17460 16776 17466 16788
rect 18049 16779 18107 16785
rect 18049 16776 18061 16779
rect 17460 16748 18061 16776
rect 17460 16736 17466 16748
rect 18049 16745 18061 16748
rect 18095 16745 18107 16779
rect 18049 16739 18107 16745
rect 18138 16736 18144 16788
rect 18196 16776 18202 16788
rect 18233 16779 18291 16785
rect 18233 16776 18245 16779
rect 18196 16748 18245 16776
rect 18196 16736 18202 16748
rect 18233 16745 18245 16748
rect 18279 16745 18291 16779
rect 23750 16776 23756 16788
rect 23711 16748 23756 16776
rect 18233 16739 18291 16745
rect 23750 16736 23756 16748
rect 23808 16736 23814 16788
rect 26970 16776 26976 16788
rect 25148 16748 26976 16776
rect 20533 16711 20591 16717
rect 20533 16677 20545 16711
rect 20579 16708 20591 16711
rect 21174 16708 21180 16720
rect 20579 16680 21180 16708
rect 20579 16677 20591 16680
rect 20533 16671 20591 16677
rect 21174 16668 21180 16680
rect 21232 16668 21238 16720
rect 15289 16643 15347 16649
rect 15289 16640 15301 16643
rect 15212 16612 15301 16640
rect 14369 16575 14427 16581
rect 14369 16541 14381 16575
rect 14415 16541 14427 16575
rect 14369 16535 14427 16541
rect 14461 16575 14519 16581
rect 14461 16541 14473 16575
rect 14507 16541 14519 16575
rect 14461 16535 14519 16541
rect 15212 16436 15240 16612
rect 15289 16609 15301 16612
rect 15335 16609 15347 16643
rect 15470 16640 15476 16652
rect 15431 16612 15476 16640
rect 15289 16603 15347 16609
rect 15470 16600 15476 16612
rect 15528 16600 15534 16652
rect 17586 16600 17592 16652
rect 17644 16640 17650 16652
rect 17862 16640 17868 16652
rect 17644 16612 17868 16640
rect 17644 16600 17650 16612
rect 17862 16600 17868 16612
rect 17920 16600 17926 16652
rect 19334 16640 19340 16652
rect 19247 16612 19340 16640
rect 15378 16572 15384 16584
rect 15339 16544 15384 16572
rect 15378 16532 15384 16544
rect 15436 16532 15442 16584
rect 15565 16575 15623 16581
rect 15565 16541 15577 16575
rect 15611 16541 15623 16575
rect 15565 16535 15623 16541
rect 15580 16504 15608 16535
rect 17310 16532 17316 16584
rect 17368 16581 17374 16584
rect 19260 16581 19288 16612
rect 19334 16600 19340 16612
rect 19392 16640 19398 16652
rect 19978 16640 19984 16652
rect 19392 16612 19984 16640
rect 19392 16600 19398 16612
rect 19978 16600 19984 16612
rect 20036 16600 20042 16652
rect 20806 16600 20812 16652
rect 20864 16640 20870 16652
rect 20993 16643 21051 16649
rect 20993 16640 21005 16643
rect 20864 16612 21005 16640
rect 20864 16600 20870 16612
rect 20993 16609 21005 16612
rect 21039 16609 21051 16643
rect 25148 16640 25176 16748
rect 26970 16736 26976 16748
rect 27028 16736 27034 16788
rect 25593 16711 25651 16717
rect 25593 16677 25605 16711
rect 25639 16708 25651 16711
rect 26326 16708 26332 16720
rect 25639 16680 26332 16708
rect 25639 16677 25651 16680
rect 25593 16671 25651 16677
rect 26326 16668 26332 16680
rect 26384 16668 26390 16720
rect 27982 16640 27988 16652
rect 20993 16603 21051 16609
rect 25056 16612 25176 16640
rect 27943 16612 27988 16640
rect 17368 16572 17380 16581
rect 19245 16575 19303 16581
rect 17368 16544 17413 16572
rect 17368 16535 17380 16544
rect 19245 16541 19257 16575
rect 19291 16541 19303 16575
rect 19245 16535 19303 16541
rect 17368 16532 17374 16535
rect 20254 16532 20260 16584
rect 20312 16572 20318 16584
rect 20349 16575 20407 16581
rect 20349 16572 20361 16575
rect 20312 16544 20361 16572
rect 20312 16532 20318 16544
rect 20349 16541 20361 16544
rect 20395 16572 20407 16575
rect 21177 16575 21235 16581
rect 21177 16572 21189 16575
rect 20395 16544 21189 16572
rect 20395 16541 20407 16544
rect 20349 16535 20407 16541
rect 21177 16541 21189 16544
rect 21223 16541 21235 16575
rect 23566 16572 23572 16584
rect 23527 16544 23572 16572
rect 21177 16535 21235 16541
rect 23566 16532 23572 16544
rect 23624 16532 23630 16584
rect 25056 16581 25084 16612
rect 27982 16600 27988 16612
rect 28040 16600 28046 16652
rect 28166 16640 28172 16652
rect 28127 16612 28172 16640
rect 28166 16600 28172 16612
rect 28224 16600 28230 16652
rect 25041 16575 25099 16581
rect 25041 16541 25053 16575
rect 25087 16541 25099 16575
rect 25498 16572 25504 16584
rect 25459 16544 25504 16572
rect 25041 16535 25099 16541
rect 25498 16532 25504 16544
rect 25556 16532 25562 16584
rect 25682 16572 25688 16584
rect 25643 16544 25688 16572
rect 25682 16532 25688 16544
rect 25740 16532 25746 16584
rect 25774 16532 25780 16584
rect 25832 16572 25838 16584
rect 26329 16575 26387 16581
rect 26329 16572 26341 16575
rect 25832 16544 26341 16572
rect 25832 16532 25838 16544
rect 26329 16541 26341 16544
rect 26375 16541 26387 16575
rect 26329 16535 26387 16541
rect 15654 16504 15660 16516
rect 15567 16476 15660 16504
rect 15654 16464 15660 16476
rect 15712 16504 15718 16516
rect 18201 16507 18259 16513
rect 18201 16504 18213 16507
rect 15712 16476 18213 16504
rect 15712 16464 15718 16476
rect 18201 16473 18213 16476
rect 18247 16473 18259 16507
rect 18201 16467 18259 16473
rect 18417 16507 18475 16513
rect 18417 16473 18429 16507
rect 18463 16473 18475 16507
rect 18417 16467 18475 16473
rect 24949 16507 25007 16513
rect 24949 16473 24961 16507
rect 24995 16504 25007 16507
rect 24995 16476 26004 16504
rect 24995 16473 25007 16476
rect 24949 16467 25007 16473
rect 16206 16436 16212 16448
rect 15212 16408 16212 16436
rect 16206 16396 16212 16408
rect 16264 16436 16270 16448
rect 18432 16436 18460 16467
rect 19334 16436 19340 16448
rect 16264 16408 18460 16436
rect 19295 16408 19340 16436
rect 16264 16396 16270 16408
rect 19334 16396 19340 16408
rect 19392 16396 19398 16448
rect 25976 16436 26004 16476
rect 27062 16436 27068 16448
rect 25976 16408 27068 16436
rect 27062 16396 27068 16408
rect 27120 16396 27126 16448
rect 1104 16346 28888 16368
rect 1104 16294 10214 16346
rect 10266 16294 10278 16346
rect 10330 16294 10342 16346
rect 10394 16294 10406 16346
rect 10458 16294 10470 16346
rect 10522 16294 19478 16346
rect 19530 16294 19542 16346
rect 19594 16294 19606 16346
rect 19658 16294 19670 16346
rect 19722 16294 19734 16346
rect 19786 16294 28888 16346
rect 1104 16272 28888 16294
rect 7282 16192 7288 16244
rect 7340 16232 7346 16244
rect 12805 16235 12863 16241
rect 12805 16232 12817 16235
rect 7340 16204 12817 16232
rect 7340 16192 7346 16204
rect 12805 16201 12817 16204
rect 12851 16201 12863 16235
rect 15654 16232 15660 16244
rect 15615 16204 15660 16232
rect 12805 16195 12863 16201
rect 15654 16192 15660 16204
rect 15712 16192 15718 16244
rect 18046 16232 18052 16244
rect 18007 16204 18052 16232
rect 18046 16192 18052 16204
rect 18104 16192 18110 16244
rect 19797 16235 19855 16241
rect 19797 16201 19809 16235
rect 19843 16232 19855 16235
rect 19886 16232 19892 16244
rect 19843 16204 19892 16232
rect 19843 16201 19855 16204
rect 19797 16195 19855 16201
rect 19886 16192 19892 16204
rect 19944 16192 19950 16244
rect 27338 16232 27344 16244
rect 25792 16204 27344 16232
rect 18417 16167 18475 16173
rect 18417 16133 18429 16167
rect 18463 16164 18475 16167
rect 19242 16164 19248 16176
rect 18463 16136 19248 16164
rect 18463 16133 18475 16136
rect 18417 16127 18475 16133
rect 19242 16124 19248 16136
rect 19300 16164 19306 16176
rect 25792 16164 25820 16204
rect 27338 16192 27344 16204
rect 27396 16192 27402 16244
rect 19300 16136 19472 16164
rect 19300 16124 19306 16136
rect 12713 16099 12771 16105
rect 12713 16065 12725 16099
rect 12759 16096 12771 16099
rect 13354 16096 13360 16108
rect 12759 16068 13360 16096
rect 12759 16065 12771 16068
rect 12713 16059 12771 16065
rect 13354 16056 13360 16068
rect 13412 16056 13418 16108
rect 15473 16099 15531 16105
rect 15473 16065 15485 16099
rect 15519 16096 15531 16099
rect 16022 16096 16028 16108
rect 15519 16068 16028 16096
rect 15519 16065 15531 16068
rect 15473 16059 15531 16065
rect 16022 16056 16028 16068
rect 16080 16056 16086 16108
rect 16206 16056 16212 16108
rect 16264 16096 16270 16108
rect 19444 16105 19472 16136
rect 25700 16136 25820 16164
rect 17129 16099 17187 16105
rect 17129 16096 17141 16099
rect 16264 16068 17141 16096
rect 16264 16056 16270 16068
rect 17129 16065 17141 16068
rect 17175 16065 17187 16099
rect 19153 16099 19211 16105
rect 19153 16096 19165 16099
rect 17129 16059 17187 16065
rect 18708 16068 19165 16096
rect 18708 16040 18736 16068
rect 19153 16065 19165 16068
rect 19199 16065 19211 16099
rect 19153 16059 19211 16065
rect 19337 16099 19395 16105
rect 19337 16065 19349 16099
rect 19383 16065 19395 16099
rect 19337 16059 19395 16065
rect 19429 16099 19487 16105
rect 19429 16065 19441 16099
rect 19475 16065 19487 16099
rect 19429 16059 19487 16065
rect 19521 16099 19579 16105
rect 19521 16065 19533 16099
rect 19567 16096 19579 16099
rect 20714 16096 20720 16108
rect 19567 16068 20720 16096
rect 19567 16065 19579 16068
rect 19521 16059 19579 16065
rect 12894 15988 12900 16040
rect 12952 16028 12958 16040
rect 12989 16031 13047 16037
rect 12989 16028 13001 16031
rect 12952 16000 13001 16028
rect 12952 15988 12958 16000
rect 12989 15997 13001 16000
rect 13035 15997 13047 16031
rect 12989 15991 13047 15997
rect 13004 15960 13032 15991
rect 14550 15988 14556 16040
rect 14608 16028 14614 16040
rect 15289 16031 15347 16037
rect 15289 16028 15301 16031
rect 14608 16000 15301 16028
rect 14608 15988 14614 16000
rect 15289 15997 15301 16000
rect 15335 15997 15347 16031
rect 15289 15991 15347 15997
rect 17589 16031 17647 16037
rect 17589 15997 17601 16031
rect 17635 16028 17647 16031
rect 18208 16031 18266 16037
rect 18208 16028 18220 16031
rect 17635 16000 18220 16028
rect 17635 15997 17647 16000
rect 17589 15991 17647 15997
rect 18208 15997 18220 16000
rect 18254 15997 18266 16031
rect 18208 15991 18266 15997
rect 18325 16031 18383 16037
rect 18325 15997 18337 16031
rect 18371 15997 18383 16031
rect 18690 16028 18696 16040
rect 18651 16000 18696 16028
rect 18325 15991 18383 15997
rect 16482 15960 16488 15972
rect 13004 15932 16488 15960
rect 16482 15920 16488 15932
rect 16540 15920 16546 15972
rect 18340 15960 18368 15991
rect 18690 15988 18696 16000
rect 18748 15988 18754 16040
rect 19352 16028 19380 16059
rect 20714 16056 20720 16068
rect 20772 16056 20778 16108
rect 25700 16105 25728 16136
rect 25866 16124 25872 16176
rect 25924 16164 25930 16176
rect 26973 16167 27031 16173
rect 26973 16164 26985 16167
rect 25924 16136 26985 16164
rect 25924 16124 25930 16136
rect 25685 16099 25743 16105
rect 25685 16065 25697 16099
rect 25731 16065 25743 16099
rect 25685 16059 25743 16065
rect 25774 16056 25780 16108
rect 25832 16096 25838 16108
rect 25976 16105 26004 16136
rect 26973 16133 26985 16136
rect 27019 16133 27031 16167
rect 28074 16164 28080 16176
rect 28035 16136 28080 16164
rect 26973 16127 27031 16133
rect 28074 16124 28080 16136
rect 28132 16124 28138 16176
rect 25961 16099 26019 16105
rect 25832 16068 25877 16096
rect 25832 16056 25838 16068
rect 25961 16065 25973 16099
rect 26007 16065 26019 16099
rect 25961 16059 26019 16065
rect 26053 16099 26111 16105
rect 26053 16065 26065 16099
rect 26099 16096 26111 16099
rect 26234 16096 26240 16108
rect 26099 16068 26240 16096
rect 26099 16065 26111 16068
rect 26053 16059 26111 16065
rect 26234 16056 26240 16068
rect 26292 16056 26298 16108
rect 27249 16099 27307 16105
rect 27249 16096 27261 16099
rect 26344 16068 27261 16096
rect 19886 16028 19892 16040
rect 19352 16000 19892 16028
rect 19352 15960 19380 16000
rect 19886 15988 19892 16000
rect 19944 15988 19950 16040
rect 25041 16031 25099 16037
rect 25041 15997 25053 16031
rect 25087 15997 25099 16031
rect 25041 15991 25099 15997
rect 18340 15932 19380 15960
rect 25056 15960 25084 15991
rect 25866 15988 25872 16040
rect 25924 16028 25930 16040
rect 26344 16028 26372 16068
rect 27249 16065 27261 16068
rect 27295 16065 27307 16099
rect 27249 16059 27307 16065
rect 26970 16028 26976 16040
rect 25924 16000 26372 16028
rect 26931 16000 26976 16028
rect 25924 15988 25930 16000
rect 26970 15988 26976 16000
rect 27028 15988 27034 16040
rect 26050 15960 26056 15972
rect 25056 15932 26056 15960
rect 26050 15920 26056 15932
rect 26108 15920 26114 15972
rect 2685 15895 2743 15901
rect 2685 15861 2697 15895
rect 2731 15892 2743 15895
rect 4338 15892 4344 15904
rect 2731 15864 4344 15892
rect 2731 15861 2743 15864
rect 2685 15855 2743 15861
rect 4338 15852 4344 15864
rect 4396 15852 4402 15904
rect 12158 15852 12164 15904
rect 12216 15892 12222 15904
rect 12345 15895 12403 15901
rect 12345 15892 12357 15895
rect 12216 15864 12357 15892
rect 12216 15852 12222 15864
rect 12345 15861 12357 15864
rect 12391 15861 12403 15895
rect 12345 15855 12403 15861
rect 17405 15895 17463 15901
rect 17405 15861 17417 15895
rect 17451 15892 17463 15895
rect 17678 15892 17684 15904
rect 17451 15864 17684 15892
rect 17451 15861 17463 15864
rect 17405 15855 17463 15861
rect 17678 15852 17684 15864
rect 17736 15852 17742 15904
rect 25501 15895 25559 15901
rect 25501 15861 25513 15895
rect 25547 15892 25559 15895
rect 26142 15892 26148 15904
rect 25547 15864 26148 15892
rect 25547 15861 25559 15864
rect 25501 15855 25559 15861
rect 26142 15852 26148 15864
rect 26200 15852 26206 15904
rect 26602 15852 26608 15904
rect 26660 15892 26666 15904
rect 27157 15895 27215 15901
rect 27157 15892 27169 15895
rect 26660 15864 27169 15892
rect 26660 15852 26666 15864
rect 27157 15861 27169 15864
rect 27203 15861 27215 15895
rect 27982 15892 27988 15904
rect 27943 15864 27988 15892
rect 27157 15855 27215 15861
rect 27982 15852 27988 15864
rect 28040 15852 28046 15904
rect 1104 15802 28888 15824
rect 1104 15750 5582 15802
rect 5634 15750 5646 15802
rect 5698 15750 5710 15802
rect 5762 15750 5774 15802
rect 5826 15750 5838 15802
rect 5890 15750 14846 15802
rect 14898 15750 14910 15802
rect 14962 15750 14974 15802
rect 15026 15750 15038 15802
rect 15090 15750 15102 15802
rect 15154 15750 24110 15802
rect 24162 15750 24174 15802
rect 24226 15750 24238 15802
rect 24290 15750 24302 15802
rect 24354 15750 24366 15802
rect 24418 15750 28888 15802
rect 1104 15728 28888 15750
rect 14090 15648 14096 15700
rect 14148 15688 14154 15700
rect 15105 15691 15163 15697
rect 15105 15688 15117 15691
rect 14148 15660 15117 15688
rect 14148 15648 14154 15660
rect 15028 15632 15056 15660
rect 15105 15657 15117 15660
rect 15151 15657 15163 15691
rect 15105 15651 15163 15657
rect 17957 15691 18015 15697
rect 17957 15657 17969 15691
rect 18003 15688 18015 15691
rect 18690 15688 18696 15700
rect 18003 15660 18696 15688
rect 18003 15657 18015 15660
rect 17957 15651 18015 15657
rect 18690 15648 18696 15660
rect 18748 15648 18754 15700
rect 19242 15688 19248 15700
rect 19203 15660 19248 15688
rect 19242 15648 19248 15660
rect 19300 15648 19306 15700
rect 19705 15691 19763 15697
rect 19705 15688 19717 15691
rect 19352 15660 19717 15688
rect 13354 15580 13360 15632
rect 13412 15620 13418 15632
rect 14182 15620 14188 15632
rect 13412 15592 14188 15620
rect 13412 15580 13418 15592
rect 14182 15580 14188 15592
rect 14240 15580 14246 15632
rect 15010 15580 15016 15632
rect 15068 15580 15074 15632
rect 17405 15623 17463 15629
rect 17405 15589 17417 15623
rect 17451 15620 17463 15623
rect 17678 15620 17684 15632
rect 17451 15592 17684 15620
rect 17451 15589 17463 15592
rect 17405 15583 17463 15589
rect 17678 15580 17684 15592
rect 17736 15580 17742 15632
rect 19150 15620 19156 15632
rect 18432 15592 19156 15620
rect 11977 15555 12035 15561
rect 11977 15521 11989 15555
rect 12023 15552 12035 15555
rect 12434 15552 12440 15564
rect 12023 15524 12440 15552
rect 12023 15521 12035 15524
rect 11977 15515 12035 15521
rect 12434 15512 12440 15524
rect 12492 15512 12498 15564
rect 14093 15555 14151 15561
rect 14093 15521 14105 15555
rect 14139 15552 14151 15555
rect 14366 15552 14372 15564
rect 14139 15524 14372 15552
rect 14139 15521 14151 15524
rect 14093 15515 14151 15521
rect 14366 15512 14372 15524
rect 14424 15512 14430 15564
rect 16206 15512 16212 15564
rect 16264 15552 16270 15564
rect 17037 15555 17095 15561
rect 17037 15552 17049 15555
rect 16264 15524 17049 15552
rect 16264 15512 16270 15524
rect 17037 15521 17049 15524
rect 17083 15521 17095 15555
rect 17037 15515 17095 15521
rect 17497 15555 17555 15561
rect 17497 15521 17509 15555
rect 17543 15552 17555 15555
rect 18233 15555 18291 15561
rect 18233 15552 18245 15555
rect 17543 15524 18245 15552
rect 17543 15521 17555 15524
rect 17497 15515 17555 15521
rect 18233 15521 18245 15524
rect 18279 15521 18291 15555
rect 18233 15515 18291 15521
rect 18432 15496 18460 15592
rect 19150 15580 19156 15592
rect 19208 15580 19214 15632
rect 19352 15552 19380 15660
rect 19705 15657 19717 15660
rect 19751 15657 19763 15691
rect 20714 15688 20720 15700
rect 20675 15660 20720 15688
rect 19705 15651 19763 15657
rect 18708 15524 19380 15552
rect 19720 15552 19748 15651
rect 20714 15648 20720 15660
rect 20772 15648 20778 15700
rect 24578 15648 24584 15700
rect 24636 15688 24642 15700
rect 25225 15691 25283 15697
rect 25225 15688 25237 15691
rect 24636 15660 25237 15688
rect 24636 15648 24642 15660
rect 25225 15657 25237 15660
rect 25271 15657 25283 15691
rect 27982 15688 27988 15700
rect 25225 15651 25283 15657
rect 25332 15660 27988 15688
rect 20622 15580 20628 15632
rect 20680 15620 20686 15632
rect 25332 15620 25360 15660
rect 27982 15648 27988 15660
rect 28040 15648 28046 15700
rect 20680 15592 25360 15620
rect 20680 15580 20686 15592
rect 22649 15555 22707 15561
rect 19720 15524 20300 15552
rect 1394 15444 1400 15496
rect 1452 15484 1458 15496
rect 1489 15487 1547 15493
rect 1489 15484 1501 15487
rect 1452 15456 1501 15484
rect 1452 15444 1458 15456
rect 1489 15453 1501 15456
rect 1535 15453 1547 15487
rect 3970 15484 3976 15496
rect 3931 15456 3976 15484
rect 1489 15447 1547 15453
rect 3970 15444 3976 15456
rect 4028 15444 4034 15496
rect 12158 15484 12164 15496
rect 12119 15456 12164 15484
rect 12158 15444 12164 15456
rect 12216 15444 12222 15496
rect 12345 15487 12403 15493
rect 12345 15453 12357 15487
rect 12391 15484 12403 15487
rect 12989 15487 13047 15493
rect 12989 15484 13001 15487
rect 12391 15456 13001 15484
rect 12391 15453 12403 15456
rect 12345 15447 12403 15453
rect 12989 15453 13001 15456
rect 13035 15453 13047 15487
rect 15013 15487 15071 15493
rect 15013 15484 15025 15487
rect 12989 15447 13047 15453
rect 14568 15456 15025 15484
rect 14568 15428 14596 15456
rect 15013 15453 15025 15456
rect 15059 15453 15071 15487
rect 15013 15447 15071 15453
rect 15378 15444 15384 15496
rect 15436 15484 15442 15496
rect 15657 15487 15715 15493
rect 15657 15484 15669 15487
rect 15436 15456 15669 15484
rect 15436 15444 15442 15456
rect 15657 15453 15669 15456
rect 15703 15453 15715 15487
rect 15657 15447 15715 15453
rect 15746 15444 15752 15496
rect 15804 15484 15810 15496
rect 15841 15487 15899 15493
rect 15841 15484 15853 15487
rect 15804 15456 15853 15484
rect 15804 15444 15810 15456
rect 15841 15453 15853 15456
rect 15887 15453 15899 15487
rect 18322 15484 18328 15496
rect 18283 15456 18328 15484
rect 15841 15447 15899 15453
rect 18322 15444 18328 15456
rect 18380 15444 18386 15496
rect 18414 15444 18420 15496
rect 18472 15484 18478 15496
rect 18708 15493 18736 15524
rect 18693 15487 18751 15493
rect 18693 15484 18705 15487
rect 18472 15456 18517 15484
rect 18616 15456 18705 15484
rect 18472 15444 18478 15456
rect 14550 15416 14556 15428
rect 14511 15388 14556 15416
rect 14550 15376 14556 15388
rect 14608 15376 14614 15428
rect 16298 15376 16304 15428
rect 16356 15416 16362 15428
rect 18616 15416 18644 15456
rect 18693 15453 18705 15456
rect 18739 15453 18751 15487
rect 19426 15484 19432 15496
rect 19387 15456 19432 15484
rect 18693 15447 18751 15453
rect 19426 15444 19432 15456
rect 19484 15444 19490 15496
rect 19518 15444 19524 15496
rect 19576 15484 19582 15496
rect 20272 15493 20300 15524
rect 22649 15521 22661 15555
rect 22695 15521 22707 15555
rect 22830 15552 22836 15564
rect 22791 15524 22836 15552
rect 22649 15515 22707 15521
rect 19797 15487 19855 15493
rect 19576 15456 19621 15484
rect 19576 15444 19582 15456
rect 19797 15453 19809 15487
rect 19843 15453 19855 15487
rect 19797 15447 19855 15453
rect 20257 15487 20315 15493
rect 20257 15453 20269 15487
rect 20303 15453 20315 15487
rect 20533 15487 20591 15493
rect 20533 15484 20545 15487
rect 20257 15447 20315 15453
rect 20456 15456 20545 15484
rect 19812 15416 19840 15447
rect 20349 15419 20407 15425
rect 20349 15416 20361 15419
rect 16356 15388 18644 15416
rect 18708 15388 20361 15416
rect 16356 15376 16362 15388
rect 18708 15360 18736 15388
rect 20349 15385 20361 15388
rect 20395 15385 20407 15419
rect 20349 15379 20407 15385
rect 3881 15351 3939 15357
rect 3881 15317 3893 15351
rect 3927 15348 3939 15351
rect 4154 15348 4160 15360
rect 3927 15320 4160 15348
rect 3927 15317 3939 15320
rect 3881 15311 3939 15317
rect 4154 15308 4160 15320
rect 4212 15308 4218 15360
rect 12802 15348 12808 15360
rect 12763 15320 12808 15348
rect 12802 15308 12808 15320
rect 12860 15308 12866 15360
rect 15470 15308 15476 15360
rect 15528 15348 15534 15360
rect 15657 15351 15715 15357
rect 15657 15348 15669 15351
rect 15528 15320 15669 15348
rect 15528 15308 15534 15320
rect 15657 15317 15669 15320
rect 15703 15317 15715 15351
rect 15657 15311 15715 15317
rect 18601 15351 18659 15357
rect 18601 15317 18613 15351
rect 18647 15348 18659 15351
rect 18690 15348 18696 15360
rect 18647 15320 18696 15348
rect 18647 15317 18659 15320
rect 18601 15311 18659 15317
rect 18690 15308 18696 15320
rect 18748 15308 18754 15360
rect 19150 15308 19156 15360
rect 19208 15348 19214 15360
rect 20456 15348 20484 15456
rect 20533 15453 20545 15456
rect 20579 15453 20591 15487
rect 22664 15484 22692 15515
rect 22830 15512 22836 15524
rect 22888 15512 22894 15564
rect 25682 15512 25688 15564
rect 25740 15552 25746 15564
rect 25869 15555 25927 15561
rect 25869 15552 25881 15555
rect 25740 15524 25881 15552
rect 25740 15512 25746 15524
rect 25869 15521 25881 15524
rect 25915 15521 25927 15555
rect 25869 15515 25927 15521
rect 26050 15512 26056 15564
rect 26108 15552 26114 15564
rect 26329 15555 26387 15561
rect 26329 15552 26341 15555
rect 26108 15524 26341 15552
rect 26108 15512 26114 15524
rect 26329 15521 26341 15524
rect 26375 15521 26387 15555
rect 28166 15552 28172 15564
rect 28127 15524 28172 15552
rect 26329 15515 26387 15521
rect 28166 15512 28172 15524
rect 28224 15512 28230 15564
rect 23566 15484 23572 15496
rect 22664 15456 23572 15484
rect 20533 15447 20591 15453
rect 23566 15444 23572 15456
rect 23624 15444 23630 15496
rect 24765 15487 24823 15493
rect 24765 15453 24777 15487
rect 24811 15484 24823 15487
rect 24854 15484 24860 15496
rect 24811 15456 24860 15484
rect 24811 15453 24823 15456
rect 24765 15447 24823 15453
rect 24854 15444 24860 15456
rect 24912 15444 24918 15496
rect 25409 15487 25467 15493
rect 25409 15453 25421 15487
rect 25455 15484 25467 15487
rect 25455 15456 26372 15484
rect 25455 15453 25467 15456
rect 25409 15447 25467 15453
rect 26344 15428 26372 15456
rect 22925 15419 22983 15425
rect 22925 15385 22937 15419
rect 22971 15416 22983 15419
rect 24118 15416 24124 15428
rect 22971 15388 24124 15416
rect 22971 15385 22983 15388
rect 22925 15379 22983 15385
rect 24118 15376 24124 15388
rect 24176 15376 24182 15428
rect 25314 15376 25320 15428
rect 25372 15416 25378 15428
rect 25501 15419 25559 15425
rect 25501 15416 25513 15419
rect 25372 15388 25513 15416
rect 25372 15376 25378 15388
rect 25501 15385 25513 15388
rect 25547 15385 25559 15419
rect 25501 15379 25559 15385
rect 25593 15419 25651 15425
rect 25593 15385 25605 15419
rect 25639 15385 25651 15419
rect 25593 15379 25651 15385
rect 25731 15419 25789 15425
rect 25731 15385 25743 15419
rect 25777 15416 25789 15419
rect 25777 15388 26188 15416
rect 25777 15385 25789 15388
rect 25731 15379 25789 15385
rect 19208 15320 20484 15348
rect 19208 15308 19214 15320
rect 23014 15308 23020 15360
rect 23072 15348 23078 15360
rect 23293 15351 23351 15357
rect 23293 15348 23305 15351
rect 23072 15320 23305 15348
rect 23072 15308 23078 15320
rect 23293 15317 23305 15320
rect 23339 15317 23351 15351
rect 23293 15311 23351 15317
rect 23658 15308 23664 15360
rect 23716 15348 23722 15360
rect 24581 15351 24639 15357
rect 24581 15348 24593 15351
rect 23716 15320 24593 15348
rect 23716 15308 23722 15320
rect 24581 15317 24593 15320
rect 24627 15317 24639 15351
rect 25608 15348 25636 15379
rect 25866 15348 25872 15360
rect 25608 15320 25872 15348
rect 24581 15311 24639 15317
rect 25866 15308 25872 15320
rect 25924 15308 25930 15360
rect 26160 15348 26188 15388
rect 26326 15376 26332 15428
rect 26384 15376 26390 15428
rect 26510 15416 26516 15428
rect 26471 15388 26516 15416
rect 26510 15376 26516 15388
rect 26568 15376 26574 15428
rect 26418 15348 26424 15360
rect 26160 15320 26424 15348
rect 26418 15308 26424 15320
rect 26476 15308 26482 15360
rect 1104 15258 28888 15280
rect 1104 15206 10214 15258
rect 10266 15206 10278 15258
rect 10330 15206 10342 15258
rect 10394 15206 10406 15258
rect 10458 15206 10470 15258
rect 10522 15206 19478 15258
rect 19530 15206 19542 15258
rect 19594 15206 19606 15258
rect 19658 15206 19670 15258
rect 19722 15206 19734 15258
rect 19786 15206 28888 15258
rect 1104 15184 28888 15206
rect 4062 15144 4068 15156
rect 2148 15116 4068 15144
rect 2148 15020 2176 15116
rect 4062 15104 4068 15116
rect 4120 15104 4126 15156
rect 13354 15144 13360 15156
rect 13315 15116 13360 15144
rect 13354 15104 13360 15116
rect 13412 15104 13418 15156
rect 18322 15104 18328 15156
rect 18380 15144 18386 15156
rect 18877 15147 18935 15153
rect 18877 15144 18889 15147
rect 18380 15116 18889 15144
rect 18380 15104 18386 15116
rect 18877 15113 18889 15116
rect 18923 15113 18935 15147
rect 18877 15107 18935 15113
rect 20625 15147 20683 15153
rect 20625 15113 20637 15147
rect 20671 15144 20683 15147
rect 23658 15144 23664 15156
rect 20671 15116 23664 15144
rect 20671 15113 20683 15116
rect 20625 15107 20683 15113
rect 23658 15104 23664 15116
rect 23716 15104 23722 15156
rect 24118 15144 24124 15156
rect 24079 15116 24124 15144
rect 24118 15104 24124 15116
rect 24176 15144 24182 15156
rect 24762 15144 24768 15156
rect 24176 15116 24768 15144
rect 24176 15104 24182 15116
rect 24762 15104 24768 15116
rect 24820 15104 24826 15156
rect 26234 15104 26240 15156
rect 26292 15144 26298 15156
rect 26329 15147 26387 15153
rect 26329 15144 26341 15147
rect 26292 15116 26341 15144
rect 26292 15104 26298 15116
rect 26329 15113 26341 15116
rect 26375 15113 26387 15147
rect 26329 15107 26387 15113
rect 26510 15104 26516 15156
rect 26568 15144 26574 15156
rect 28077 15147 28135 15153
rect 28077 15144 28089 15147
rect 26568 15116 28089 15144
rect 26568 15104 26574 15116
rect 28077 15113 28089 15116
rect 28123 15113 28135 15147
rect 28077 15107 28135 15113
rect 4154 15076 4160 15088
rect 4115 15048 4160 15076
rect 4154 15036 4160 15048
rect 4212 15036 4218 15088
rect 12244 15079 12302 15085
rect 12244 15045 12256 15079
rect 12290 15076 12302 15079
rect 12802 15076 12808 15088
rect 12290 15048 12808 15076
rect 12290 15045 12302 15048
rect 12244 15039 12302 15045
rect 12802 15036 12808 15048
rect 12860 15036 12866 15088
rect 19337 15079 19395 15085
rect 19337 15045 19349 15079
rect 19383 15076 19395 15079
rect 19978 15076 19984 15088
rect 19383 15048 19984 15076
rect 19383 15045 19395 15048
rect 19337 15039 19395 15045
rect 19978 15036 19984 15048
rect 20036 15036 20042 15088
rect 22278 15036 22284 15088
rect 22336 15076 22342 15088
rect 22986 15079 23044 15085
rect 22986 15076 22998 15079
rect 22336 15048 22998 15076
rect 22336 15036 22342 15048
rect 22986 15045 22998 15048
rect 23032 15045 23044 15079
rect 22986 15039 23044 15045
rect 25314 15036 25320 15088
rect 25372 15076 25378 15088
rect 25590 15076 25596 15088
rect 25372 15048 25596 15076
rect 25372 15036 25378 15048
rect 25590 15036 25596 15048
rect 25648 15076 25654 15088
rect 25648 15048 27384 15076
rect 25648 15036 25654 15048
rect 1949 15011 2007 15017
rect 1949 14977 1961 15011
rect 1995 15008 2007 15011
rect 2130 15008 2136 15020
rect 1995 14980 2136 15008
rect 1995 14977 2007 14980
rect 1949 14971 2007 14977
rect 2130 14968 2136 14980
rect 2188 14968 2194 15020
rect 4338 14968 4344 15020
rect 4396 15008 4402 15020
rect 4396 14980 4441 15008
rect 4396 14968 4402 14980
rect 11882 14968 11888 15020
rect 11940 15008 11946 15020
rect 11977 15011 12035 15017
rect 11977 15008 11989 15011
rect 11940 14980 11989 15008
rect 11940 14968 11946 14980
rect 11977 14977 11989 14980
rect 12023 14977 12035 15011
rect 15010 15008 15016 15020
rect 14971 14980 15016 15008
rect 11977 14971 12035 14977
rect 15010 14968 15016 14980
rect 15068 14968 15074 15020
rect 15197 15011 15255 15017
rect 15197 14977 15209 15011
rect 15243 15008 15255 15011
rect 15286 15008 15292 15020
rect 15243 14980 15292 15008
rect 15243 14977 15255 14980
rect 15197 14971 15255 14977
rect 15286 14968 15292 14980
rect 15344 14968 15350 15020
rect 20530 15008 20536 15020
rect 20491 14980 20536 15008
rect 20530 14968 20536 14980
rect 20588 14968 20594 15020
rect 22094 14968 22100 15020
rect 22152 15008 22158 15020
rect 26237 15011 26295 15017
rect 22152 14980 22197 15008
rect 22152 14968 22158 14980
rect 26237 14977 26249 15011
rect 26283 14977 26295 15011
rect 26418 15008 26424 15020
rect 26379 14980 26424 15008
rect 26237 14971 26295 14977
rect 2774 14940 2780 14952
rect 2735 14912 2780 14940
rect 2774 14900 2780 14912
rect 2832 14900 2838 14952
rect 16482 14900 16488 14952
rect 16540 14940 16546 14952
rect 20254 14940 20260 14952
rect 16540 14912 20260 14940
rect 16540 14900 16546 14912
rect 20254 14900 20260 14912
rect 20312 14940 20318 14952
rect 20717 14943 20775 14949
rect 20717 14940 20729 14943
rect 20312 14912 20729 14940
rect 20312 14900 20318 14912
rect 20717 14909 20729 14912
rect 20763 14909 20775 14943
rect 20717 14903 20775 14909
rect 21818 14900 21824 14952
rect 21876 14940 21882 14952
rect 22741 14943 22799 14949
rect 22741 14940 22753 14943
rect 21876 14912 22753 14940
rect 21876 14900 21882 14912
rect 22741 14909 22753 14912
rect 22787 14909 22799 14943
rect 22741 14903 22799 14909
rect 24949 14943 25007 14949
rect 24949 14909 24961 14943
rect 24995 14940 25007 14943
rect 25130 14940 25136 14952
rect 24995 14912 25136 14940
rect 24995 14909 25007 14912
rect 24949 14903 25007 14909
rect 25130 14900 25136 14912
rect 25188 14900 25194 14952
rect 25225 14943 25283 14949
rect 25225 14909 25237 14943
rect 25271 14940 25283 14943
rect 25774 14940 25780 14952
rect 25271 14912 25780 14940
rect 25271 14909 25283 14912
rect 25225 14903 25283 14909
rect 25774 14900 25780 14912
rect 25832 14940 25838 14952
rect 26252 14940 26280 14971
rect 26418 14968 26424 14980
rect 26476 14968 26482 15020
rect 27356 15017 27384 15048
rect 27341 15011 27399 15017
rect 27341 14977 27353 15011
rect 27387 14977 27399 15011
rect 27341 14971 27399 14977
rect 27985 15011 28043 15017
rect 27985 14977 27997 15011
rect 28031 14977 28043 15011
rect 27985 14971 28043 14977
rect 25832 14912 26280 14940
rect 25832 14900 25838 14912
rect 19061 14875 19119 14881
rect 19061 14841 19073 14875
rect 19107 14872 19119 14875
rect 20530 14872 20536 14884
rect 19107 14844 20536 14872
rect 19107 14841 19119 14844
rect 19061 14835 19119 14841
rect 19352 14816 19380 14844
rect 20530 14832 20536 14844
rect 20588 14832 20594 14884
rect 22278 14872 22284 14884
rect 22239 14844 22284 14872
rect 22278 14832 22284 14844
rect 22336 14832 22342 14884
rect 26252 14872 26280 14912
rect 26326 14900 26332 14952
rect 26384 14940 26390 14952
rect 27157 14943 27215 14949
rect 27157 14940 27169 14943
rect 26384 14912 27169 14940
rect 26384 14900 26390 14912
rect 27157 14909 27169 14912
rect 27203 14909 27215 14943
rect 27157 14903 27215 14909
rect 27246 14900 27252 14952
rect 27304 14940 27310 14952
rect 27304 14912 27349 14940
rect 27304 14900 27310 14912
rect 27430 14900 27436 14952
rect 27488 14940 27494 14952
rect 27488 14912 27533 14940
rect 27488 14900 27494 14912
rect 26878 14872 26884 14884
rect 26252 14844 26884 14872
rect 26878 14832 26884 14844
rect 26936 14832 26942 14884
rect 27522 14872 27528 14884
rect 27356 14844 27528 14872
rect 27356 14816 27384 14844
rect 27522 14832 27528 14844
rect 27580 14872 27586 14884
rect 28000 14872 28028 14971
rect 27580 14844 28028 14872
rect 27580 14832 27586 14844
rect 1578 14764 1584 14816
rect 1636 14804 1642 14816
rect 1857 14807 1915 14813
rect 1857 14804 1869 14807
rect 1636 14776 1869 14804
rect 1636 14764 1642 14776
rect 1857 14773 1869 14776
rect 1903 14773 1915 14807
rect 1857 14767 1915 14773
rect 15105 14807 15163 14813
rect 15105 14773 15117 14807
rect 15151 14804 15163 14807
rect 15194 14804 15200 14816
rect 15151 14776 15200 14804
rect 15151 14773 15163 14776
rect 15105 14767 15163 14773
rect 15194 14764 15200 14776
rect 15252 14764 15258 14816
rect 19334 14764 19340 14816
rect 19392 14764 19398 14816
rect 19978 14764 19984 14816
rect 20036 14804 20042 14816
rect 20165 14807 20223 14813
rect 20165 14804 20177 14807
rect 20036 14776 20177 14804
rect 20036 14764 20042 14776
rect 20165 14773 20177 14776
rect 20211 14773 20223 14807
rect 20165 14767 20223 14773
rect 24854 14764 24860 14816
rect 24912 14804 24918 14816
rect 25222 14804 25228 14816
rect 24912 14776 25228 14804
rect 24912 14764 24918 14776
rect 25222 14764 25228 14776
rect 25280 14764 25286 14816
rect 26510 14764 26516 14816
rect 26568 14804 26574 14816
rect 26973 14807 27031 14813
rect 26973 14804 26985 14807
rect 26568 14776 26985 14804
rect 26568 14764 26574 14776
rect 26973 14773 26985 14776
rect 27019 14773 27031 14807
rect 26973 14767 27031 14773
rect 27338 14764 27344 14816
rect 27396 14764 27402 14816
rect 1104 14714 28888 14736
rect 1104 14662 5582 14714
rect 5634 14662 5646 14714
rect 5698 14662 5710 14714
rect 5762 14662 5774 14714
rect 5826 14662 5838 14714
rect 5890 14662 14846 14714
rect 14898 14662 14910 14714
rect 14962 14662 14974 14714
rect 15026 14662 15038 14714
rect 15090 14662 15102 14714
rect 15154 14662 24110 14714
rect 24162 14662 24174 14714
rect 24226 14662 24238 14714
rect 24290 14662 24302 14714
rect 24354 14662 24366 14714
rect 24418 14662 28888 14714
rect 1104 14640 28888 14662
rect 15289 14603 15347 14609
rect 15289 14569 15301 14603
rect 15335 14600 15347 14603
rect 15470 14600 15476 14612
rect 15335 14572 15476 14600
rect 15335 14569 15347 14572
rect 15289 14563 15347 14569
rect 15470 14560 15476 14572
rect 15528 14560 15534 14612
rect 16025 14603 16083 14609
rect 16025 14569 16037 14603
rect 16071 14600 16083 14603
rect 16850 14600 16856 14612
rect 16071 14572 16856 14600
rect 16071 14569 16083 14572
rect 16025 14563 16083 14569
rect 16850 14560 16856 14572
rect 16908 14560 16914 14612
rect 22094 14560 22100 14612
rect 22152 14600 22158 14612
rect 22833 14603 22891 14609
rect 22833 14600 22845 14603
rect 22152 14572 22845 14600
rect 22152 14560 22158 14572
rect 22833 14569 22845 14572
rect 22879 14569 22891 14603
rect 25130 14600 25136 14612
rect 25091 14572 25136 14600
rect 22833 14563 22891 14569
rect 25130 14560 25136 14572
rect 25188 14560 25194 14612
rect 25869 14603 25927 14609
rect 25869 14569 25881 14603
rect 25915 14600 25927 14603
rect 27430 14600 27436 14612
rect 25915 14572 27436 14600
rect 25915 14569 25927 14572
rect 25869 14563 25927 14569
rect 27430 14560 27436 14572
rect 27488 14560 27494 14612
rect 22373 14535 22431 14541
rect 22373 14501 22385 14535
rect 22419 14532 22431 14535
rect 22738 14532 22744 14544
rect 22419 14504 22744 14532
rect 22419 14501 22431 14504
rect 22373 14495 22431 14501
rect 22738 14492 22744 14504
rect 22796 14492 22802 14544
rect 24946 14532 24952 14544
rect 24504 14504 24952 14532
rect 24504 14476 24532 14504
rect 24946 14492 24952 14504
rect 25004 14492 25010 14544
rect 1394 14464 1400 14476
rect 1355 14436 1400 14464
rect 1394 14424 1400 14436
rect 1452 14424 1458 14476
rect 1578 14464 1584 14476
rect 1539 14436 1584 14464
rect 1578 14424 1584 14436
rect 1636 14424 1642 14476
rect 1854 14464 1860 14476
rect 1815 14436 1860 14464
rect 1854 14424 1860 14436
rect 1912 14424 1918 14476
rect 19334 14424 19340 14476
rect 19392 14464 19398 14476
rect 19797 14467 19855 14473
rect 19797 14464 19809 14467
rect 19392 14436 19809 14464
rect 19392 14424 19398 14436
rect 19797 14433 19809 14436
rect 19843 14464 19855 14467
rect 20806 14464 20812 14476
rect 19843 14436 20812 14464
rect 19843 14433 19855 14436
rect 19797 14427 19855 14433
rect 20806 14424 20812 14436
rect 20864 14424 20870 14476
rect 24486 14464 24492 14476
rect 24447 14436 24492 14464
rect 24486 14424 24492 14436
rect 24544 14424 24550 14476
rect 24670 14464 24676 14476
rect 24631 14436 24676 14464
rect 24670 14424 24676 14436
rect 24728 14424 24734 14476
rect 27522 14464 27528 14476
rect 27483 14436 27528 14464
rect 27522 14424 27528 14436
rect 27580 14424 27586 14476
rect 15562 14356 15568 14408
rect 15620 14396 15626 14408
rect 15933 14399 15991 14405
rect 15933 14396 15945 14399
rect 15620 14368 15945 14396
rect 15620 14356 15626 14368
rect 15933 14365 15945 14368
rect 15979 14396 15991 14399
rect 16114 14396 16120 14408
rect 15979 14368 16120 14396
rect 15979 14365 15991 14368
rect 15933 14359 15991 14365
rect 16114 14356 16120 14368
rect 16172 14356 16178 14408
rect 19978 14396 19984 14408
rect 19939 14368 19984 14396
rect 19978 14356 19984 14368
rect 20036 14356 20042 14408
rect 20990 14396 20996 14408
rect 20903 14368 20996 14396
rect 20990 14356 20996 14368
rect 21048 14396 21054 14408
rect 21818 14396 21824 14408
rect 21048 14368 21824 14396
rect 21048 14356 21054 14368
rect 21818 14356 21824 14368
rect 21876 14356 21882 14408
rect 23014 14396 23020 14408
rect 22975 14368 23020 14396
rect 23014 14356 23020 14368
rect 23072 14356 23078 14408
rect 23201 14399 23259 14405
rect 23201 14365 23213 14399
rect 23247 14396 23259 14399
rect 23382 14396 23388 14408
rect 23247 14368 23388 14396
rect 23247 14365 23259 14368
rect 23201 14359 23259 14365
rect 23382 14356 23388 14368
rect 23440 14356 23446 14408
rect 24762 14396 24768 14408
rect 24723 14368 24768 14396
rect 24762 14356 24768 14368
rect 24820 14356 24826 14408
rect 25590 14396 25596 14408
rect 25551 14368 25596 14396
rect 25590 14356 25596 14368
rect 25648 14356 25654 14408
rect 25866 14396 25872 14408
rect 25827 14368 25872 14396
rect 25866 14356 25872 14368
rect 25924 14356 25930 14408
rect 28166 14356 28172 14408
rect 28224 14396 28230 14408
rect 28224 14368 28269 14396
rect 28224 14356 28230 14368
rect 15194 14288 15200 14340
rect 15252 14337 15258 14340
rect 15252 14331 15315 14337
rect 15252 14297 15269 14331
rect 15303 14297 15315 14331
rect 15252 14291 15315 14297
rect 15252 14288 15258 14291
rect 15378 14288 15384 14340
rect 15436 14328 15442 14340
rect 15473 14331 15531 14337
rect 15473 14328 15485 14331
rect 15436 14300 15485 14328
rect 15436 14288 15442 14300
rect 15473 14297 15485 14300
rect 15519 14328 15531 14331
rect 16666 14328 16672 14340
rect 15519 14300 16672 14328
rect 15519 14297 15531 14300
rect 15473 14291 15531 14297
rect 16666 14288 16672 14300
rect 16724 14288 16730 14340
rect 21266 14337 21272 14340
rect 21260 14328 21272 14337
rect 21227 14300 21272 14328
rect 21260 14291 21272 14300
rect 21266 14288 21272 14291
rect 21324 14288 21330 14340
rect 27890 14288 27896 14340
rect 27948 14328 27954 14340
rect 27985 14331 28043 14337
rect 27985 14328 27997 14331
rect 27948 14300 27997 14328
rect 27948 14288 27954 14300
rect 27985 14297 27997 14300
rect 28031 14297 28043 14331
rect 27985 14291 28043 14297
rect 14274 14220 14280 14272
rect 14332 14260 14338 14272
rect 15105 14263 15163 14269
rect 15105 14260 15117 14263
rect 14332 14232 15117 14260
rect 14332 14220 14338 14232
rect 15105 14229 15117 14232
rect 15151 14229 15163 14263
rect 15105 14223 15163 14229
rect 20070 14220 20076 14272
rect 20128 14260 20134 14272
rect 20165 14263 20223 14269
rect 20165 14260 20177 14263
rect 20128 14232 20177 14260
rect 20128 14220 20134 14232
rect 20165 14229 20177 14232
rect 20211 14229 20223 14263
rect 20165 14223 20223 14229
rect 25685 14263 25743 14269
rect 25685 14229 25697 14263
rect 25731 14260 25743 14263
rect 25774 14260 25780 14272
rect 25731 14232 25780 14260
rect 25731 14229 25743 14232
rect 25685 14223 25743 14229
rect 25774 14220 25780 14232
rect 25832 14260 25838 14272
rect 26602 14260 26608 14272
rect 25832 14232 26608 14260
rect 25832 14220 25838 14232
rect 26602 14220 26608 14232
rect 26660 14220 26666 14272
rect 1104 14170 28888 14192
rect 1104 14118 10214 14170
rect 10266 14118 10278 14170
rect 10330 14118 10342 14170
rect 10394 14118 10406 14170
rect 10458 14118 10470 14170
rect 10522 14118 19478 14170
rect 19530 14118 19542 14170
rect 19594 14118 19606 14170
rect 19658 14118 19670 14170
rect 19722 14118 19734 14170
rect 19786 14118 28888 14170
rect 1104 14096 28888 14118
rect 16666 14016 16672 14068
rect 16724 14056 16730 14068
rect 17247 14059 17305 14065
rect 16724 14028 17080 14056
rect 16724 14016 16730 14028
rect 14734 13988 14740 14000
rect 13372 13960 14740 13988
rect 11882 13880 11888 13932
rect 11940 13920 11946 13932
rect 13372 13929 13400 13960
rect 14734 13948 14740 13960
rect 14792 13948 14798 14000
rect 15565 13991 15623 13997
rect 15565 13957 15577 13991
rect 15611 13988 15623 13991
rect 16850 13988 16856 14000
rect 15611 13960 16856 13988
rect 15611 13957 15623 13960
rect 15565 13951 15623 13957
rect 16850 13948 16856 13960
rect 16908 13948 16914 14000
rect 17052 13997 17080 14028
rect 17247 14025 17259 14059
rect 17293 14056 17305 14059
rect 17862 14056 17868 14068
rect 17293 14028 17868 14056
rect 17293 14025 17305 14028
rect 17247 14019 17305 14025
rect 17862 14016 17868 14028
rect 17920 14056 17926 14068
rect 17957 14059 18015 14065
rect 17957 14056 17969 14059
rect 17920 14028 17969 14056
rect 17920 14016 17926 14028
rect 17957 14025 17969 14028
rect 18003 14025 18015 14059
rect 18690 14056 18696 14068
rect 18651 14028 18696 14056
rect 17957 14019 18015 14025
rect 18690 14016 18696 14028
rect 18748 14016 18754 14068
rect 20530 14016 20536 14068
rect 20588 14056 20594 14068
rect 20901 14059 20959 14065
rect 20901 14056 20913 14059
rect 20588 14028 20913 14056
rect 20588 14016 20594 14028
rect 20901 14025 20913 14028
rect 20947 14025 20959 14059
rect 20901 14019 20959 14025
rect 25130 14016 25136 14068
rect 25188 14016 25194 14068
rect 25317 14059 25375 14065
rect 25317 14025 25329 14059
rect 25363 14056 25375 14059
rect 25590 14056 25596 14068
rect 25363 14028 25596 14056
rect 25363 14025 25375 14028
rect 25317 14019 25375 14025
rect 25590 14016 25596 14028
rect 25648 14016 25654 14068
rect 27890 14056 27896 14068
rect 27851 14028 27896 14056
rect 27890 14016 27896 14028
rect 27948 14016 27954 14068
rect 17037 13991 17095 13997
rect 17037 13957 17049 13991
rect 17083 13957 17095 13991
rect 20990 13988 20996 14000
rect 17037 13951 17095 13957
rect 19536 13960 20996 13988
rect 13357 13923 13415 13929
rect 13357 13920 13369 13923
rect 11940 13892 13369 13920
rect 11940 13880 11946 13892
rect 13357 13889 13369 13892
rect 13403 13889 13415 13923
rect 13357 13883 13415 13889
rect 13624 13923 13682 13929
rect 13624 13889 13636 13923
rect 13670 13920 13682 13923
rect 14090 13920 14096 13932
rect 13670 13892 14096 13920
rect 13670 13889 13682 13892
rect 13624 13883 13682 13889
rect 14090 13880 14096 13892
rect 14148 13880 14154 13932
rect 15381 13923 15439 13929
rect 15381 13889 15393 13923
rect 15427 13920 15439 13923
rect 15470 13920 15476 13932
rect 15427 13892 15476 13920
rect 15427 13889 15439 13892
rect 15381 13883 15439 13889
rect 15470 13880 15476 13892
rect 15528 13880 15534 13932
rect 17770 13880 17776 13932
rect 17828 13920 17834 13932
rect 17865 13923 17923 13929
rect 17865 13920 17877 13923
rect 17828 13892 17877 13920
rect 17828 13880 17834 13892
rect 17865 13889 17877 13892
rect 17911 13889 17923 13923
rect 17865 13883 17923 13889
rect 18049 13923 18107 13929
rect 18049 13889 18061 13923
rect 18095 13920 18107 13923
rect 18322 13920 18328 13932
rect 18095 13892 18328 13920
rect 18095 13889 18107 13892
rect 18049 13883 18107 13889
rect 18322 13880 18328 13892
rect 18380 13920 18386 13932
rect 19536 13929 19564 13960
rect 20990 13948 20996 13960
rect 21048 13948 21054 14000
rect 24949 13991 25007 13997
rect 24949 13957 24961 13991
rect 24995 13988 25007 13991
rect 25148 13988 25176 14016
rect 24995 13960 25176 13988
rect 24995 13957 25007 13960
rect 24949 13951 25007 13957
rect 25866 13948 25872 14000
rect 25924 13988 25930 14000
rect 26973 13991 27031 13997
rect 26973 13988 26985 13991
rect 25924 13960 26985 13988
rect 25924 13948 25930 13960
rect 26973 13957 26985 13960
rect 27019 13957 27031 13991
rect 26973 13951 27031 13957
rect 27246 13948 27252 14000
rect 27304 13988 27310 14000
rect 27341 13991 27399 13997
rect 27341 13988 27353 13991
rect 27304 13960 27353 13988
rect 27304 13948 27310 13960
rect 27341 13957 27353 13960
rect 27387 13957 27399 13991
rect 27341 13951 27399 13957
rect 19794 13929 19800 13932
rect 18601 13923 18659 13929
rect 18601 13920 18613 13923
rect 18380 13892 18613 13920
rect 18380 13880 18386 13892
rect 18601 13889 18613 13892
rect 18647 13889 18659 13923
rect 18601 13883 18659 13889
rect 19521 13923 19579 13929
rect 19521 13889 19533 13923
rect 19567 13889 19579 13923
rect 19521 13883 19579 13889
rect 19788 13883 19800 13929
rect 19852 13920 19858 13932
rect 23290 13920 23296 13932
rect 19852 13892 19888 13920
rect 23251 13892 23296 13920
rect 19794 13880 19800 13883
rect 19852 13880 19858 13892
rect 23290 13880 23296 13892
rect 23348 13880 23354 13932
rect 23382 13880 23388 13932
rect 23440 13920 23446 13932
rect 25133 13923 25191 13929
rect 23440 13892 23485 13920
rect 23440 13880 23446 13892
rect 25133 13889 25145 13923
rect 25179 13889 25191 13923
rect 25133 13883 25191 13889
rect 1486 13852 1492 13864
rect 1447 13824 1492 13852
rect 1486 13812 1492 13824
rect 1544 13812 1550 13864
rect 1670 13852 1676 13864
rect 1631 13824 1676 13852
rect 1670 13812 1676 13824
rect 1728 13812 1734 13864
rect 1946 13852 1952 13864
rect 1907 13824 1952 13852
rect 1946 13812 1952 13824
rect 2004 13812 2010 13864
rect 14550 13812 14556 13864
rect 14608 13852 14614 13864
rect 14608 13824 14780 13852
rect 14608 13812 14614 13824
rect 14752 13793 14780 13824
rect 23014 13812 23020 13864
rect 23072 13852 23078 13864
rect 23109 13855 23167 13861
rect 23109 13852 23121 13855
rect 23072 13824 23121 13852
rect 23072 13812 23078 13824
rect 23109 13821 23121 13824
rect 23155 13821 23167 13855
rect 25148 13852 25176 13883
rect 25406 13880 25412 13932
rect 25464 13920 25470 13932
rect 25777 13923 25835 13929
rect 25777 13920 25789 13923
rect 25464 13892 25789 13920
rect 25464 13880 25470 13892
rect 25777 13889 25789 13892
rect 25823 13889 25835 13923
rect 25777 13883 25835 13889
rect 25961 13923 26019 13929
rect 25961 13889 25973 13923
rect 26007 13889 26019 13923
rect 25961 13883 26019 13889
rect 27157 13923 27215 13929
rect 27157 13889 27169 13923
rect 27203 13889 27215 13923
rect 27798 13920 27804 13932
rect 27759 13892 27804 13920
rect 27157 13883 27215 13889
rect 25498 13852 25504 13864
rect 25148 13824 25504 13852
rect 23109 13815 23167 13821
rect 25498 13812 25504 13824
rect 25556 13852 25562 13864
rect 25976 13852 26004 13883
rect 25556 13824 26004 13852
rect 27172 13852 27200 13883
rect 27798 13880 27804 13892
rect 27856 13880 27862 13932
rect 27246 13852 27252 13864
rect 27172 13824 27252 13852
rect 25556 13812 25562 13824
rect 14737 13787 14795 13793
rect 14737 13753 14749 13787
rect 14783 13753 14795 13787
rect 14737 13747 14795 13753
rect 25682 13744 25688 13796
rect 25740 13784 25746 13796
rect 27172 13784 27200 13824
rect 27246 13812 27252 13824
rect 27304 13812 27310 13864
rect 25740 13756 27200 13784
rect 25740 13744 25746 13756
rect 15562 13676 15568 13728
rect 15620 13716 15626 13728
rect 15749 13719 15807 13725
rect 15749 13716 15761 13719
rect 15620 13688 15761 13716
rect 15620 13676 15626 13688
rect 15749 13685 15761 13688
rect 15795 13685 15807 13719
rect 15749 13679 15807 13685
rect 17126 13676 17132 13728
rect 17184 13716 17190 13728
rect 17221 13719 17279 13725
rect 17221 13716 17233 13719
rect 17184 13688 17233 13716
rect 17184 13676 17190 13688
rect 17221 13685 17233 13688
rect 17267 13685 17279 13719
rect 17402 13716 17408 13728
rect 17363 13688 17408 13716
rect 17221 13679 17279 13685
rect 17402 13676 17408 13688
rect 17460 13676 17466 13728
rect 25958 13716 25964 13728
rect 25919 13688 25964 13716
rect 25958 13676 25964 13688
rect 26016 13676 26022 13728
rect 1104 13626 28888 13648
rect 1104 13574 5582 13626
rect 5634 13574 5646 13626
rect 5698 13574 5710 13626
rect 5762 13574 5774 13626
rect 5826 13574 5838 13626
rect 5890 13574 14846 13626
rect 14898 13574 14910 13626
rect 14962 13574 14974 13626
rect 15026 13574 15038 13626
rect 15090 13574 15102 13626
rect 15154 13574 24110 13626
rect 24162 13574 24174 13626
rect 24226 13574 24238 13626
rect 24290 13574 24302 13626
rect 24354 13574 24366 13626
rect 24418 13574 28888 13626
rect 1104 13552 28888 13574
rect 1670 13472 1676 13524
rect 1728 13512 1734 13524
rect 1949 13515 2007 13521
rect 1949 13512 1961 13515
rect 1728 13484 1961 13512
rect 1728 13472 1734 13484
rect 1949 13481 1961 13484
rect 1995 13481 2007 13515
rect 14090 13512 14096 13524
rect 14051 13484 14096 13512
rect 1949 13475 2007 13481
rect 14090 13472 14096 13484
rect 14148 13472 14154 13524
rect 15565 13515 15623 13521
rect 15565 13481 15577 13515
rect 15611 13512 15623 13515
rect 16301 13515 16359 13521
rect 16301 13512 16313 13515
rect 15611 13484 16313 13512
rect 15611 13481 15623 13484
rect 15565 13475 15623 13481
rect 16301 13481 16313 13484
rect 16347 13481 16359 13515
rect 16301 13475 16359 13481
rect 19794 13472 19800 13524
rect 19852 13512 19858 13524
rect 19889 13515 19947 13521
rect 19889 13512 19901 13515
rect 19852 13484 19901 13512
rect 19852 13472 19858 13484
rect 19889 13481 19901 13484
rect 19935 13481 19947 13515
rect 25682 13512 25688 13524
rect 19889 13475 19947 13481
rect 24780 13484 25688 13512
rect 21174 13404 21180 13456
rect 21232 13444 21238 13456
rect 21232 13416 22094 13444
rect 21232 13404 21238 13416
rect 21358 13336 21364 13388
rect 21416 13376 21422 13388
rect 21545 13379 21603 13385
rect 21545 13376 21557 13379
rect 21416 13348 21557 13376
rect 21416 13336 21422 13348
rect 21545 13345 21557 13348
rect 21591 13345 21603 13379
rect 21545 13339 21603 13345
rect 21729 13379 21787 13385
rect 21729 13345 21741 13379
rect 21775 13376 21787 13379
rect 22066 13376 22094 13416
rect 23109 13379 23167 13385
rect 23109 13376 23121 13379
rect 21775 13348 21864 13376
rect 21775 13345 21787 13348
rect 21729 13339 21787 13345
rect 2041 13311 2099 13317
rect 2041 13277 2053 13311
rect 2087 13308 2099 13311
rect 2130 13308 2136 13320
rect 2087 13280 2136 13308
rect 2087 13277 2099 13280
rect 2041 13271 2099 13277
rect 2130 13268 2136 13280
rect 2188 13308 2194 13320
rect 2774 13308 2780 13320
rect 2188 13280 2780 13308
rect 2188 13268 2194 13280
rect 2774 13268 2780 13280
rect 2832 13268 2838 13320
rect 14274 13308 14280 13320
rect 14235 13280 14280 13308
rect 14274 13268 14280 13280
rect 14332 13268 14338 13320
rect 15470 13268 15476 13320
rect 15528 13308 15534 13320
rect 16209 13311 16267 13317
rect 16209 13308 16221 13311
rect 15528 13280 16221 13308
rect 15528 13268 15534 13280
rect 16209 13277 16221 13280
rect 16255 13277 16267 13311
rect 16209 13271 16267 13277
rect 16393 13311 16451 13317
rect 16393 13277 16405 13311
rect 16439 13308 16451 13311
rect 16850 13308 16856 13320
rect 16439 13280 16856 13308
rect 16439 13277 16451 13280
rect 16393 13271 16451 13277
rect 16850 13268 16856 13280
rect 16908 13268 16914 13320
rect 16945 13311 17003 13317
rect 16945 13277 16957 13311
rect 16991 13308 17003 13311
rect 17586 13308 17592 13320
rect 16991 13280 17592 13308
rect 16991 13277 17003 13280
rect 16945 13271 17003 13277
rect 17328 13252 17356 13280
rect 17586 13268 17592 13280
rect 17644 13268 17650 13320
rect 20070 13308 20076 13320
rect 20031 13280 20076 13308
rect 20070 13268 20076 13280
rect 20128 13268 20134 13320
rect 15378 13240 15384 13252
rect 15339 13212 15384 13240
rect 15378 13200 15384 13212
rect 15436 13200 15442 13252
rect 17218 13249 17224 13252
rect 17212 13240 17224 13249
rect 17179 13212 17224 13240
rect 17212 13203 17224 13212
rect 17218 13200 17224 13203
rect 17276 13200 17282 13252
rect 17310 13200 17316 13252
rect 17368 13200 17374 13252
rect 21453 13243 21511 13249
rect 21453 13209 21465 13243
rect 21499 13240 21511 13243
rect 21836 13240 21864 13348
rect 22066 13348 23121 13376
rect 22066 13320 22094 13348
rect 23109 13345 23121 13348
rect 23155 13345 23167 13379
rect 23109 13339 23167 13345
rect 22002 13268 22008 13320
rect 22060 13280 22094 13320
rect 22833 13311 22891 13317
rect 22060 13268 22066 13280
rect 22833 13277 22845 13311
rect 22879 13308 22891 13311
rect 23382 13308 23388 13320
rect 22879 13280 23388 13308
rect 22879 13277 22891 13280
rect 22833 13271 22891 13277
rect 23382 13268 23388 13280
rect 23440 13268 23446 13320
rect 24670 13268 24676 13320
rect 24728 13308 24734 13320
rect 24780 13317 24808 13484
rect 25682 13472 25688 13484
rect 25740 13472 25746 13524
rect 25774 13472 25780 13524
rect 25832 13512 25838 13524
rect 25869 13515 25927 13521
rect 25869 13512 25881 13515
rect 25832 13484 25881 13512
rect 25832 13472 25838 13484
rect 25869 13481 25881 13484
rect 25915 13481 25927 13515
rect 25869 13475 25927 13481
rect 24857 13447 24915 13453
rect 24857 13413 24869 13447
rect 24903 13444 24915 13447
rect 26970 13444 26976 13456
rect 24903 13416 26976 13444
rect 24903 13413 24915 13416
rect 24857 13407 24915 13413
rect 26970 13404 26976 13416
rect 27028 13404 27034 13456
rect 25958 13376 25964 13388
rect 24964 13348 25964 13376
rect 24964 13317 24992 13348
rect 25958 13336 25964 13348
rect 26016 13336 26022 13388
rect 27522 13376 27528 13388
rect 27483 13348 27528 13376
rect 27522 13336 27528 13348
rect 27580 13336 27586 13388
rect 24765 13311 24823 13317
rect 24765 13308 24777 13311
rect 24728 13280 24777 13308
rect 24728 13268 24734 13280
rect 24765 13277 24777 13280
rect 24811 13277 24823 13311
rect 24765 13271 24823 13277
rect 24949 13311 25007 13317
rect 24949 13277 24961 13311
rect 24995 13277 25007 13311
rect 24949 13271 25007 13277
rect 25222 13268 25228 13320
rect 25280 13308 25286 13320
rect 25409 13311 25467 13317
rect 25409 13308 25421 13311
rect 25280 13280 25421 13308
rect 25280 13268 25286 13280
rect 25409 13277 25421 13280
rect 25455 13308 25467 13311
rect 25498 13308 25504 13320
rect 25455 13280 25504 13308
rect 25455 13277 25467 13280
rect 25409 13271 25467 13277
rect 25498 13268 25504 13280
rect 25556 13268 25562 13320
rect 26234 13268 26240 13320
rect 26292 13308 26298 13320
rect 26329 13311 26387 13317
rect 26329 13308 26341 13311
rect 26292 13280 26341 13308
rect 26292 13268 26298 13280
rect 26329 13277 26341 13280
rect 26375 13277 26387 13311
rect 26329 13271 26387 13277
rect 23566 13240 23572 13252
rect 21499 13212 21772 13240
rect 21836 13212 23572 13240
rect 21499 13209 21511 13212
rect 21453 13203 21511 13209
rect 15562 13132 15568 13184
rect 15620 13181 15626 13184
rect 15620 13175 15639 13181
rect 15627 13141 15639 13175
rect 15746 13172 15752 13184
rect 15707 13144 15752 13172
rect 15620 13135 15639 13141
rect 15620 13132 15626 13135
rect 15746 13132 15752 13144
rect 15804 13132 15810 13184
rect 18322 13172 18328 13184
rect 18283 13144 18328 13172
rect 18322 13132 18328 13144
rect 18380 13132 18386 13184
rect 20990 13132 20996 13184
rect 21048 13172 21054 13184
rect 21085 13175 21143 13181
rect 21085 13172 21097 13175
rect 21048 13144 21097 13172
rect 21048 13132 21054 13144
rect 21085 13141 21097 13144
rect 21131 13141 21143 13175
rect 21744 13172 21772 13212
rect 23566 13200 23572 13212
rect 23624 13240 23630 13252
rect 24026 13240 24032 13252
rect 23624 13212 24032 13240
rect 23624 13200 23630 13212
rect 24026 13200 24032 13212
rect 24084 13200 24090 13252
rect 26513 13243 26571 13249
rect 26513 13209 26525 13243
rect 26559 13240 26571 13243
rect 28074 13240 28080 13252
rect 26559 13212 28080 13240
rect 26559 13209 26571 13212
rect 26513 13203 26571 13209
rect 28074 13200 28080 13212
rect 28132 13200 28138 13252
rect 23198 13172 23204 13184
rect 21744 13144 23204 13172
rect 21085 13135 21143 13141
rect 23198 13132 23204 13144
rect 23256 13132 23262 13184
rect 1104 13082 28888 13104
rect 1104 13030 10214 13082
rect 10266 13030 10278 13082
rect 10330 13030 10342 13082
rect 10394 13030 10406 13082
rect 10458 13030 10470 13082
rect 10522 13030 19478 13082
rect 19530 13030 19542 13082
rect 19594 13030 19606 13082
rect 19658 13030 19670 13082
rect 19722 13030 19734 13082
rect 19786 13030 28888 13082
rect 1104 13008 28888 13030
rect 16114 12968 16120 12980
rect 16075 12940 16120 12968
rect 16114 12928 16120 12940
rect 16172 12928 16178 12980
rect 23198 12968 23204 12980
rect 23159 12940 23204 12968
rect 23198 12928 23204 12940
rect 23256 12968 23262 12980
rect 24305 12971 24363 12977
rect 24305 12968 24317 12971
rect 23256 12940 24317 12968
rect 23256 12928 23262 12940
rect 24305 12937 24317 12940
rect 24351 12937 24363 12971
rect 24670 12968 24676 12980
rect 24631 12940 24676 12968
rect 24305 12931 24363 12937
rect 24670 12928 24676 12940
rect 24728 12928 24734 12980
rect 28074 12968 28080 12980
rect 28035 12940 28080 12968
rect 28074 12928 28080 12940
rect 28132 12928 28138 12980
rect 17310 12900 17316 12912
rect 14936 12872 17316 12900
rect 1486 12792 1492 12844
rect 1544 12832 1550 12844
rect 1581 12835 1639 12841
rect 1581 12832 1593 12835
rect 1544 12804 1593 12832
rect 1544 12792 1550 12804
rect 1581 12801 1593 12804
rect 1627 12801 1639 12835
rect 14734 12832 14740 12844
rect 14647 12804 14740 12832
rect 1581 12795 1639 12801
rect 14734 12792 14740 12804
rect 14792 12832 14798 12844
rect 14936 12832 14964 12872
rect 17310 12860 17316 12872
rect 17368 12860 17374 12912
rect 17497 12903 17555 12909
rect 17497 12869 17509 12903
rect 17543 12900 17555 12903
rect 18322 12900 18328 12912
rect 17543 12872 18328 12900
rect 17543 12869 17555 12872
rect 17497 12863 17555 12869
rect 18322 12860 18328 12872
rect 18380 12860 18386 12912
rect 14792 12804 14964 12832
rect 15004 12835 15062 12841
rect 14792 12792 14798 12804
rect 15004 12801 15016 12835
rect 15050 12832 15062 12835
rect 15562 12832 15568 12844
rect 15050 12804 15568 12832
rect 15050 12801 15062 12804
rect 15004 12795 15062 12801
rect 15562 12792 15568 12804
rect 15620 12792 15626 12844
rect 17681 12835 17739 12841
rect 17681 12801 17693 12835
rect 17727 12832 17739 12835
rect 17770 12832 17776 12844
rect 17727 12804 17776 12832
rect 17727 12801 17739 12804
rect 17681 12795 17739 12801
rect 17770 12792 17776 12804
rect 17828 12792 17834 12844
rect 20806 12832 20812 12844
rect 20767 12804 20812 12832
rect 20806 12792 20812 12804
rect 20864 12792 20870 12844
rect 20990 12832 20996 12844
rect 20951 12804 20996 12832
rect 20990 12792 20996 12804
rect 21048 12792 21054 12844
rect 22094 12841 22100 12844
rect 22088 12795 22100 12841
rect 22152 12832 22158 12844
rect 22152 12804 22188 12832
rect 22094 12792 22100 12795
rect 22152 12792 22158 12804
rect 23842 12792 23848 12844
rect 23900 12832 23906 12844
rect 24213 12835 24271 12841
rect 24213 12832 24225 12835
rect 23900 12804 24225 12832
rect 23900 12792 23906 12804
rect 24213 12801 24225 12804
rect 24259 12801 24271 12835
rect 24213 12795 24271 12801
rect 25406 12792 25412 12844
rect 25464 12832 25470 12844
rect 25593 12835 25651 12841
rect 25593 12832 25605 12835
rect 25464 12804 25605 12832
rect 25464 12792 25470 12804
rect 25593 12801 25605 12804
rect 25639 12832 25651 12835
rect 25682 12832 25688 12844
rect 25639 12804 25688 12832
rect 25639 12801 25651 12804
rect 25593 12795 25651 12801
rect 25682 12792 25688 12804
rect 25740 12792 25746 12844
rect 25866 12832 25872 12844
rect 25827 12804 25872 12832
rect 25866 12792 25872 12804
rect 25924 12832 25930 12844
rect 27157 12835 27215 12841
rect 27157 12832 27169 12835
rect 25924 12804 27169 12832
rect 25924 12792 25930 12804
rect 27157 12801 27169 12804
rect 27203 12801 27215 12835
rect 27157 12795 27215 12801
rect 27433 12835 27491 12841
rect 27433 12801 27445 12835
rect 27479 12832 27491 12835
rect 27706 12832 27712 12844
rect 27479 12804 27712 12832
rect 27479 12801 27491 12804
rect 27433 12795 27491 12801
rect 27706 12792 27712 12804
rect 27764 12792 27770 12844
rect 27982 12832 27988 12844
rect 27943 12804 27988 12832
rect 27982 12792 27988 12804
rect 28040 12792 28046 12844
rect 17126 12724 17132 12776
rect 17184 12764 17190 12776
rect 17313 12767 17371 12773
rect 17313 12764 17325 12767
rect 17184 12736 17325 12764
rect 17184 12724 17190 12736
rect 17313 12733 17325 12736
rect 17359 12733 17371 12767
rect 21818 12764 21824 12776
rect 21779 12736 21824 12764
rect 17313 12727 17371 12733
rect 21818 12724 21824 12736
rect 21876 12724 21882 12776
rect 24121 12767 24179 12773
rect 24121 12733 24133 12767
rect 24167 12764 24179 12767
rect 24486 12764 24492 12776
rect 24167 12736 24492 12764
rect 24167 12733 24179 12736
rect 24121 12727 24179 12733
rect 24486 12724 24492 12736
rect 24544 12724 24550 12776
rect 25958 12724 25964 12776
rect 26016 12764 26022 12776
rect 27341 12767 27399 12773
rect 27341 12764 27353 12767
rect 26016 12736 27353 12764
rect 26016 12724 26022 12736
rect 27341 12733 27353 12736
rect 27387 12733 27399 12767
rect 27341 12727 27399 12733
rect 26878 12656 26884 12708
rect 26936 12696 26942 12708
rect 27249 12699 27307 12705
rect 27249 12696 27261 12699
rect 26936 12668 27261 12696
rect 26936 12656 26942 12668
rect 27249 12665 27261 12668
rect 27295 12665 27307 12699
rect 27249 12659 27307 12665
rect 21082 12588 21088 12640
rect 21140 12628 21146 12640
rect 21177 12631 21235 12637
rect 21177 12628 21189 12631
rect 21140 12600 21189 12628
rect 21140 12588 21146 12600
rect 21177 12597 21189 12600
rect 21223 12597 21235 12631
rect 26970 12628 26976 12640
rect 26931 12600 26976 12628
rect 21177 12591 21235 12597
rect 26970 12588 26976 12600
rect 27028 12588 27034 12640
rect 1104 12538 28888 12560
rect 1104 12486 5582 12538
rect 5634 12486 5646 12538
rect 5698 12486 5710 12538
rect 5762 12486 5774 12538
rect 5826 12486 5838 12538
rect 5890 12486 14846 12538
rect 14898 12486 14910 12538
rect 14962 12486 14974 12538
rect 15026 12486 15038 12538
rect 15090 12486 15102 12538
rect 15154 12486 24110 12538
rect 24162 12486 24174 12538
rect 24226 12486 24238 12538
rect 24290 12486 24302 12538
rect 24354 12486 24366 12538
rect 24418 12486 28888 12538
rect 1104 12464 28888 12486
rect 15562 12424 15568 12436
rect 15523 12396 15568 12424
rect 15562 12384 15568 12396
rect 15620 12384 15626 12436
rect 17218 12424 17224 12436
rect 17179 12396 17224 12424
rect 17218 12384 17224 12396
rect 17276 12384 17282 12436
rect 21269 12427 21327 12433
rect 21269 12393 21281 12427
rect 21315 12424 21327 12427
rect 22094 12424 22100 12436
rect 21315 12396 22100 12424
rect 21315 12393 21327 12396
rect 21269 12387 21327 12393
rect 22094 12384 22100 12396
rect 22152 12384 22158 12436
rect 23842 12424 23848 12436
rect 23803 12396 23848 12424
rect 23842 12384 23848 12396
rect 23900 12384 23906 12436
rect 27706 12424 27712 12436
rect 27667 12396 27712 12424
rect 27706 12384 27712 12396
rect 27764 12384 27770 12436
rect 26326 12316 26332 12368
rect 26384 12356 26390 12368
rect 26881 12359 26939 12365
rect 26881 12356 26893 12359
rect 26384 12328 26893 12356
rect 26384 12316 26390 12328
rect 26881 12325 26893 12328
rect 26927 12325 26939 12359
rect 26881 12319 26939 12325
rect 20714 12248 20720 12300
rect 20772 12288 20778 12300
rect 21818 12288 21824 12300
rect 20772 12260 21824 12288
rect 20772 12248 20778 12260
rect 21818 12248 21824 12260
rect 21876 12288 21882 12300
rect 22465 12291 22523 12297
rect 22465 12288 22477 12291
rect 21876 12260 22477 12288
rect 21876 12248 21882 12260
rect 22465 12257 22477 12260
rect 22511 12257 22523 12291
rect 22465 12251 22523 12257
rect 26142 12248 26148 12300
rect 26200 12288 26206 12300
rect 26421 12291 26479 12297
rect 26421 12288 26433 12291
rect 26200 12260 26433 12288
rect 26200 12248 26206 12260
rect 26421 12257 26433 12260
rect 26467 12257 26479 12291
rect 26421 12251 26479 12257
rect 27338 12248 27344 12300
rect 27396 12288 27402 12300
rect 27706 12288 27712 12300
rect 27396 12260 27712 12288
rect 27396 12248 27402 12260
rect 27706 12248 27712 12260
rect 27764 12248 27770 12300
rect 1486 12220 1492 12232
rect 1447 12192 1492 12220
rect 1486 12180 1492 12192
rect 1544 12180 1550 12232
rect 15746 12220 15752 12232
rect 15707 12192 15752 12220
rect 15746 12180 15752 12192
rect 15804 12180 15810 12232
rect 17402 12220 17408 12232
rect 17363 12192 17408 12220
rect 17402 12180 17408 12192
rect 17460 12180 17466 12232
rect 18690 12180 18696 12232
rect 18748 12220 18754 12232
rect 19245 12223 19303 12229
rect 19245 12220 19257 12223
rect 18748 12192 19257 12220
rect 18748 12180 18754 12192
rect 19245 12189 19257 12192
rect 19291 12189 19303 12223
rect 21082 12220 21088 12232
rect 21043 12192 21088 12220
rect 19245 12183 19303 12189
rect 21082 12180 21088 12192
rect 21140 12180 21146 12232
rect 24581 12223 24639 12229
rect 24581 12220 24593 12223
rect 22066 12192 24593 12220
rect 3326 12112 3332 12164
rect 3384 12152 3390 12164
rect 22066 12152 22094 12192
rect 24581 12189 24593 12192
rect 24627 12189 24639 12223
rect 26878 12220 26884 12232
rect 26839 12192 26884 12220
rect 24581 12183 24639 12189
rect 26878 12180 26884 12192
rect 26936 12180 26942 12232
rect 27157 12223 27215 12229
rect 27157 12189 27169 12223
rect 27203 12189 27215 12223
rect 27157 12183 27215 12189
rect 3384 12124 22094 12152
rect 22732 12155 22790 12161
rect 3384 12112 3390 12124
rect 22732 12121 22744 12155
rect 22778 12152 22790 12155
rect 22830 12152 22836 12164
rect 22778 12124 22836 12152
rect 22778 12121 22790 12124
rect 22732 12115 22790 12121
rect 22830 12112 22836 12124
rect 22888 12112 22894 12164
rect 24946 12112 24952 12164
rect 25004 12152 25010 12164
rect 26237 12155 26295 12161
rect 26237 12152 26249 12155
rect 25004 12124 26249 12152
rect 25004 12112 25010 12124
rect 26237 12121 26249 12124
rect 26283 12121 26295 12155
rect 26237 12115 26295 12121
rect 26418 12112 26424 12164
rect 26476 12152 26482 12164
rect 27172 12152 27200 12183
rect 27246 12180 27252 12232
rect 27304 12220 27310 12232
rect 27617 12223 27675 12229
rect 27617 12220 27629 12223
rect 27304 12192 27629 12220
rect 27304 12180 27310 12192
rect 27617 12189 27629 12192
rect 27663 12189 27675 12223
rect 27617 12183 27675 12189
rect 27801 12223 27859 12229
rect 27801 12189 27813 12223
rect 27847 12189 27859 12223
rect 27801 12183 27859 12189
rect 27816 12152 27844 12183
rect 26476 12124 27844 12152
rect 26476 12112 26482 12124
rect 19334 12084 19340 12096
rect 19295 12056 19340 12084
rect 19334 12044 19340 12056
rect 19392 12044 19398 12096
rect 25866 12044 25872 12096
rect 25924 12084 25930 12096
rect 27065 12087 27123 12093
rect 27065 12084 27077 12087
rect 25924 12056 27077 12084
rect 25924 12044 25930 12056
rect 27065 12053 27077 12056
rect 27111 12053 27123 12087
rect 27065 12047 27123 12053
rect 1104 11994 28888 12016
rect 1104 11942 10214 11994
rect 10266 11942 10278 11994
rect 10330 11942 10342 11994
rect 10394 11942 10406 11994
rect 10458 11942 10470 11994
rect 10522 11942 19478 11994
rect 19530 11942 19542 11994
rect 19594 11942 19606 11994
rect 19658 11942 19670 11994
rect 19722 11942 19734 11994
rect 19786 11942 28888 11994
rect 1104 11920 28888 11942
rect 18414 11840 18420 11892
rect 18472 11880 18478 11892
rect 19153 11883 19211 11889
rect 19153 11880 19165 11883
rect 18472 11852 19165 11880
rect 18472 11840 18478 11852
rect 19153 11849 19165 11852
rect 19199 11849 19211 11883
rect 19153 11843 19211 11849
rect 19613 11883 19671 11889
rect 19613 11849 19625 11883
rect 19659 11880 19671 11883
rect 19886 11880 19892 11892
rect 19659 11852 19892 11880
rect 19659 11849 19671 11852
rect 19613 11843 19671 11849
rect 19886 11840 19892 11852
rect 19944 11840 19950 11892
rect 22830 11880 22836 11892
rect 22791 11852 22836 11880
rect 22830 11840 22836 11852
rect 22888 11840 22894 11892
rect 23290 11840 23296 11892
rect 23348 11880 23354 11892
rect 23477 11883 23535 11889
rect 23477 11880 23489 11883
rect 23348 11852 23489 11880
rect 23348 11840 23354 11852
rect 23477 11849 23489 11852
rect 23523 11849 23535 11883
rect 23934 11880 23940 11892
rect 23895 11852 23940 11880
rect 23477 11843 23535 11849
rect 23934 11840 23940 11852
rect 23992 11840 23998 11892
rect 24946 11880 24952 11892
rect 24907 11852 24952 11880
rect 24946 11840 24952 11852
rect 25004 11840 25010 11892
rect 25961 11883 26019 11889
rect 25961 11849 25973 11883
rect 26007 11880 26019 11883
rect 26418 11880 26424 11892
rect 26007 11852 26424 11880
rect 26007 11849 26019 11852
rect 25961 11843 26019 11849
rect 26418 11840 26424 11852
rect 26476 11840 26482 11892
rect 17681 11815 17739 11821
rect 17681 11781 17693 11815
rect 17727 11812 17739 11815
rect 19334 11812 19340 11824
rect 17727 11784 19340 11812
rect 17727 11781 17739 11784
rect 17681 11775 17739 11781
rect 19334 11772 19340 11784
rect 19392 11812 19398 11824
rect 19797 11815 19855 11821
rect 19797 11812 19809 11815
rect 19392 11784 19809 11812
rect 19392 11772 19398 11784
rect 19797 11781 19809 11784
rect 19843 11781 19855 11815
rect 22002 11812 22008 11824
rect 19797 11775 19855 11781
rect 20548 11784 22008 11812
rect 1486 11744 1492 11756
rect 1447 11716 1492 11744
rect 1486 11704 1492 11716
rect 1544 11704 1550 11756
rect 15470 11704 15476 11756
rect 15528 11744 15534 11756
rect 17313 11747 17371 11753
rect 17313 11744 17325 11747
rect 15528 11716 17325 11744
rect 15528 11704 15534 11716
rect 17313 11713 17325 11716
rect 17359 11713 17371 11747
rect 17313 11707 17371 11713
rect 17773 11747 17831 11753
rect 17773 11713 17785 11747
rect 17819 11744 17831 11747
rect 17862 11744 17868 11756
rect 17819 11716 17868 11744
rect 17819 11713 17831 11716
rect 17773 11707 17831 11713
rect 17862 11704 17868 11716
rect 17920 11704 17926 11756
rect 18690 11744 18696 11756
rect 18651 11716 18696 11744
rect 18690 11704 18696 11716
rect 18748 11704 18754 11756
rect 19978 11744 19984 11756
rect 19939 11716 19984 11744
rect 19978 11704 19984 11716
rect 20036 11704 20042 11756
rect 20548 11753 20576 11784
rect 22002 11772 22008 11784
rect 22060 11772 22066 11824
rect 23842 11812 23848 11824
rect 23803 11784 23848 11812
rect 23842 11772 23848 11784
rect 23900 11772 23906 11824
rect 25222 11772 25228 11824
rect 25280 11812 25286 11824
rect 25593 11815 25651 11821
rect 25593 11812 25605 11815
rect 25280 11784 25605 11812
rect 25280 11772 25286 11784
rect 25593 11781 25605 11784
rect 25639 11781 25651 11815
rect 25593 11775 25651 11781
rect 25682 11772 25688 11824
rect 25740 11812 25746 11824
rect 25777 11815 25835 11821
rect 25777 11812 25789 11815
rect 25740 11784 25789 11812
rect 25740 11772 25746 11784
rect 25777 11781 25789 11784
rect 25823 11781 25835 11815
rect 25777 11775 25835 11781
rect 20533 11747 20591 11753
rect 20533 11713 20545 11747
rect 20579 11713 20591 11747
rect 20533 11707 20591 11713
rect 20625 11747 20683 11753
rect 20625 11713 20637 11747
rect 20671 11744 20683 11747
rect 20898 11744 20904 11756
rect 20671 11716 20904 11744
rect 20671 11713 20683 11716
rect 20625 11707 20683 11713
rect 20898 11704 20904 11716
rect 20956 11704 20962 11756
rect 23014 11744 23020 11756
rect 22975 11716 23020 11744
rect 23014 11704 23020 11716
rect 23072 11704 23078 11756
rect 24857 11747 24915 11753
rect 24857 11713 24869 11747
rect 24903 11744 24915 11747
rect 25038 11744 25044 11756
rect 24903 11716 25044 11744
rect 24903 11713 24915 11716
rect 24857 11707 24915 11713
rect 25038 11704 25044 11716
rect 25096 11704 25102 11756
rect 27985 11747 28043 11753
rect 27985 11713 27997 11747
rect 28031 11744 28043 11747
rect 28166 11744 28172 11756
rect 28031 11716 28172 11744
rect 28031 11713 28043 11716
rect 27985 11707 28043 11713
rect 28166 11704 28172 11716
rect 28224 11704 28230 11756
rect 1673 11679 1731 11685
rect 1673 11645 1685 11679
rect 1719 11676 1731 11679
rect 1854 11676 1860 11688
rect 1719 11648 1860 11676
rect 1719 11645 1731 11648
rect 1673 11639 1731 11645
rect 1854 11636 1860 11648
rect 1912 11636 1918 11688
rect 1946 11636 1952 11688
rect 2004 11676 2010 11688
rect 24026 11676 24032 11688
rect 2004 11648 2049 11676
rect 23987 11648 24032 11676
rect 2004 11636 2010 11648
rect 24026 11636 24032 11648
rect 24084 11636 24090 11688
rect 19061 11611 19119 11617
rect 19061 11577 19073 11611
rect 19107 11608 19119 11611
rect 19334 11608 19340 11620
rect 19107 11580 19340 11608
rect 19107 11577 19119 11580
rect 19061 11571 19119 11577
rect 19334 11568 19340 11580
rect 19392 11568 19398 11620
rect 17497 11543 17555 11549
rect 17497 11509 17509 11543
rect 17543 11540 17555 11543
rect 17586 11540 17592 11552
rect 17543 11512 17592 11540
rect 17543 11509 17555 11512
rect 17497 11503 17555 11509
rect 17586 11500 17592 11512
rect 17644 11500 17650 11552
rect 20809 11543 20867 11549
rect 20809 11509 20821 11543
rect 20855 11540 20867 11543
rect 21358 11540 21364 11552
rect 20855 11512 21364 11540
rect 20855 11509 20867 11512
rect 20809 11503 20867 11509
rect 21358 11500 21364 11512
rect 21416 11500 21422 11552
rect 27341 11543 27399 11549
rect 27341 11509 27353 11543
rect 27387 11540 27399 11543
rect 27890 11540 27896 11552
rect 27387 11512 27896 11540
rect 27387 11509 27399 11512
rect 27341 11503 27399 11509
rect 27890 11500 27896 11512
rect 27948 11500 27954 11552
rect 1104 11450 28888 11472
rect 1104 11398 5582 11450
rect 5634 11398 5646 11450
rect 5698 11398 5710 11450
rect 5762 11398 5774 11450
rect 5826 11398 5838 11450
rect 5890 11398 14846 11450
rect 14898 11398 14910 11450
rect 14962 11398 14974 11450
rect 15026 11398 15038 11450
rect 15090 11398 15102 11450
rect 15154 11398 24110 11450
rect 24162 11398 24174 11450
rect 24226 11398 24238 11450
rect 24290 11398 24302 11450
rect 24354 11398 24366 11450
rect 24418 11398 28888 11450
rect 1104 11376 28888 11398
rect 1854 11336 1860 11348
rect 1815 11308 1860 11336
rect 1854 11296 1860 11308
rect 1912 11296 1918 11348
rect 18690 11336 18696 11348
rect 18651 11308 18696 11336
rect 18690 11296 18696 11308
rect 18748 11296 18754 11348
rect 25869 11339 25927 11345
rect 25869 11305 25881 11339
rect 25915 11336 25927 11339
rect 26234 11336 26240 11348
rect 25915 11308 26240 11336
rect 25915 11305 25927 11308
rect 25869 11299 25927 11305
rect 26234 11296 26240 11308
rect 26292 11296 26298 11348
rect 21177 11271 21235 11277
rect 21177 11237 21189 11271
rect 21223 11237 21235 11271
rect 21177 11231 21235 11237
rect 13814 11160 13820 11212
rect 13872 11200 13878 11212
rect 16942 11200 16948 11212
rect 13872 11172 16948 11200
rect 13872 11160 13878 11172
rect 1949 11135 2007 11141
rect 1949 11101 1961 11135
rect 1995 11132 2007 11135
rect 2038 11132 2044 11144
rect 1995 11104 2044 11132
rect 1995 11101 2007 11104
rect 1949 11095 2007 11101
rect 2038 11092 2044 11104
rect 2096 11092 2102 11144
rect 15396 11141 15424 11172
rect 16942 11160 16948 11172
rect 17000 11160 17006 11212
rect 17310 11200 17316 11212
rect 17271 11172 17316 11200
rect 17310 11160 17316 11172
rect 17368 11160 17374 11212
rect 20714 11200 20720 11212
rect 20675 11172 20720 11200
rect 20714 11160 20720 11172
rect 20772 11160 20778 11212
rect 15381 11135 15439 11141
rect 15381 11101 15393 11135
rect 15427 11101 15439 11135
rect 15381 11095 15439 11101
rect 16485 11135 16543 11141
rect 16485 11101 16497 11135
rect 16531 11132 16543 11135
rect 16574 11132 16580 11144
rect 16531 11104 16580 11132
rect 16531 11101 16543 11104
rect 16485 11095 16543 11101
rect 16574 11092 16580 11104
rect 16632 11092 16638 11144
rect 17586 11141 17592 11144
rect 16669 11135 16727 11141
rect 16669 11101 16681 11135
rect 16715 11101 16727 11135
rect 17580 11132 17592 11141
rect 17547 11104 17592 11132
rect 16669 11095 16727 11101
rect 17580 11095 17592 11104
rect 16684 11064 16712 11095
rect 17586 11092 17592 11095
rect 17644 11092 17650 11144
rect 20461 11135 20519 11141
rect 20461 11101 20473 11135
rect 20507 11132 20519 11135
rect 21192 11132 21220 11231
rect 27522 11200 27528 11212
rect 27483 11172 27528 11200
rect 27522 11160 27528 11172
rect 27580 11160 27586 11212
rect 27890 11160 27896 11212
rect 27948 11200 27954 11212
rect 28169 11203 28227 11209
rect 28169 11200 28181 11203
rect 27948 11172 28181 11200
rect 27948 11160 27954 11172
rect 28169 11169 28181 11172
rect 28215 11169 28227 11203
rect 28169 11163 28227 11169
rect 21358 11132 21364 11144
rect 20507 11104 21220 11132
rect 21319 11104 21364 11132
rect 20507 11101 20519 11104
rect 20461 11095 20519 11101
rect 21358 11092 21364 11104
rect 21416 11092 21422 11144
rect 19242 11064 19248 11076
rect 16684 11036 19248 11064
rect 19242 11024 19248 11036
rect 19300 11024 19306 11076
rect 27982 11064 27988 11076
rect 27943 11036 27988 11064
rect 27982 11024 27988 11036
rect 28040 11024 28046 11076
rect 15562 10996 15568 11008
rect 15523 10968 15568 10996
rect 15562 10956 15568 10968
rect 15620 10956 15626 11008
rect 15930 10956 15936 11008
rect 15988 10996 15994 11008
rect 16301 10999 16359 11005
rect 16301 10996 16313 10999
rect 15988 10968 16313 10996
rect 15988 10956 15994 10968
rect 16301 10965 16313 10968
rect 16347 10965 16359 10999
rect 19334 10996 19340 11008
rect 19295 10968 19340 10996
rect 16301 10959 16359 10965
rect 19334 10956 19340 10968
rect 19392 10956 19398 11008
rect 1104 10906 28888 10928
rect 1104 10854 10214 10906
rect 10266 10854 10278 10906
rect 10330 10854 10342 10906
rect 10394 10854 10406 10906
rect 10458 10854 10470 10906
rect 10522 10854 19478 10906
rect 19530 10854 19542 10906
rect 19594 10854 19606 10906
rect 19658 10854 19670 10906
rect 19722 10854 19734 10906
rect 19786 10854 28888 10906
rect 1104 10832 28888 10854
rect 17678 10752 17684 10804
rect 17736 10792 17742 10804
rect 18049 10795 18107 10801
rect 18049 10792 18061 10795
rect 17736 10764 18061 10792
rect 17736 10752 17742 10764
rect 18049 10761 18061 10764
rect 18095 10761 18107 10795
rect 18049 10755 18107 10761
rect 19334 10752 19340 10804
rect 19392 10792 19398 10804
rect 19978 10792 19984 10804
rect 19392 10764 19984 10792
rect 19392 10752 19398 10764
rect 19978 10752 19984 10764
rect 20036 10792 20042 10804
rect 20533 10795 20591 10801
rect 20533 10792 20545 10795
rect 20036 10764 20545 10792
rect 20036 10752 20042 10764
rect 20533 10761 20545 10764
rect 20579 10761 20591 10795
rect 20898 10792 20904 10804
rect 20859 10764 20904 10792
rect 20533 10755 20591 10761
rect 20898 10752 20904 10764
rect 20956 10752 20962 10804
rect 27801 10795 27859 10801
rect 27801 10761 27813 10795
rect 27847 10792 27859 10795
rect 27982 10792 27988 10804
rect 27847 10764 27988 10792
rect 27847 10761 27859 10764
rect 27801 10755 27859 10761
rect 27982 10752 27988 10764
rect 28040 10752 28046 10804
rect 17310 10724 17316 10736
rect 16684 10696 17316 10724
rect 15930 10656 15936 10668
rect 15891 10628 15936 10656
rect 15930 10616 15936 10628
rect 15988 10616 15994 10668
rect 16684 10665 16712 10696
rect 17310 10684 17316 10696
rect 17368 10684 17374 10736
rect 16669 10659 16727 10665
rect 16669 10625 16681 10659
rect 16715 10625 16727 10659
rect 16925 10659 16983 10665
rect 16925 10656 16937 10659
rect 16669 10619 16727 10625
rect 16776 10628 16937 10656
rect 16776 10588 16804 10628
rect 16925 10625 16937 10628
rect 16971 10625 16983 10659
rect 16925 10619 16983 10625
rect 27614 10616 27620 10668
rect 27672 10656 27678 10668
rect 27709 10659 27767 10665
rect 27709 10656 27721 10659
rect 27672 10628 27721 10656
rect 27672 10616 27678 10628
rect 27709 10625 27721 10628
rect 27755 10625 27767 10659
rect 27709 10619 27767 10625
rect 20254 10588 20260 10600
rect 16132 10560 16804 10588
rect 20215 10560 20260 10588
rect 16132 10529 16160 10560
rect 20254 10548 20260 10560
rect 20312 10548 20318 10600
rect 20438 10588 20444 10600
rect 20399 10560 20444 10588
rect 20438 10548 20444 10560
rect 20496 10548 20502 10600
rect 25958 10588 25964 10600
rect 25919 10560 25964 10588
rect 25958 10548 25964 10560
rect 26016 10548 26022 10600
rect 26234 10548 26240 10600
rect 26292 10588 26298 10600
rect 26421 10591 26479 10597
rect 26292 10560 26337 10588
rect 26292 10548 26298 10560
rect 26421 10557 26433 10591
rect 26467 10588 26479 10591
rect 27065 10591 27123 10597
rect 27065 10588 27077 10591
rect 26467 10560 27077 10588
rect 26467 10557 26479 10560
rect 26421 10551 26479 10557
rect 27065 10557 27077 10560
rect 27111 10557 27123 10591
rect 27065 10551 27123 10557
rect 16117 10523 16175 10529
rect 16117 10489 16129 10523
rect 16163 10489 16175 10523
rect 16117 10483 16175 10489
rect 1394 10412 1400 10464
rect 1452 10452 1458 10464
rect 1489 10455 1547 10461
rect 1489 10452 1501 10455
rect 1452 10424 1501 10452
rect 1452 10412 1458 10424
rect 1489 10421 1501 10424
rect 1535 10421 1547 10455
rect 1489 10415 1547 10421
rect 1104 10362 28888 10384
rect 1104 10310 5582 10362
rect 5634 10310 5646 10362
rect 5698 10310 5710 10362
rect 5762 10310 5774 10362
rect 5826 10310 5838 10362
rect 5890 10310 14846 10362
rect 14898 10310 14910 10362
rect 14962 10310 14974 10362
rect 15026 10310 15038 10362
rect 15090 10310 15102 10362
rect 15154 10310 24110 10362
rect 24162 10310 24174 10362
rect 24226 10310 24238 10362
rect 24290 10310 24302 10362
rect 24354 10310 24366 10362
rect 24418 10310 28888 10362
rect 1104 10288 28888 10310
rect 16574 10208 16580 10260
rect 16632 10248 16638 10260
rect 16761 10251 16819 10257
rect 16761 10248 16773 10251
rect 16632 10220 16773 10248
rect 16632 10208 16638 10220
rect 16761 10217 16773 10220
rect 16807 10217 16819 10251
rect 16761 10211 16819 10217
rect 28350 10180 28356 10192
rect 2424 10152 28356 10180
rect 1762 10044 1768 10056
rect 1723 10016 1768 10044
rect 1762 10004 1768 10016
rect 1820 10004 1826 10056
rect 2424 10053 2452 10152
rect 28350 10140 28356 10152
rect 28408 10140 28414 10192
rect 15562 10072 15568 10124
rect 15620 10112 15626 10124
rect 17405 10115 17463 10121
rect 17405 10112 17417 10115
rect 15620 10084 17417 10112
rect 15620 10072 15626 10084
rect 17405 10081 17417 10084
rect 17451 10112 17463 10115
rect 20254 10112 20260 10124
rect 17451 10084 20260 10112
rect 17451 10081 17463 10084
rect 17405 10075 17463 10081
rect 20254 10072 20260 10084
rect 20312 10072 20318 10124
rect 25314 10112 25320 10124
rect 25275 10084 25320 10112
rect 25314 10072 25320 10084
rect 25372 10072 25378 10124
rect 26789 10115 26847 10121
rect 26789 10112 26801 10115
rect 25424 10084 26801 10112
rect 2409 10047 2467 10053
rect 2409 10013 2421 10047
rect 2455 10013 2467 10047
rect 2409 10007 2467 10013
rect 3053 10047 3111 10053
rect 3053 10013 3065 10047
rect 3099 10044 3111 10047
rect 3786 10044 3792 10056
rect 3099 10016 3792 10044
rect 3099 10013 3111 10016
rect 3053 10007 3111 10013
rect 3786 10004 3792 10016
rect 3844 10004 3850 10056
rect 17129 10047 17187 10053
rect 17129 10013 17141 10047
rect 17175 10044 17187 10047
rect 17678 10044 17684 10056
rect 17175 10016 17684 10044
rect 17175 10013 17187 10016
rect 17129 10007 17187 10013
rect 17678 10004 17684 10016
rect 17736 10004 17742 10056
rect 24673 10047 24731 10053
rect 24673 10013 24685 10047
rect 24719 10044 24731 10047
rect 25038 10044 25044 10056
rect 24719 10016 25044 10044
rect 24719 10013 24731 10016
rect 24673 10007 24731 10013
rect 25038 10004 25044 10016
rect 25096 10004 25102 10056
rect 24581 9979 24639 9985
rect 24581 9945 24593 9979
rect 24627 9976 24639 9979
rect 25424 9976 25452 10084
rect 26789 10081 26801 10084
rect 26835 10081 26847 10115
rect 26970 10112 26976 10124
rect 26931 10084 26976 10112
rect 26789 10075 26847 10081
rect 26970 10072 26976 10084
rect 27028 10072 27034 10124
rect 27433 10047 27491 10053
rect 27433 10013 27445 10047
rect 27479 10013 27491 10047
rect 27433 10007 27491 10013
rect 24627 9948 25452 9976
rect 24627 9945 24639 9948
rect 24581 9939 24639 9945
rect 1578 9868 1584 9920
rect 1636 9908 1642 9920
rect 1673 9911 1731 9917
rect 1673 9908 1685 9911
rect 1636 9880 1685 9908
rect 1636 9868 1642 9880
rect 1673 9877 1685 9880
rect 1719 9877 1731 9911
rect 1673 9871 1731 9877
rect 2317 9911 2375 9917
rect 2317 9877 2329 9911
rect 2363 9908 2375 9911
rect 3602 9908 3608 9920
rect 2363 9880 3608 9908
rect 2363 9877 2375 9880
rect 2317 9871 2375 9877
rect 3602 9868 3608 9880
rect 3660 9868 3666 9920
rect 17221 9911 17279 9917
rect 17221 9877 17233 9911
rect 17267 9908 17279 9911
rect 17494 9908 17500 9920
rect 17267 9880 17500 9908
rect 17267 9877 17279 9880
rect 17221 9871 17279 9877
rect 17494 9868 17500 9880
rect 17552 9868 17558 9920
rect 25038 9868 25044 9920
rect 25096 9908 25102 9920
rect 27448 9908 27476 10007
rect 25096 9880 27476 9908
rect 25096 9868 25102 9880
rect 27522 9868 27528 9920
rect 27580 9908 27586 9920
rect 27580 9880 27625 9908
rect 27580 9868 27586 9880
rect 1104 9818 28888 9840
rect 1104 9766 10214 9818
rect 10266 9766 10278 9818
rect 10330 9766 10342 9818
rect 10394 9766 10406 9818
rect 10458 9766 10470 9818
rect 10522 9766 19478 9818
rect 19530 9766 19542 9818
rect 19594 9766 19606 9818
rect 19658 9766 19670 9818
rect 19722 9766 19734 9818
rect 19786 9766 28888 9818
rect 1104 9744 28888 9766
rect 26234 9664 26240 9716
rect 26292 9704 26298 9716
rect 27157 9707 27215 9713
rect 27157 9704 27169 9707
rect 26292 9676 27169 9704
rect 26292 9664 26298 9676
rect 27157 9673 27169 9676
rect 27203 9673 27215 9707
rect 27157 9667 27215 9673
rect 3602 9636 3608 9648
rect 3563 9608 3608 9636
rect 3602 9596 3608 9608
rect 3660 9596 3666 9648
rect 6886 9608 27752 9636
rect 3786 9528 3792 9580
rect 3844 9568 3850 9580
rect 3844 9540 3889 9568
rect 3844 9528 3850 9540
rect 3234 9500 3240 9512
rect 3195 9472 3240 9500
rect 3234 9460 3240 9472
rect 3292 9460 3298 9512
rect 2958 9392 2964 9444
rect 3016 9432 3022 9444
rect 6886 9432 6914 9608
rect 26421 9571 26479 9577
rect 26421 9537 26433 9571
rect 26467 9568 26479 9571
rect 26510 9568 26516 9580
rect 26467 9540 26516 9568
rect 26467 9537 26479 9540
rect 26421 9531 26479 9537
rect 26510 9528 26516 9540
rect 26568 9528 26574 9580
rect 27724 9577 27752 9608
rect 27249 9571 27307 9577
rect 27249 9537 27261 9571
rect 27295 9537 27307 9571
rect 27249 9531 27307 9537
rect 27709 9571 27767 9577
rect 27709 9537 27721 9571
rect 27755 9537 27767 9571
rect 27709 9531 27767 9537
rect 24854 9500 24860 9512
rect 24815 9472 24860 9500
rect 24854 9460 24860 9472
rect 24912 9460 24918 9512
rect 25222 9460 25228 9512
rect 25280 9500 25286 9512
rect 26237 9503 26295 9509
rect 26237 9500 26249 9503
rect 25280 9472 26249 9500
rect 25280 9460 25286 9472
rect 26237 9469 26249 9472
rect 26283 9469 26295 9503
rect 27264 9500 27292 9531
rect 28258 9500 28264 9512
rect 27264 9472 28264 9500
rect 26237 9463 26295 9469
rect 28258 9460 28264 9472
rect 28316 9460 28322 9512
rect 27801 9435 27859 9441
rect 27801 9432 27813 9435
rect 3016 9404 6914 9432
rect 26206 9404 27813 9432
rect 3016 9392 3022 9404
rect 25498 9324 25504 9376
rect 25556 9364 25562 9376
rect 26206 9364 26234 9404
rect 27801 9401 27813 9404
rect 27847 9401 27859 9435
rect 27801 9395 27859 9401
rect 25556 9336 26234 9364
rect 25556 9324 25562 9336
rect 1104 9274 28888 9296
rect 1104 9222 5582 9274
rect 5634 9222 5646 9274
rect 5698 9222 5710 9274
rect 5762 9222 5774 9274
rect 5826 9222 5838 9274
rect 5890 9222 14846 9274
rect 14898 9222 14910 9274
rect 14962 9222 14974 9274
rect 15026 9222 15038 9274
rect 15090 9222 15102 9274
rect 15154 9222 24110 9274
rect 24162 9222 24174 9274
rect 24226 9222 24238 9274
rect 24290 9222 24302 9274
rect 24354 9222 24366 9274
rect 24418 9222 28888 9274
rect 1104 9200 28888 9222
rect 25222 9160 25228 9172
rect 25183 9132 25228 9160
rect 25222 9120 25228 9132
rect 25280 9120 25286 9172
rect 1394 9024 1400 9036
rect 1355 8996 1400 9024
rect 1394 8984 1400 8996
rect 1452 8984 1458 9036
rect 1578 9024 1584 9036
rect 1539 8996 1584 9024
rect 1578 8984 1584 8996
rect 1636 8984 1642 9036
rect 1854 9024 1860 9036
rect 1815 8996 1860 9024
rect 1854 8984 1860 8996
rect 1912 8984 1918 9036
rect 26326 9024 26332 9036
rect 26287 8996 26332 9024
rect 26326 8984 26332 8996
rect 26384 8984 26390 9036
rect 26513 9027 26571 9033
rect 26513 8993 26525 9027
rect 26559 9024 26571 9027
rect 27522 9024 27528 9036
rect 26559 8996 27528 9024
rect 26559 8993 26571 8996
rect 26513 8987 26571 8993
rect 27522 8984 27528 8996
rect 27580 8984 27586 9036
rect 24578 8916 24584 8968
rect 24636 8956 24642 8968
rect 24673 8959 24731 8965
rect 24673 8956 24685 8959
rect 24636 8928 24685 8956
rect 24636 8916 24642 8928
rect 24673 8925 24685 8928
rect 24719 8925 24731 8959
rect 24673 8919 24731 8925
rect 25038 8916 25044 8968
rect 25096 8956 25102 8968
rect 25133 8959 25191 8965
rect 25133 8956 25145 8959
rect 25096 8928 25145 8956
rect 25096 8916 25102 8928
rect 25133 8925 25145 8928
rect 25179 8925 25191 8959
rect 25133 8919 25191 8925
rect 28169 8891 28227 8897
rect 28169 8857 28181 8891
rect 28215 8888 28227 8891
rect 28994 8888 29000 8900
rect 28215 8860 29000 8888
rect 28215 8857 28227 8860
rect 28169 8851 28227 8857
rect 28994 8848 29000 8860
rect 29052 8848 29058 8900
rect 1104 8730 28888 8752
rect 1104 8678 10214 8730
rect 10266 8678 10278 8730
rect 10330 8678 10342 8730
rect 10394 8678 10406 8730
rect 10458 8678 10470 8730
rect 10522 8678 19478 8730
rect 19530 8678 19542 8730
rect 19594 8678 19606 8730
rect 19658 8678 19670 8730
rect 19722 8678 19734 8730
rect 19786 8678 28888 8730
rect 1104 8656 28888 8678
rect 27154 8440 27160 8492
rect 27212 8480 27218 8492
rect 27341 8483 27399 8489
rect 27341 8480 27353 8483
rect 27212 8452 27353 8480
rect 27212 8440 27218 8452
rect 27341 8449 27353 8452
rect 27387 8449 27399 8483
rect 27341 8443 27399 8449
rect 2958 8412 2964 8424
rect 2919 8384 2964 8412
rect 2958 8372 2964 8384
rect 3016 8372 3022 8424
rect 3142 8412 3148 8424
rect 3103 8384 3148 8412
rect 3142 8372 3148 8384
rect 3200 8372 3206 8424
rect 3421 8415 3479 8421
rect 3421 8381 3433 8415
rect 3467 8381 3479 8415
rect 25958 8412 25964 8424
rect 25919 8384 25964 8412
rect 3421 8375 3479 8381
rect 3436 8288 3464 8375
rect 25958 8372 25964 8384
rect 26016 8372 26022 8424
rect 26234 8372 26240 8424
rect 26292 8412 26298 8424
rect 26418 8412 26424 8424
rect 26292 8384 26337 8412
rect 26379 8384 26424 8412
rect 26292 8372 26298 8384
rect 26418 8372 26424 8384
rect 26476 8372 26482 8424
rect 27249 8347 27307 8353
rect 27249 8313 27261 8347
rect 27295 8344 27307 8347
rect 27890 8344 27896 8356
rect 27295 8316 27896 8344
rect 27295 8313 27307 8316
rect 27249 8307 27307 8313
rect 27890 8304 27896 8316
rect 27948 8304 27954 8356
rect 1486 8236 1492 8288
rect 1544 8276 1550 8288
rect 1581 8279 1639 8285
rect 1581 8276 1593 8279
rect 1544 8248 1593 8276
rect 1544 8236 1550 8248
rect 1581 8245 1593 8248
rect 1627 8245 1639 8279
rect 1581 8239 1639 8245
rect 3418 8236 3424 8288
rect 3476 8236 3482 8288
rect 27982 8276 27988 8288
rect 27943 8248 27988 8276
rect 27982 8236 27988 8248
rect 28040 8236 28046 8288
rect 1104 8186 28888 8208
rect 1104 8134 5582 8186
rect 5634 8134 5646 8186
rect 5698 8134 5710 8186
rect 5762 8134 5774 8186
rect 5826 8134 5838 8186
rect 5890 8134 14846 8186
rect 14898 8134 14910 8186
rect 14962 8134 14974 8186
rect 15026 8134 15038 8186
rect 15090 8134 15102 8186
rect 15154 8134 24110 8186
rect 24162 8134 24174 8186
rect 24226 8134 24238 8186
rect 24290 8134 24302 8186
rect 24354 8134 24366 8186
rect 24418 8134 28888 8186
rect 1104 8112 28888 8134
rect 1670 8032 1676 8084
rect 1728 8072 1734 8084
rect 1949 8075 2007 8081
rect 1949 8072 1961 8075
rect 1728 8044 1961 8072
rect 1728 8032 1734 8044
rect 1949 8041 1961 8044
rect 1995 8041 2007 8075
rect 2958 8072 2964 8084
rect 2919 8044 2964 8072
rect 1949 8035 2007 8041
rect 2958 8032 2964 8044
rect 3016 8032 3022 8084
rect 3142 8032 3148 8084
rect 3200 8072 3206 8084
rect 3881 8075 3939 8081
rect 3881 8072 3893 8075
rect 3200 8044 3893 8072
rect 3200 8032 3206 8044
rect 3881 8041 3893 8044
rect 3927 8041 3939 8075
rect 3881 8035 3939 8041
rect 25777 8075 25835 8081
rect 25777 8041 25789 8075
rect 25823 8072 25835 8075
rect 26234 8072 26240 8084
rect 25823 8044 26240 8072
rect 25823 8041 25835 8044
rect 25777 8035 25835 8041
rect 26234 8032 26240 8044
rect 26292 8032 26298 8084
rect 27522 7936 27528 7948
rect 27483 7908 27528 7936
rect 27522 7896 27528 7908
rect 27580 7896 27586 7948
rect 27982 7896 27988 7948
rect 28040 7936 28046 7948
rect 28169 7939 28227 7945
rect 28169 7936 28181 7939
rect 28040 7908 28181 7936
rect 28040 7896 28046 7908
rect 28169 7905 28181 7908
rect 28215 7905 28227 7939
rect 28169 7899 28227 7905
rect 2038 7868 2044 7880
rect 1999 7840 2044 7868
rect 2038 7828 2044 7840
rect 2096 7828 2102 7880
rect 3973 7871 4031 7877
rect 3973 7837 3985 7871
rect 4019 7837 4031 7871
rect 3973 7831 4031 7837
rect 4617 7871 4675 7877
rect 4617 7837 4629 7871
rect 4663 7868 4675 7871
rect 18690 7868 18696 7880
rect 4663 7840 18696 7868
rect 4663 7837 4675 7840
rect 4617 7831 4675 7837
rect 3988 7800 4016 7831
rect 18690 7828 18696 7840
rect 18748 7868 18754 7880
rect 25685 7871 25743 7877
rect 25685 7868 25697 7871
rect 18748 7840 25697 7868
rect 18748 7828 18754 7840
rect 25685 7837 25697 7840
rect 25731 7837 25743 7871
rect 25685 7831 25743 7837
rect 9214 7800 9220 7812
rect 3988 7772 9220 7800
rect 9214 7760 9220 7772
rect 9272 7760 9278 7812
rect 27890 7760 27896 7812
rect 27948 7800 27954 7812
rect 27985 7803 28043 7809
rect 27985 7800 27997 7803
rect 27948 7772 27997 7800
rect 27948 7760 27954 7772
rect 27985 7769 27997 7772
rect 28031 7769 28043 7803
rect 27985 7763 28043 7769
rect 3970 7692 3976 7744
rect 4028 7732 4034 7744
rect 4525 7735 4583 7741
rect 4525 7732 4537 7735
rect 4028 7704 4537 7732
rect 4028 7692 4034 7704
rect 4525 7701 4537 7704
rect 4571 7701 4583 7735
rect 4525 7695 4583 7701
rect 1104 7642 28888 7664
rect 1104 7590 10214 7642
rect 10266 7590 10278 7642
rect 10330 7590 10342 7642
rect 10394 7590 10406 7642
rect 10458 7590 10470 7642
rect 10522 7590 19478 7642
rect 19530 7590 19542 7642
rect 19594 7590 19606 7642
rect 19658 7590 19670 7642
rect 19722 7590 19734 7642
rect 19786 7590 28888 7642
rect 1104 7568 28888 7590
rect 3970 7460 3976 7472
rect 3931 7432 3976 7460
rect 3970 7420 3976 7432
rect 4028 7420 4034 7472
rect 24765 7463 24823 7469
rect 24765 7429 24777 7463
rect 24811 7460 24823 7463
rect 25498 7460 25504 7472
rect 24811 7432 25504 7460
rect 24811 7429 24823 7432
rect 24765 7423 24823 7429
rect 25498 7420 25504 7432
rect 25556 7420 25562 7472
rect 1486 7392 1492 7404
rect 1447 7364 1492 7392
rect 1486 7352 1492 7364
rect 1544 7352 1550 7404
rect 24578 7392 24584 7404
rect 24539 7364 24584 7392
rect 24578 7352 24584 7364
rect 24636 7352 24642 7404
rect 26418 7352 26424 7404
rect 26476 7392 26482 7404
rect 26973 7395 27031 7401
rect 26973 7392 26985 7395
rect 26476 7364 26985 7392
rect 26476 7352 26482 7364
rect 26973 7361 26985 7364
rect 27019 7361 27031 7395
rect 26973 7355 27031 7361
rect 1670 7324 1676 7336
rect 1631 7296 1676 7324
rect 1670 7284 1676 7296
rect 1728 7284 1734 7336
rect 2866 7324 2872 7336
rect 2827 7296 2872 7324
rect 2866 7284 2872 7296
rect 2924 7284 2930 7336
rect 3786 7324 3792 7336
rect 3747 7296 3792 7324
rect 3786 7284 3792 7296
rect 3844 7284 3850 7336
rect 4154 7284 4160 7336
rect 4212 7324 4218 7336
rect 4249 7327 4307 7333
rect 4249 7324 4261 7327
rect 4212 7296 4261 7324
rect 4212 7284 4218 7296
rect 4249 7293 4261 7296
rect 4295 7293 4307 7327
rect 26142 7324 26148 7336
rect 26103 7296 26148 7324
rect 4249 7287 4307 7293
rect 26142 7284 26148 7296
rect 26200 7284 26206 7336
rect 28077 7191 28135 7197
rect 28077 7157 28089 7191
rect 28123 7188 28135 7191
rect 28166 7188 28172 7200
rect 28123 7160 28172 7188
rect 28123 7157 28135 7160
rect 28077 7151 28135 7157
rect 28166 7148 28172 7160
rect 28224 7148 28230 7200
rect 1104 7098 28888 7120
rect 1104 7046 5582 7098
rect 5634 7046 5646 7098
rect 5698 7046 5710 7098
rect 5762 7046 5774 7098
rect 5826 7046 5838 7098
rect 5890 7046 14846 7098
rect 14898 7046 14910 7098
rect 14962 7046 14974 7098
rect 15026 7046 15038 7098
rect 15090 7046 15102 7098
rect 15154 7046 24110 7098
rect 24162 7046 24174 7098
rect 24226 7046 24238 7098
rect 24290 7046 24302 7098
rect 24354 7046 24366 7098
rect 24418 7046 28888 7098
rect 1104 7024 28888 7046
rect 1670 6944 1676 6996
rect 1728 6984 1734 6996
rect 1949 6987 2007 6993
rect 1949 6984 1961 6987
rect 1728 6956 1961 6984
rect 1728 6944 1734 6956
rect 1949 6953 1961 6956
rect 1995 6953 2007 6987
rect 3786 6984 3792 6996
rect 3747 6956 3792 6984
rect 1949 6947 2007 6953
rect 3786 6944 3792 6956
rect 3844 6944 3850 6996
rect 3418 6808 3424 6860
rect 3476 6848 3482 6860
rect 24854 6848 24860 6860
rect 3476 6820 24860 6848
rect 3476 6808 3482 6820
rect 24854 6808 24860 6820
rect 24912 6808 24918 6860
rect 27522 6848 27528 6860
rect 27483 6820 27528 6848
rect 27522 6808 27528 6820
rect 27580 6808 27586 6860
rect 28166 6848 28172 6860
rect 28127 6820 28172 6848
rect 28166 6808 28172 6820
rect 28224 6808 28230 6860
rect 2038 6780 2044 6792
rect 1999 6752 2044 6780
rect 2038 6740 2044 6752
rect 2096 6780 2102 6792
rect 6178 6780 6184 6792
rect 2096 6752 6184 6780
rect 2096 6740 2102 6752
rect 6178 6740 6184 6752
rect 6236 6740 6242 6792
rect 27798 6672 27804 6724
rect 27856 6712 27862 6724
rect 27985 6715 28043 6721
rect 27985 6712 27997 6715
rect 27856 6684 27997 6712
rect 27856 6672 27862 6684
rect 27985 6681 27997 6684
rect 28031 6681 28043 6715
rect 27985 6675 28043 6681
rect 1104 6554 28888 6576
rect 1104 6502 10214 6554
rect 10266 6502 10278 6554
rect 10330 6502 10342 6554
rect 10394 6502 10406 6554
rect 10458 6502 10470 6554
rect 10522 6502 19478 6554
rect 19530 6502 19542 6554
rect 19594 6502 19606 6554
rect 19658 6502 19670 6554
rect 19722 6502 19734 6554
rect 19786 6502 28888 6554
rect 1104 6480 28888 6502
rect 27798 6440 27804 6452
rect 27759 6412 27804 6440
rect 27798 6400 27804 6412
rect 27856 6400 27862 6452
rect 27614 6264 27620 6316
rect 27672 6304 27678 6316
rect 27709 6307 27767 6313
rect 27709 6304 27721 6307
rect 27672 6276 27721 6304
rect 27672 6264 27678 6276
rect 27709 6273 27721 6276
rect 27755 6273 27767 6307
rect 27709 6267 27767 6273
rect 1673 6239 1731 6245
rect 1673 6205 1685 6239
rect 1719 6236 1731 6239
rect 2133 6239 2191 6245
rect 2133 6236 2145 6239
rect 1719 6208 2145 6236
rect 1719 6205 1731 6208
rect 1673 6199 1731 6205
rect 2133 6205 2145 6208
rect 2179 6205 2191 6239
rect 2314 6236 2320 6248
rect 2275 6208 2320 6236
rect 2133 6199 2191 6205
rect 2314 6196 2320 6208
rect 2372 6196 2378 6248
rect 2590 6236 2596 6248
rect 2551 6208 2596 6236
rect 2590 6196 2596 6208
rect 2648 6196 2654 6248
rect 26326 6060 26332 6112
rect 26384 6100 26390 6112
rect 27065 6103 27123 6109
rect 27065 6100 27077 6103
rect 26384 6072 27077 6100
rect 26384 6060 26390 6072
rect 27065 6069 27077 6072
rect 27111 6069 27123 6103
rect 27065 6063 27123 6069
rect 1104 6010 28888 6032
rect 1104 5958 5582 6010
rect 5634 5958 5646 6010
rect 5698 5958 5710 6010
rect 5762 5958 5774 6010
rect 5826 5958 5838 6010
rect 5890 5958 14846 6010
rect 14898 5958 14910 6010
rect 14962 5958 14974 6010
rect 15026 5958 15038 6010
rect 15090 5958 15102 6010
rect 15154 5958 24110 6010
rect 24162 5958 24174 6010
rect 24226 5958 24238 6010
rect 24290 5958 24302 6010
rect 24354 5958 24366 6010
rect 24418 5958 28888 6010
rect 1104 5936 28888 5958
rect 2225 5899 2283 5905
rect 2225 5865 2237 5899
rect 2271 5896 2283 5899
rect 2314 5896 2320 5908
rect 2271 5868 2320 5896
rect 2271 5865 2283 5868
rect 2225 5859 2283 5865
rect 2314 5856 2320 5868
rect 2372 5856 2378 5908
rect 27614 5828 27620 5840
rect 22066 5800 27620 5828
rect 18417 5763 18475 5769
rect 18417 5760 18429 5763
rect 6886 5732 18429 5760
rect 2317 5695 2375 5701
rect 2317 5661 2329 5695
rect 2363 5692 2375 5695
rect 2961 5695 3019 5701
rect 2961 5692 2973 5695
rect 2363 5664 2973 5692
rect 2363 5661 2375 5664
rect 2317 5655 2375 5661
rect 2961 5661 2973 5664
rect 3007 5692 3019 5695
rect 6886 5692 6914 5732
rect 18417 5729 18429 5732
rect 18463 5760 18475 5763
rect 22066 5760 22094 5800
rect 27614 5788 27620 5800
rect 27672 5788 27678 5840
rect 26326 5760 26332 5772
rect 18463 5732 22094 5760
rect 26287 5732 26332 5760
rect 18463 5729 18475 5732
rect 18417 5723 18475 5729
rect 26326 5720 26332 5732
rect 26384 5720 26390 5772
rect 3007 5664 6914 5692
rect 18233 5695 18291 5701
rect 3007 5661 3019 5664
rect 2961 5655 3019 5661
rect 18233 5661 18245 5695
rect 18279 5692 18291 5695
rect 18598 5692 18604 5704
rect 18279 5664 18604 5692
rect 18279 5661 18291 5664
rect 18233 5655 18291 5661
rect 18598 5652 18604 5664
rect 18656 5692 18662 5704
rect 22738 5692 22744 5704
rect 18656 5664 22744 5692
rect 18656 5652 18662 5664
rect 22738 5652 22744 5664
rect 22796 5652 22802 5704
rect 26510 5624 26516 5636
rect 26471 5596 26516 5624
rect 26510 5584 26516 5596
rect 26568 5584 26574 5636
rect 28166 5624 28172 5636
rect 28127 5596 28172 5624
rect 28166 5584 28172 5596
rect 28224 5584 28230 5636
rect 2866 5556 2872 5568
rect 2827 5528 2872 5556
rect 2866 5516 2872 5528
rect 2924 5516 2930 5568
rect 1104 5466 28888 5488
rect 1104 5414 10214 5466
rect 10266 5414 10278 5466
rect 10330 5414 10342 5466
rect 10394 5414 10406 5466
rect 10458 5414 10470 5466
rect 10522 5414 19478 5466
rect 19530 5414 19542 5466
rect 19594 5414 19606 5466
rect 19658 5414 19670 5466
rect 19722 5414 19734 5466
rect 19786 5414 28888 5466
rect 1104 5392 28888 5414
rect 26510 5312 26516 5364
rect 26568 5352 26574 5364
rect 27525 5355 27583 5361
rect 27525 5352 27537 5355
rect 26568 5324 27537 5352
rect 26568 5312 26574 5324
rect 27525 5321 27537 5324
rect 27571 5321 27583 5355
rect 27525 5315 27583 5321
rect 2685 5287 2743 5293
rect 2685 5253 2697 5287
rect 2731 5284 2743 5287
rect 2866 5284 2872 5296
rect 2731 5256 2872 5284
rect 2731 5253 2743 5256
rect 2685 5247 2743 5253
rect 2866 5244 2872 5256
rect 2924 5244 2930 5296
rect 17865 5219 17923 5225
rect 17865 5185 17877 5219
rect 17911 5216 17923 5219
rect 18598 5216 18604 5228
rect 17911 5188 18604 5216
rect 17911 5185 17923 5188
rect 17865 5179 17923 5185
rect 18598 5176 18604 5188
rect 18656 5176 18662 5228
rect 22738 5216 22744 5228
rect 22699 5188 22744 5216
rect 22738 5176 22744 5188
rect 22796 5176 22802 5228
rect 27617 5219 27675 5225
rect 27617 5185 27629 5219
rect 27663 5216 27675 5219
rect 27890 5216 27896 5228
rect 27663 5188 27896 5216
rect 27663 5185 27675 5188
rect 27617 5179 27675 5185
rect 2041 5151 2099 5157
rect 2041 5117 2053 5151
rect 2087 5148 2099 5151
rect 2501 5151 2559 5157
rect 2501 5148 2513 5151
rect 2087 5120 2513 5148
rect 2087 5117 2099 5120
rect 2041 5111 2099 5117
rect 2501 5117 2513 5120
rect 2547 5117 2559 5151
rect 3142 5148 3148 5160
rect 3103 5120 3148 5148
rect 2501 5111 2559 5117
rect 3142 5108 3148 5120
rect 3200 5108 3206 5160
rect 19334 5108 19340 5160
rect 19392 5148 19398 5160
rect 27632 5148 27660 5179
rect 27890 5176 27896 5188
rect 27948 5176 27954 5228
rect 19392 5120 27660 5148
rect 19392 5108 19398 5120
rect 4985 5015 5043 5021
rect 4985 4981 4997 5015
rect 5031 5012 5043 5015
rect 6270 5012 6276 5024
rect 5031 4984 6276 5012
rect 5031 4981 5043 4984
rect 4985 4975 5043 4981
rect 6270 4972 6276 4984
rect 6328 4972 6334 5024
rect 17678 5012 17684 5024
rect 17639 4984 17684 5012
rect 17678 4972 17684 4984
rect 17736 4972 17742 5024
rect 22830 5012 22836 5024
rect 22791 4984 22836 5012
rect 22830 4972 22836 4984
rect 22888 4972 22894 5024
rect 1104 4922 28888 4944
rect 1104 4870 5582 4922
rect 5634 4870 5646 4922
rect 5698 4870 5710 4922
rect 5762 4870 5774 4922
rect 5826 4870 5838 4922
rect 5890 4870 14846 4922
rect 14898 4870 14910 4922
rect 14962 4870 14974 4922
rect 15026 4870 15038 4922
rect 15090 4870 15102 4922
rect 15154 4870 24110 4922
rect 24162 4870 24174 4922
rect 24226 4870 24238 4922
rect 24290 4870 24302 4922
rect 24354 4870 24366 4922
rect 24418 4870 28888 4922
rect 1104 4848 28888 4870
rect 2774 4632 2780 4684
rect 2832 4672 2838 4684
rect 3237 4675 3295 4681
rect 3237 4672 3249 4675
rect 2832 4644 3249 4672
rect 2832 4632 2838 4644
rect 3237 4641 3249 4644
rect 3283 4641 3295 4675
rect 3237 4635 3295 4641
rect 3326 4632 3332 4684
rect 3384 4672 3390 4684
rect 4433 4675 4491 4681
rect 4433 4672 4445 4675
rect 3384 4644 4445 4672
rect 3384 4632 3390 4644
rect 4433 4641 4445 4644
rect 4479 4641 4491 4675
rect 6270 4672 6276 4684
rect 6231 4644 6276 4672
rect 4433 4635 4491 4641
rect 6270 4632 6276 4644
rect 6328 4632 6334 4684
rect 21358 4672 21364 4684
rect 21319 4644 21364 4672
rect 21358 4632 21364 4644
rect 21416 4632 21422 4684
rect 27430 4672 27436 4684
rect 27391 4644 27436 4672
rect 27430 4632 27436 4644
rect 27488 4632 27494 4684
rect 27985 4675 28043 4681
rect 27985 4641 27997 4675
rect 28031 4672 28043 4675
rect 28534 4672 28540 4684
rect 28031 4644 28540 4672
rect 28031 4641 28043 4644
rect 27985 4635 28043 4641
rect 28534 4632 28540 4644
rect 28592 4632 28598 4684
rect 20714 4604 20720 4616
rect 20675 4576 20720 4604
rect 20714 4564 20720 4576
rect 20772 4564 20778 4616
rect 28166 4564 28172 4616
rect 28224 4604 28230 4616
rect 28224 4576 28269 4604
rect 28224 4564 28230 4576
rect 1394 4536 1400 4548
rect 1355 4508 1400 4536
rect 1394 4496 1400 4508
rect 1452 4496 1458 4548
rect 2958 4496 2964 4548
rect 3016 4536 3022 4548
rect 3053 4539 3111 4545
rect 3053 4536 3065 4539
rect 3016 4508 3065 4536
rect 3016 4496 3022 4508
rect 3053 4505 3065 4508
rect 3099 4505 3111 4539
rect 3053 4499 3111 4505
rect 6089 4539 6147 4545
rect 6089 4505 6101 4539
rect 6135 4536 6147 4539
rect 17678 4536 17684 4548
rect 6135 4508 17684 4536
rect 6135 4505 6147 4508
rect 6089 4499 6147 4505
rect 17678 4496 17684 4508
rect 17736 4496 17742 4548
rect 20898 4536 20904 4548
rect 20859 4508 20904 4536
rect 20898 4496 20904 4508
rect 20956 4496 20962 4548
rect 1104 4378 28888 4400
rect 1104 4326 10214 4378
rect 10266 4326 10278 4378
rect 10330 4326 10342 4378
rect 10394 4326 10406 4378
rect 10458 4326 10470 4378
rect 10522 4326 19478 4378
rect 19530 4326 19542 4378
rect 19594 4326 19606 4378
rect 19658 4326 19670 4378
rect 19722 4326 19734 4378
rect 19786 4326 28888 4378
rect 1104 4304 28888 4326
rect 20898 4264 20904 4276
rect 20859 4236 20904 4264
rect 20898 4224 20904 4236
rect 20956 4224 20962 4276
rect 19705 4199 19763 4205
rect 19705 4165 19717 4199
rect 19751 4196 19763 4199
rect 19751 4168 19932 4196
rect 19751 4165 19763 4168
rect 19705 4159 19763 4165
rect 1765 4131 1823 4137
rect 1765 4097 1777 4131
rect 1811 4128 1823 4131
rect 1946 4128 1952 4140
rect 1811 4100 1952 4128
rect 1811 4097 1823 4100
rect 1765 4091 1823 4097
rect 1946 4088 1952 4100
rect 2004 4088 2010 4140
rect 2409 4131 2467 4137
rect 2409 4097 2421 4131
rect 2455 4128 2467 4131
rect 2774 4128 2780 4140
rect 2455 4100 2780 4128
rect 2455 4097 2467 4100
rect 2409 4091 2467 4097
rect 2774 4088 2780 4100
rect 2832 4088 2838 4140
rect 5258 4128 5264 4140
rect 5219 4100 5264 4128
rect 5258 4088 5264 4100
rect 5316 4088 5322 4140
rect 9214 4128 9220 4140
rect 9127 4100 9220 4128
rect 9214 4088 9220 4100
rect 9272 4088 9278 4140
rect 10505 4131 10563 4137
rect 10505 4097 10517 4131
rect 10551 4128 10563 4131
rect 12894 4128 12900 4140
rect 10551 4100 12900 4128
rect 10551 4097 10563 4100
rect 10505 4091 10563 4097
rect 12894 4088 12900 4100
rect 12952 4088 12958 4140
rect 19904 4128 19932 4168
rect 20622 4128 20628 4140
rect 19904 4100 20628 4128
rect 20622 4088 20628 4100
rect 20680 4088 20686 4140
rect 20809 4131 20867 4137
rect 20809 4097 20821 4131
rect 20855 4128 20867 4131
rect 22738 4128 22744 4140
rect 20855 4100 22744 4128
rect 20855 4097 20867 4100
rect 20809 4091 20867 4097
rect 22738 4088 22744 4100
rect 22796 4088 22802 4140
rect 28077 4131 28135 4137
rect 28077 4097 28089 4131
rect 28123 4128 28135 4131
rect 28166 4128 28172 4140
rect 28123 4100 28172 4128
rect 28123 4097 28135 4100
rect 28077 4091 28135 4097
rect 28166 4088 28172 4100
rect 28224 4088 28230 4140
rect 2866 4060 2872 4072
rect 2827 4032 2872 4060
rect 2866 4020 2872 4032
rect 2924 4020 2930 4072
rect 3050 4060 3056 4072
rect 3011 4032 3056 4060
rect 3050 4020 3056 4032
rect 3108 4020 3114 4072
rect 3234 4020 3240 4072
rect 3292 4060 3298 4072
rect 3329 4063 3387 4069
rect 3329 4060 3341 4063
rect 3292 4032 3341 4060
rect 3292 4020 3298 4032
rect 3329 4029 3341 4032
rect 3375 4029 3387 4063
rect 3329 4023 3387 4029
rect 1673 3995 1731 4001
rect 1673 3961 1685 3995
rect 1719 3992 1731 3995
rect 2958 3992 2964 4004
rect 1719 3964 2964 3992
rect 1719 3961 1731 3964
rect 1673 3955 1731 3961
rect 2958 3952 2964 3964
rect 3016 3952 3022 4004
rect 9232 3992 9260 4088
rect 12618 4020 12624 4072
rect 12676 4060 12682 4072
rect 12989 4063 13047 4069
rect 12989 4060 13001 4063
rect 12676 4032 13001 4060
rect 12676 4020 12682 4032
rect 12989 4029 13001 4032
rect 13035 4029 13047 4063
rect 13170 4060 13176 4072
rect 13131 4032 13176 4060
rect 12989 4023 13047 4029
rect 13170 4020 13176 4032
rect 13228 4020 13234 4072
rect 13538 4060 13544 4072
rect 13499 4032 13544 4060
rect 13538 4020 13544 4032
rect 13596 4020 13602 4072
rect 18046 4060 18052 4072
rect 18007 4032 18052 4060
rect 18046 4020 18052 4032
rect 18104 4020 18110 4072
rect 18230 4020 18236 4072
rect 18288 4060 18294 4072
rect 19610 4060 19616 4072
rect 18288 4032 19616 4060
rect 18288 4020 18294 4032
rect 19610 4020 19616 4032
rect 19668 4020 19674 4072
rect 19886 4060 19892 4072
rect 19847 4032 19892 4060
rect 19886 4020 19892 4032
rect 19944 4020 19950 4072
rect 20714 4020 20720 4072
rect 20772 4060 20778 4072
rect 21821 4063 21879 4069
rect 21821 4060 21833 4063
rect 20772 4032 21833 4060
rect 20772 4020 20778 4032
rect 21821 4029 21833 4032
rect 21867 4029 21879 4063
rect 21821 4023 21879 4029
rect 26786 3992 26792 4004
rect 9232 3964 22094 3992
rect 5350 3924 5356 3936
rect 5311 3896 5356 3924
rect 5350 3884 5356 3896
rect 5408 3884 5414 3936
rect 6362 3924 6368 3936
rect 6323 3896 6368 3924
rect 6362 3884 6368 3896
rect 6420 3884 6426 3936
rect 7469 3927 7527 3933
rect 7469 3893 7481 3927
rect 7515 3924 7527 3927
rect 8662 3924 8668 3936
rect 7515 3896 8668 3924
rect 7515 3893 7527 3896
rect 7469 3887 7527 3893
rect 8662 3884 8668 3896
rect 8720 3884 8726 3936
rect 9306 3924 9312 3936
rect 9267 3896 9312 3924
rect 9306 3884 9312 3896
rect 9364 3884 9370 3936
rect 10597 3927 10655 3933
rect 10597 3893 10609 3927
rect 10643 3924 10655 3927
rect 11698 3924 11704 3936
rect 10643 3896 11704 3924
rect 10643 3893 10655 3896
rect 10597 3887 10655 3893
rect 11698 3884 11704 3896
rect 11756 3884 11762 3936
rect 12894 3884 12900 3936
rect 12952 3924 12958 3936
rect 19978 3924 19984 3936
rect 12952 3896 19984 3924
rect 12952 3884 12958 3896
rect 19978 3884 19984 3896
rect 20036 3884 20042 3936
rect 22066 3924 22094 3964
rect 26206 3964 26792 3992
rect 26206 3924 26234 3964
rect 26786 3952 26792 3964
rect 26844 3952 26850 4004
rect 26418 3924 26424 3936
rect 22066 3896 26234 3924
rect 26379 3896 26424 3924
rect 26418 3884 26424 3896
rect 26476 3884 26482 3936
rect 26970 3924 26976 3936
rect 26931 3896 26976 3924
rect 26970 3884 26976 3896
rect 27028 3884 27034 3936
rect 1104 3834 28888 3856
rect 1104 3782 5582 3834
rect 5634 3782 5646 3834
rect 5698 3782 5710 3834
rect 5762 3782 5774 3834
rect 5826 3782 5838 3834
rect 5890 3782 14846 3834
rect 14898 3782 14910 3834
rect 14962 3782 14974 3834
rect 15026 3782 15038 3834
rect 15090 3782 15102 3834
rect 15154 3782 24110 3834
rect 24162 3782 24174 3834
rect 24226 3782 24238 3834
rect 24290 3782 24302 3834
rect 24354 3782 24366 3834
rect 24418 3782 28888 3834
rect 1104 3760 28888 3782
rect 2869 3723 2927 3729
rect 2869 3689 2881 3723
rect 2915 3720 2927 3723
rect 3050 3720 3056 3732
rect 2915 3692 3056 3720
rect 2915 3689 2927 3692
rect 2869 3683 2927 3689
rect 3050 3680 3056 3692
rect 3108 3680 3114 3732
rect 5442 3680 5448 3732
rect 5500 3720 5506 3732
rect 12618 3720 12624 3732
rect 5500 3692 11836 3720
rect 12579 3692 12624 3720
rect 5500 3680 5506 3692
rect 11808 3652 11836 3692
rect 12618 3680 12624 3692
rect 12676 3680 12682 3732
rect 13170 3720 13176 3732
rect 13131 3692 13176 3720
rect 13170 3680 13176 3692
rect 13228 3680 13234 3732
rect 18325 3723 18383 3729
rect 18325 3689 18337 3723
rect 18371 3720 18383 3723
rect 19886 3720 19892 3732
rect 18371 3692 19892 3720
rect 18371 3689 18383 3692
rect 18325 3683 18383 3689
rect 19886 3680 19892 3692
rect 19944 3680 19950 3732
rect 4356 3624 11744 3652
rect 11808 3624 19564 3652
rect 4356 3584 4384 3624
rect 5350 3584 5356 3596
rect 2240 3556 4384 3584
rect 5311 3556 5356 3584
rect 1581 3519 1639 3525
rect 1581 3485 1593 3519
rect 1627 3516 1639 3519
rect 1670 3516 1676 3528
rect 1627 3488 1676 3516
rect 1627 3485 1639 3488
rect 1581 3479 1639 3485
rect 1670 3476 1676 3488
rect 1728 3476 1734 3528
rect 2240 3525 2268 3556
rect 2225 3519 2283 3525
rect 2225 3485 2237 3519
rect 2271 3485 2283 3519
rect 2774 3516 2780 3528
rect 2735 3488 2780 3516
rect 2225 3479 2283 3485
rect 2774 3476 2780 3488
rect 2832 3476 2838 3528
rect 4356 3525 4384 3556
rect 5350 3544 5356 3556
rect 5408 3544 5414 3596
rect 5902 3584 5908 3596
rect 5863 3556 5908 3584
rect 5902 3544 5908 3556
rect 5960 3544 5966 3596
rect 9306 3584 9312 3596
rect 9267 3556 9312 3584
rect 9306 3544 9312 3556
rect 9364 3544 9370 3596
rect 9674 3584 9680 3596
rect 9635 3556 9680 3584
rect 9674 3544 9680 3556
rect 9732 3544 9738 3596
rect 11716 3584 11744 3624
rect 19288 3584 19294 3596
rect 11716 3556 19294 3584
rect 19288 3544 19294 3556
rect 19346 3544 19352 3596
rect 4341 3519 4399 3525
rect 4341 3485 4353 3519
rect 4387 3485 4399 3519
rect 5166 3516 5172 3528
rect 5127 3488 5172 3516
rect 4341 3479 4399 3485
rect 5166 3476 5172 3488
rect 5224 3476 5230 3528
rect 7469 3519 7527 3525
rect 7469 3516 7481 3519
rect 6886 3488 7481 3516
rect 2792 3448 2820 3476
rect 6886 3448 6914 3488
rect 7469 3485 7481 3488
rect 7515 3485 7527 3519
rect 7469 3479 7527 3485
rect 8389 3519 8447 3525
rect 8389 3485 8401 3519
rect 8435 3516 8447 3519
rect 9125 3519 9183 3525
rect 9125 3516 9137 3519
rect 8435 3488 9137 3516
rect 8435 3485 8447 3488
rect 8389 3479 8447 3485
rect 9125 3485 9137 3488
rect 9171 3485 9183 3519
rect 9125 3479 9183 3485
rect 11514 3476 11520 3528
rect 11572 3516 11578 3528
rect 11609 3519 11667 3525
rect 11609 3516 11621 3519
rect 11572 3488 11621 3516
rect 11572 3476 11578 3488
rect 11609 3485 11621 3488
rect 11655 3485 11667 3519
rect 13078 3516 13084 3528
rect 13039 3488 13084 3516
rect 11609 3479 11667 3485
rect 13078 3476 13084 3488
rect 13136 3476 13142 3528
rect 14642 3516 14648 3528
rect 14603 3488 14648 3516
rect 14642 3476 14648 3488
rect 14700 3476 14706 3528
rect 15105 3519 15163 3525
rect 15105 3485 15117 3519
rect 15151 3485 15163 3519
rect 16298 3516 16304 3528
rect 16259 3488 16304 3516
rect 15105 3479 15163 3485
rect 2792 3420 6914 3448
rect 14274 3408 14280 3460
rect 14332 3448 14338 3460
rect 15120 3448 15148 3479
rect 16298 3476 16304 3488
rect 16356 3476 16362 3528
rect 16666 3476 16672 3528
rect 16724 3516 16730 3528
rect 19536 3525 19564 3624
rect 20622 3612 20628 3664
rect 20680 3652 20686 3664
rect 25409 3655 25467 3661
rect 25409 3652 25421 3655
rect 20680 3624 25421 3652
rect 20680 3612 20686 3624
rect 25409 3621 25421 3624
rect 25455 3621 25467 3655
rect 28442 3652 28448 3664
rect 25409 3615 25467 3621
rect 26206 3624 28448 3652
rect 21910 3584 21916 3596
rect 21871 3556 21916 3584
rect 21910 3544 21916 3556
rect 21968 3544 21974 3596
rect 16945 3519 17003 3525
rect 16945 3516 16957 3519
rect 16724 3488 16957 3516
rect 16724 3476 16730 3488
rect 16945 3485 16957 3488
rect 16991 3485 17003 3519
rect 16945 3479 17003 3485
rect 19521 3519 19579 3525
rect 19521 3485 19533 3519
rect 19567 3485 19579 3519
rect 19521 3479 19579 3485
rect 14332 3420 15148 3448
rect 19536 3448 19564 3479
rect 19610 3476 19616 3528
rect 19668 3516 19674 3528
rect 20625 3519 20683 3525
rect 20625 3516 20637 3519
rect 19668 3488 20637 3516
rect 19668 3476 19674 3488
rect 20625 3485 20637 3488
rect 20671 3485 20683 3519
rect 21266 3516 21272 3528
rect 21227 3488 21272 3516
rect 20625 3479 20683 3485
rect 21266 3476 21272 3488
rect 21324 3476 21330 3528
rect 24026 3476 24032 3528
rect 24084 3516 24090 3528
rect 24397 3519 24455 3525
rect 24397 3516 24409 3519
rect 24084 3488 24409 3516
rect 24084 3476 24090 3488
rect 24397 3485 24409 3488
rect 24443 3485 24455 3519
rect 24397 3479 24455 3485
rect 25501 3519 25559 3525
rect 25501 3485 25513 3519
rect 25547 3516 25559 3519
rect 26206 3516 26234 3624
rect 28442 3612 28448 3624
rect 28500 3612 28506 3664
rect 26329 3587 26387 3593
rect 26329 3553 26341 3587
rect 26375 3584 26387 3587
rect 26970 3584 26976 3596
rect 26375 3556 26976 3584
rect 26375 3553 26387 3556
rect 26329 3547 26387 3553
rect 26970 3544 26976 3556
rect 27028 3544 27034 3596
rect 27522 3584 27528 3596
rect 27483 3556 27528 3584
rect 27522 3544 27528 3556
rect 27580 3544 27586 3596
rect 25547 3488 26234 3516
rect 25547 3485 25559 3488
rect 25501 3479 25559 3485
rect 20717 3451 20775 3457
rect 19536 3420 19748 3448
rect 14332 3408 14338 3420
rect 1854 3340 1860 3392
rect 1912 3380 1918 3392
rect 2133 3383 2191 3389
rect 2133 3380 2145 3383
rect 1912 3352 2145 3380
rect 1912 3340 1918 3352
rect 2133 3349 2145 3352
rect 2179 3349 2191 3383
rect 2133 3343 2191 3349
rect 4154 3340 4160 3392
rect 4212 3380 4218 3392
rect 4249 3383 4307 3389
rect 4249 3380 4261 3383
rect 4212 3352 4261 3380
rect 4212 3340 4218 3352
rect 4249 3349 4261 3352
rect 4295 3349 4307 3383
rect 4249 3343 4307 3349
rect 7561 3383 7619 3389
rect 7561 3349 7573 3383
rect 7607 3380 7619 3383
rect 8846 3380 8852 3392
rect 7607 3352 8852 3380
rect 7607 3349 7619 3352
rect 7561 3343 7619 3349
rect 8846 3340 8852 3352
rect 8904 3340 8910 3392
rect 14458 3340 14464 3392
rect 14516 3380 14522 3392
rect 14553 3383 14611 3389
rect 14553 3380 14565 3383
rect 14516 3352 14565 3380
rect 14516 3340 14522 3352
rect 14553 3349 14565 3352
rect 14599 3349 14611 3383
rect 14553 3343 14611 3349
rect 16393 3383 16451 3389
rect 16393 3349 16405 3383
rect 16439 3380 16451 3383
rect 16850 3380 16856 3392
rect 16439 3352 16856 3380
rect 16439 3349 16451 3352
rect 16393 3343 16451 3349
rect 16850 3340 16856 3352
rect 16908 3340 16914 3392
rect 19334 3340 19340 3392
rect 19392 3380 19398 3392
rect 19613 3383 19671 3389
rect 19613 3380 19625 3383
rect 19392 3352 19625 3380
rect 19392 3340 19398 3352
rect 19613 3349 19625 3352
rect 19659 3349 19671 3383
rect 19720 3380 19748 3420
rect 20717 3417 20729 3451
rect 20763 3448 20775 3451
rect 21453 3451 21511 3457
rect 21453 3448 21465 3451
rect 20763 3420 21465 3448
rect 20763 3417 20775 3420
rect 20717 3411 20775 3417
rect 21453 3417 21465 3420
rect 21499 3417 21511 3451
rect 21453 3411 21511 3417
rect 26513 3451 26571 3457
rect 26513 3417 26525 3451
rect 26559 3448 26571 3451
rect 27062 3448 27068 3460
rect 26559 3420 27068 3448
rect 26559 3417 26571 3420
rect 26513 3411 26571 3417
rect 27062 3408 27068 3420
rect 27120 3408 27126 3460
rect 26970 3380 26976 3392
rect 19720 3352 26976 3380
rect 19613 3343 19671 3349
rect 26970 3340 26976 3352
rect 27028 3340 27034 3392
rect 1104 3290 28888 3312
rect 1104 3238 10214 3290
rect 10266 3238 10278 3290
rect 10330 3238 10342 3290
rect 10394 3238 10406 3290
rect 10458 3238 10470 3290
rect 10522 3238 19478 3290
rect 19530 3238 19542 3290
rect 19594 3238 19606 3290
rect 19658 3238 19670 3290
rect 19722 3238 19734 3290
rect 19786 3238 28888 3290
rect 1104 3216 28888 3238
rect 658 3136 664 3188
rect 716 3176 722 3188
rect 2590 3176 2596 3188
rect 716 3148 2596 3176
rect 716 3136 722 3148
rect 2590 3136 2596 3148
rect 2648 3136 2654 3188
rect 13078 3176 13084 3188
rect 2700 3148 13084 3176
rect 1854 3108 1860 3120
rect 1815 3080 1860 3108
rect 1854 3068 1860 3080
rect 1912 3068 1918 3120
rect 1946 3068 1952 3120
rect 2004 3108 2010 3120
rect 2700 3108 2728 3148
rect 13078 3136 13084 3148
rect 13136 3136 13142 3188
rect 19978 3136 19984 3188
rect 20036 3176 20042 3188
rect 27062 3176 27068 3188
rect 20036 3148 26234 3176
rect 27023 3148 27068 3176
rect 20036 3136 20042 3148
rect 4154 3108 4160 3120
rect 2004 3080 2728 3108
rect 4115 3080 4160 3108
rect 2004 3068 2010 3080
rect 4154 3068 4160 3080
rect 4212 3068 4218 3120
rect 8846 3108 8852 3120
rect 8807 3080 8852 3108
rect 8846 3068 8852 3080
rect 8904 3068 8910 3120
rect 11698 3108 11704 3120
rect 11659 3080 11704 3108
rect 11698 3068 11704 3080
rect 11756 3068 11762 3120
rect 14458 3108 14464 3120
rect 14419 3080 14464 3108
rect 14458 3068 14464 3080
rect 14516 3068 14522 3120
rect 16850 3108 16856 3120
rect 16811 3080 16856 3108
rect 16850 3068 16856 3080
rect 16908 3068 16914 3120
rect 19334 3068 19340 3120
rect 19392 3108 19398 3120
rect 19613 3111 19671 3117
rect 19613 3108 19625 3111
rect 19392 3080 19625 3108
rect 19392 3068 19398 3080
rect 19613 3077 19625 3080
rect 19659 3077 19671 3111
rect 19613 3071 19671 3077
rect 23477 3111 23535 3117
rect 23477 3077 23489 3111
rect 23523 3108 23535 3111
rect 24213 3111 24271 3117
rect 24213 3108 24225 3111
rect 23523 3080 24225 3108
rect 23523 3077 23535 3080
rect 23477 3071 23535 3077
rect 24213 3077 24225 3080
rect 24259 3077 24271 3111
rect 26206 3108 26234 3148
rect 27062 3136 27068 3148
rect 27120 3136 27126 3188
rect 28074 3108 28080 3120
rect 26206 3080 28080 3108
rect 24213 3071 24271 3077
rect 28074 3068 28080 3080
rect 28132 3068 28138 3120
rect 1670 3040 1676 3052
rect 1631 3012 1676 3040
rect 1670 3000 1676 3012
rect 1728 3000 1734 3052
rect 6362 3040 6368 3052
rect 6323 3012 6368 3040
rect 6362 3000 6368 3012
rect 6420 3000 6426 3052
rect 8662 3040 8668 3052
rect 8623 3012 8668 3040
rect 8662 3000 8668 3012
rect 8720 3000 8726 3052
rect 11514 3040 11520 3052
rect 11475 3012 11520 3040
rect 11514 3000 11520 3012
rect 11572 3000 11578 3052
rect 14274 3040 14280 3052
rect 14235 3012 14280 3040
rect 14274 3000 14280 3012
rect 14332 3000 14338 3052
rect 16666 3040 16672 3052
rect 16627 3012 16672 3040
rect 16666 3000 16672 3012
rect 16724 3000 16730 3052
rect 21266 3000 21272 3052
rect 21324 3040 21330 3052
rect 21821 3043 21879 3049
rect 21821 3040 21833 3043
rect 21324 3012 21833 3040
rect 21324 3000 21330 3012
rect 21821 3009 21833 3012
rect 21867 3009 21879 3043
rect 22830 3040 22836 3052
rect 21821 3003 21879 3009
rect 22066 3012 22836 3040
rect 2774 2972 2780 2984
rect 2735 2944 2780 2972
rect 2774 2932 2780 2944
rect 2832 2932 2838 2984
rect 3970 2972 3976 2984
rect 3931 2944 3976 2972
rect 3970 2932 3976 2944
rect 4028 2932 4034 2984
rect 4522 2972 4528 2984
rect 4483 2944 4528 2972
rect 4522 2932 4528 2944
rect 4580 2932 4586 2984
rect 6546 2972 6552 2984
rect 6507 2944 6552 2972
rect 6546 2932 6552 2944
rect 6604 2932 6610 2984
rect 6825 2975 6883 2981
rect 6825 2941 6837 2975
rect 6871 2941 6883 2975
rect 6825 2935 6883 2941
rect 6454 2864 6460 2916
rect 6512 2904 6518 2916
rect 6840 2904 6868 2935
rect 8386 2932 8392 2984
rect 8444 2972 8450 2984
rect 9125 2975 9183 2981
rect 9125 2972 9137 2975
rect 8444 2944 9137 2972
rect 8444 2932 8450 2944
rect 9125 2941 9137 2944
rect 9171 2941 9183 2975
rect 9125 2935 9183 2941
rect 11977 2975 12035 2981
rect 11977 2941 11989 2975
rect 12023 2941 12035 2975
rect 14734 2972 14740 2984
rect 14695 2944 14740 2972
rect 11977 2935 12035 2941
rect 6512 2876 6868 2904
rect 6512 2864 6518 2876
rect 10962 2864 10968 2916
rect 11020 2904 11026 2916
rect 11992 2904 12020 2935
rect 14734 2932 14740 2944
rect 14792 2932 14798 2984
rect 17129 2975 17187 2981
rect 17129 2972 17141 2975
rect 16776 2944 17141 2972
rect 16776 2916 16804 2944
rect 17129 2941 17141 2944
rect 17175 2941 17187 2975
rect 19426 2972 19432 2984
rect 19387 2944 19432 2972
rect 17129 2935 17187 2941
rect 19426 2932 19432 2944
rect 19484 2932 19490 2984
rect 19978 2972 19984 2984
rect 19939 2944 19984 2972
rect 19978 2932 19984 2944
rect 20036 2932 20042 2984
rect 11020 2876 12020 2904
rect 11020 2864 11026 2876
rect 16758 2864 16764 2916
rect 16816 2864 16822 2916
rect 2590 2796 2596 2848
rect 2648 2836 2654 2848
rect 3142 2836 3148 2848
rect 2648 2808 3148 2836
rect 2648 2796 2654 2808
rect 3142 2796 3148 2808
rect 3200 2796 3206 2848
rect 16022 2796 16028 2848
rect 16080 2836 16086 2848
rect 16298 2836 16304 2848
rect 16080 2808 16304 2836
rect 16080 2796 16086 2808
rect 16298 2796 16304 2808
rect 16356 2836 16362 2848
rect 22066 2836 22094 3012
rect 22830 3000 22836 3012
rect 22888 3040 22894 3052
rect 23385 3043 23443 3049
rect 23385 3040 23397 3043
rect 22888 3012 23397 3040
rect 22888 3000 22894 3012
rect 23385 3009 23397 3012
rect 23431 3009 23443 3043
rect 24026 3040 24032 3052
rect 23987 3012 24032 3040
rect 23385 3003 23443 3009
rect 24026 3000 24032 3012
rect 24084 3000 24090 3052
rect 26970 3040 26976 3052
rect 26931 3012 26976 3040
rect 26970 3000 26976 3012
rect 27028 3000 27034 3052
rect 27706 3000 27712 3052
rect 27764 3040 27770 3052
rect 27801 3043 27859 3049
rect 27801 3040 27813 3043
rect 27764 3012 27813 3040
rect 27764 3000 27770 3012
rect 27801 3009 27813 3012
rect 27847 3009 27859 3043
rect 27801 3003 27859 3009
rect 25130 2972 25136 2984
rect 25091 2944 25136 2972
rect 25130 2932 25136 2944
rect 25188 2932 25194 2984
rect 16356 2808 22094 2836
rect 16356 2796 16362 2808
rect 26234 2796 26240 2848
rect 26292 2836 26298 2848
rect 27709 2839 27767 2845
rect 27709 2836 27721 2839
rect 26292 2808 27721 2836
rect 26292 2796 26298 2808
rect 27709 2805 27721 2808
rect 27755 2805 27767 2839
rect 27709 2799 27767 2805
rect 1104 2746 28888 2768
rect 1104 2694 5582 2746
rect 5634 2694 5646 2746
rect 5698 2694 5710 2746
rect 5762 2694 5774 2746
rect 5826 2694 5838 2746
rect 5890 2694 14846 2746
rect 14898 2694 14910 2746
rect 14962 2694 14974 2746
rect 15026 2694 15038 2746
rect 15090 2694 15102 2746
rect 15154 2694 24110 2746
rect 24162 2694 24174 2746
rect 24226 2694 24238 2746
rect 24290 2694 24302 2746
rect 24354 2694 24366 2746
rect 24418 2694 28888 2746
rect 1104 2672 28888 2694
rect 2866 2632 2872 2644
rect 2827 2604 2872 2632
rect 2866 2592 2872 2604
rect 2924 2592 2930 2644
rect 3970 2592 3976 2644
rect 4028 2632 4034 2644
rect 4065 2635 4123 2641
rect 4065 2632 4077 2635
rect 4028 2604 4077 2632
rect 4028 2592 4034 2604
rect 4065 2601 4077 2604
rect 4111 2601 4123 2635
rect 4065 2595 4123 2601
rect 5166 2592 5172 2644
rect 5224 2632 5230 2644
rect 5261 2635 5319 2641
rect 5261 2632 5273 2635
rect 5224 2604 5273 2632
rect 5224 2592 5230 2604
rect 5261 2601 5273 2604
rect 5307 2601 5319 2635
rect 5261 2595 5319 2601
rect 6457 2635 6515 2641
rect 6457 2601 6469 2635
rect 6503 2632 6515 2635
rect 6546 2632 6552 2644
rect 6503 2604 6552 2632
rect 6503 2601 6515 2604
rect 6457 2595 6515 2601
rect 6546 2592 6552 2604
rect 6604 2592 6610 2644
rect 9490 2632 9496 2644
rect 9451 2604 9496 2632
rect 9490 2592 9496 2604
rect 9548 2592 9554 2644
rect 16850 2632 16856 2644
rect 16811 2604 16856 2632
rect 16850 2592 16856 2604
rect 16908 2592 16914 2644
rect 17494 2632 17500 2644
rect 17455 2604 17500 2632
rect 17494 2592 17500 2604
rect 17552 2592 17558 2644
rect 19426 2632 19432 2644
rect 19387 2604 19432 2632
rect 19426 2592 19432 2604
rect 19484 2592 19490 2644
rect 20438 2592 20444 2644
rect 20496 2632 20502 2644
rect 20496 2604 27476 2632
rect 20496 2592 20502 2604
rect 3418 2524 3424 2576
rect 3476 2564 3482 2576
rect 25314 2564 25320 2576
rect 3476 2536 25320 2564
rect 3476 2524 3482 2536
rect 25314 2524 25320 2536
rect 25372 2524 25378 2576
rect 25958 2496 25964 2508
rect 25919 2468 25964 2496
rect 25958 2456 25964 2468
rect 26016 2456 26022 2508
rect 26234 2456 26240 2508
rect 26292 2496 26298 2508
rect 26418 2496 26424 2508
rect 26292 2468 26337 2496
rect 26379 2468 26424 2496
rect 26292 2456 26298 2468
rect 26418 2456 26424 2468
rect 26476 2456 26482 2508
rect 27448 2505 27476 2604
rect 27433 2499 27491 2505
rect 27433 2465 27445 2499
rect 27479 2465 27491 2499
rect 27433 2459 27491 2465
rect 6178 2388 6184 2440
rect 6236 2428 6242 2440
rect 6365 2431 6423 2437
rect 6365 2428 6377 2431
rect 6236 2400 6377 2428
rect 6236 2388 6242 2400
rect 6365 2397 6377 2400
rect 6411 2428 6423 2431
rect 16022 2428 16028 2440
rect 6411 2400 16028 2428
rect 6411 2397 6423 2400
rect 6365 2391 6423 2397
rect 16022 2388 16028 2400
rect 16080 2388 16086 2440
rect 16114 2388 16120 2440
rect 16172 2428 16178 2440
rect 16669 2431 16727 2437
rect 16669 2428 16681 2431
rect 16172 2400 16681 2428
rect 16172 2388 16178 2400
rect 16669 2397 16681 2400
rect 16715 2397 16727 2431
rect 16669 2391 16727 2397
rect 17402 2388 17408 2440
rect 17460 2428 17466 2440
rect 17681 2431 17739 2437
rect 17681 2428 17693 2431
rect 17460 2400 17693 2428
rect 17460 2388 17466 2400
rect 17681 2397 17693 2400
rect 17727 2397 17739 2431
rect 17681 2391 17739 2397
rect 27062 2388 27068 2440
rect 27120 2428 27126 2440
rect 27157 2431 27215 2437
rect 27157 2428 27169 2431
rect 27120 2400 27169 2428
rect 27120 2388 27126 2400
rect 27157 2397 27169 2400
rect 27203 2397 27215 2431
rect 27157 2391 27215 2397
rect 9030 2320 9036 2372
rect 9088 2360 9094 2372
rect 9401 2363 9459 2369
rect 9401 2360 9413 2363
rect 9088 2332 9413 2360
rect 9088 2320 9094 2332
rect 9401 2329 9413 2332
rect 9447 2329 9459 2363
rect 9401 2323 9459 2329
rect 1104 2202 28888 2224
rect 1104 2150 10214 2202
rect 10266 2150 10278 2202
rect 10330 2150 10342 2202
rect 10394 2150 10406 2202
rect 10458 2150 10470 2202
rect 10522 2150 19478 2202
rect 19530 2150 19542 2202
rect 19594 2150 19606 2202
rect 19658 2150 19670 2202
rect 19722 2150 19734 2202
rect 19786 2150 28888 2202
rect 1104 2128 28888 2150
<< via1 >>
rect 5582 47302 5634 47354
rect 5646 47302 5698 47354
rect 5710 47302 5762 47354
rect 5774 47302 5826 47354
rect 5838 47302 5890 47354
rect 14846 47302 14898 47354
rect 14910 47302 14962 47354
rect 14974 47302 15026 47354
rect 15038 47302 15090 47354
rect 15102 47302 15154 47354
rect 24110 47302 24162 47354
rect 24174 47302 24226 47354
rect 24238 47302 24290 47354
rect 24302 47302 24354 47354
rect 24366 47302 24418 47354
rect 23204 47107 23256 47116
rect 23204 47073 23213 47107
rect 23213 47073 23247 47107
rect 23247 47073 23256 47107
rect 23204 47064 23256 47073
rect 28356 47064 28408 47116
rect 1676 46996 1728 47048
rect 3608 46996 3660 47048
rect 3792 47039 3844 47048
rect 3792 47005 3801 47039
rect 3801 47005 3835 47039
rect 3835 47005 3844 47039
rect 3792 46996 3844 47005
rect 6092 46996 6144 47048
rect 2596 46860 2648 46912
rect 3056 46860 3108 46912
rect 6552 46903 6604 46912
rect 6552 46869 6561 46903
rect 6561 46869 6595 46903
rect 6595 46869 6604 46903
rect 6552 46860 6604 46869
rect 6644 46860 6696 46912
rect 7840 47039 7892 47048
rect 7840 47005 7849 47039
rect 7849 47005 7883 47039
rect 7883 47005 7892 47039
rect 7840 46996 7892 47005
rect 13820 46996 13872 47048
rect 16672 47039 16724 47048
rect 16672 47005 16681 47039
rect 16681 47005 16715 47039
rect 16715 47005 16724 47039
rect 16672 46996 16724 47005
rect 18144 47039 18196 47048
rect 18144 47005 18153 47039
rect 18153 47005 18187 47039
rect 18187 47005 18196 47039
rect 18144 46996 18196 47005
rect 19340 46996 19392 47048
rect 21916 46996 21968 47048
rect 28172 46996 28224 47048
rect 22744 46928 22796 46980
rect 26240 46971 26292 46980
rect 26240 46937 26249 46971
rect 26249 46937 26283 46971
rect 26283 46937 26292 46971
rect 26240 46928 26292 46937
rect 7288 46903 7340 46912
rect 7288 46869 7297 46903
rect 7297 46869 7331 46903
rect 7331 46869 7340 46903
rect 7288 46860 7340 46869
rect 11612 46860 11664 46912
rect 12532 46860 12584 46912
rect 27068 46860 27120 46912
rect 28080 46860 28132 46912
rect 10214 46758 10266 46810
rect 10278 46758 10330 46810
rect 10342 46758 10394 46810
rect 10406 46758 10458 46810
rect 10470 46758 10522 46810
rect 19478 46758 19530 46810
rect 19542 46758 19594 46810
rect 19606 46758 19658 46810
rect 19670 46758 19722 46810
rect 19734 46758 19786 46810
rect 23848 46656 23900 46708
rect 26240 46656 26292 46708
rect 25596 46631 25648 46640
rect 25596 46597 25605 46631
rect 25605 46597 25639 46631
rect 25639 46597 25648 46631
rect 25596 46588 25648 46597
rect 1676 46563 1728 46572
rect 1676 46529 1685 46563
rect 1685 46529 1719 46563
rect 1719 46529 1728 46563
rect 1676 46520 1728 46529
rect 3608 46520 3660 46572
rect 7840 46563 7892 46572
rect 7840 46529 7849 46563
rect 7849 46529 7883 46563
rect 7883 46529 7892 46563
rect 7840 46520 7892 46529
rect 13820 46563 13872 46572
rect 13820 46529 13829 46563
rect 13829 46529 13863 46563
rect 13863 46529 13872 46563
rect 13820 46520 13872 46529
rect 16672 46563 16724 46572
rect 16672 46529 16681 46563
rect 16681 46529 16715 46563
rect 16715 46529 16724 46563
rect 16672 46520 16724 46529
rect 19340 46520 19392 46572
rect 26976 46563 27028 46572
rect 26976 46529 26985 46563
rect 26985 46529 27019 46563
rect 27019 46529 27028 46563
rect 26976 46520 27028 46529
rect 2136 46452 2188 46504
rect 4160 46495 4212 46504
rect 1308 46384 1360 46436
rect 4160 46461 4169 46495
rect 4169 46461 4203 46495
rect 4203 46461 4212 46495
rect 4160 46452 4212 46461
rect 8024 46495 8076 46504
rect 2320 46384 2372 46436
rect 8024 46461 8033 46495
rect 8033 46461 8067 46495
rect 8067 46461 8076 46495
rect 8024 46452 8076 46461
rect 8392 46495 8444 46504
rect 8392 46461 8401 46495
rect 8401 46461 8435 46495
rect 8435 46461 8444 46495
rect 8392 46452 8444 46461
rect 11704 46495 11756 46504
rect 11704 46461 11713 46495
rect 11713 46461 11747 46495
rect 11747 46461 11756 46495
rect 11704 46452 11756 46461
rect 13452 46452 13504 46504
rect 16856 46495 16908 46504
rect 13544 46384 13596 46436
rect 16856 46461 16865 46495
rect 16865 46461 16899 46495
rect 16899 46461 16908 46495
rect 16856 46452 16908 46461
rect 16764 46384 16816 46436
rect 19984 46495 20036 46504
rect 19984 46461 19993 46495
rect 19993 46461 20027 46495
rect 20027 46461 20036 46495
rect 19984 46452 20036 46461
rect 23756 46495 23808 46504
rect 23756 46461 23765 46495
rect 23765 46461 23799 46495
rect 23799 46461 23808 46495
rect 23756 46452 23808 46461
rect 23940 46495 23992 46504
rect 23940 46461 23949 46495
rect 23949 46461 23983 46495
rect 23983 46461 23992 46495
rect 23940 46452 23992 46461
rect 19340 46384 19392 46436
rect 9588 46316 9640 46368
rect 10968 46316 11020 46368
rect 17592 46316 17644 46368
rect 22008 46316 22060 46368
rect 26424 46316 26476 46368
rect 27896 46359 27948 46368
rect 27896 46325 27905 46359
rect 27905 46325 27939 46359
rect 27939 46325 27948 46359
rect 27896 46316 27948 46325
rect 5582 46214 5634 46266
rect 5646 46214 5698 46266
rect 5710 46214 5762 46266
rect 5774 46214 5826 46266
rect 5838 46214 5890 46266
rect 14846 46214 14898 46266
rect 14910 46214 14962 46266
rect 14974 46214 15026 46266
rect 15038 46214 15090 46266
rect 15102 46214 15154 46266
rect 24110 46214 24162 46266
rect 24174 46214 24226 46266
rect 24238 46214 24290 46266
rect 24302 46214 24354 46266
rect 24366 46214 24418 46266
rect 2136 46155 2188 46164
rect 2136 46121 2145 46155
rect 2145 46121 2179 46155
rect 2179 46121 2188 46155
rect 2136 46112 2188 46121
rect 4160 46112 4212 46164
rect 8024 46155 8076 46164
rect 8024 46121 8033 46155
rect 8033 46121 8067 46155
rect 8067 46121 8076 46155
rect 8024 46112 8076 46121
rect 13452 46155 13504 46164
rect 13452 46121 13461 46155
rect 13461 46121 13495 46155
rect 13495 46121 13504 46155
rect 13452 46112 13504 46121
rect 16856 46112 16908 46164
rect 23756 46112 23808 46164
rect 1584 45951 1636 45960
rect 1584 45917 1593 45951
rect 1593 45917 1627 45951
rect 1627 45917 1636 45951
rect 1584 45908 1636 45917
rect 4988 46044 5040 46096
rect 3792 46019 3844 46028
rect 3792 45985 3801 46019
rect 3801 45985 3835 46019
rect 3835 45985 3844 46019
rect 3792 45976 3844 45985
rect 4068 45976 4120 46028
rect 26976 46044 27028 46096
rect 9588 46019 9640 46028
rect 9588 45985 9597 46019
rect 9597 45985 9631 46019
rect 9631 45985 9640 46019
rect 9588 45976 9640 45985
rect 10140 46019 10192 46028
rect 10140 45985 10149 46019
rect 10149 45985 10183 46019
rect 10183 45985 10192 46019
rect 10140 45976 10192 45985
rect 4528 45840 4580 45892
rect 9864 45840 9916 45892
rect 20168 45976 20220 46028
rect 21272 46019 21324 46028
rect 21272 45985 21281 46019
rect 21281 45985 21315 46019
rect 21315 45985 21324 46019
rect 21272 45976 21324 45985
rect 22008 46019 22060 46028
rect 22008 45985 22017 46019
rect 22017 45985 22051 46019
rect 22051 45985 22060 46019
rect 22008 45976 22060 45985
rect 22560 46019 22612 46028
rect 22560 45985 22569 46019
rect 22569 45985 22603 46019
rect 22603 45985 22612 46019
rect 22560 45976 22612 45985
rect 26148 45976 26200 46028
rect 28172 46019 28224 46028
rect 28172 45985 28181 46019
rect 28181 45985 28215 46019
rect 28215 45985 28224 46019
rect 28172 45976 28224 45985
rect 14280 45951 14332 45960
rect 14280 45917 14289 45951
rect 14289 45917 14323 45951
rect 14323 45917 14332 45951
rect 14280 45908 14332 45917
rect 18236 45951 18288 45960
rect 14464 45883 14516 45892
rect 14464 45849 14473 45883
rect 14473 45849 14507 45883
rect 14507 45849 14516 45883
rect 14464 45840 14516 45849
rect 14740 45840 14792 45892
rect 18236 45917 18245 45951
rect 18245 45917 18279 45951
rect 18279 45917 18288 45951
rect 18236 45908 18288 45917
rect 25780 45908 25832 45960
rect 19892 45883 19944 45892
rect 18052 45772 18104 45824
rect 18328 45815 18380 45824
rect 18328 45781 18337 45815
rect 18337 45781 18371 45815
rect 18371 45781 18380 45815
rect 18328 45772 18380 45781
rect 19892 45849 19901 45883
rect 19901 45849 19935 45883
rect 19935 45849 19944 45883
rect 19892 45840 19944 45849
rect 22192 45883 22244 45892
rect 22192 45849 22201 45883
rect 22201 45849 22235 45883
rect 22235 45849 22244 45883
rect 22192 45840 22244 45849
rect 27528 45840 27580 45892
rect 26240 45772 26292 45824
rect 26884 45772 26936 45824
rect 27436 45772 27488 45824
rect 10214 45670 10266 45722
rect 10278 45670 10330 45722
rect 10342 45670 10394 45722
rect 10406 45670 10458 45722
rect 10470 45670 10522 45722
rect 19478 45670 19530 45722
rect 19542 45670 19594 45722
rect 19606 45670 19658 45722
rect 19670 45670 19722 45722
rect 19734 45670 19786 45722
rect 9864 45611 9916 45620
rect 9864 45577 9873 45611
rect 9873 45577 9907 45611
rect 9907 45577 9916 45611
rect 9864 45568 9916 45577
rect 14464 45611 14516 45620
rect 14464 45577 14473 45611
rect 14473 45577 14507 45611
rect 14507 45577 14516 45611
rect 14464 45568 14516 45577
rect 18052 45568 18104 45620
rect 19892 45568 19944 45620
rect 22192 45568 22244 45620
rect 4528 45543 4580 45552
rect 4528 45509 4537 45543
rect 4537 45509 4571 45543
rect 4571 45509 4580 45543
rect 4528 45500 4580 45509
rect 11704 45500 11756 45552
rect 18328 45543 18380 45552
rect 18328 45509 18337 45543
rect 18337 45509 18371 45543
rect 18371 45509 18380 45543
rect 18328 45500 18380 45509
rect 19524 45500 19576 45552
rect 22744 45543 22796 45552
rect 22744 45509 22753 45543
rect 22753 45509 22787 45543
rect 22787 45509 22796 45543
rect 22744 45500 22796 45509
rect 23940 45500 23992 45552
rect 26240 45543 26292 45552
rect 26240 45509 26249 45543
rect 26249 45509 26283 45543
rect 26283 45509 26292 45543
rect 27528 45543 27580 45552
rect 26240 45500 26292 45509
rect 27528 45509 27537 45543
rect 27537 45509 27571 45543
rect 27571 45509 27580 45543
rect 27528 45500 27580 45509
rect 1584 45475 1636 45484
rect 1584 45441 1593 45475
rect 1593 45441 1627 45475
rect 1627 45441 1636 45475
rect 1584 45432 1636 45441
rect 5448 45432 5500 45484
rect 9956 45475 10008 45484
rect 9956 45441 9965 45475
rect 9965 45441 9999 45475
rect 9999 45441 10008 45475
rect 9956 45432 10008 45441
rect 14372 45475 14424 45484
rect 14372 45441 14381 45475
rect 14381 45441 14415 45475
rect 14415 45441 14424 45475
rect 14372 45432 14424 45441
rect 18144 45475 18196 45484
rect 18144 45441 18153 45475
rect 18153 45441 18187 45475
rect 18187 45441 18196 45475
rect 18144 45432 18196 45441
rect 20444 45475 20496 45484
rect 20444 45441 20453 45475
rect 20453 45441 20487 45475
rect 20487 45441 20496 45475
rect 20444 45432 20496 45441
rect 22008 45475 22060 45484
rect 22008 45441 22017 45475
rect 22017 45441 22051 45475
rect 22051 45441 22060 45475
rect 22008 45432 22060 45441
rect 23296 45475 23348 45484
rect 1952 45364 2004 45416
rect 20 45296 72 45348
rect 14280 45364 14332 45416
rect 18696 45407 18748 45416
rect 18696 45373 18705 45407
rect 18705 45373 18739 45407
rect 18739 45373 18748 45407
rect 18696 45364 18748 45373
rect 23296 45441 23305 45475
rect 23305 45441 23339 45475
rect 23339 45441 23348 45475
rect 23296 45432 23348 45441
rect 26424 45475 26476 45484
rect 26424 45441 26433 45475
rect 26433 45441 26467 45475
rect 26467 45441 26476 45475
rect 27436 45475 27488 45484
rect 26424 45432 26476 45441
rect 27436 45441 27445 45475
rect 27445 45441 27479 45475
rect 27479 45441 27488 45475
rect 27436 45432 27488 45441
rect 5448 45296 5500 45348
rect 25780 45364 25832 45416
rect 25964 45407 26016 45416
rect 25964 45373 25973 45407
rect 25973 45373 26007 45407
rect 26007 45373 26016 45407
rect 25964 45364 26016 45373
rect 5582 45126 5634 45178
rect 5646 45126 5698 45178
rect 5710 45126 5762 45178
rect 5774 45126 5826 45178
rect 5838 45126 5890 45178
rect 14846 45126 14898 45178
rect 14910 45126 14962 45178
rect 14974 45126 15026 45178
rect 15038 45126 15090 45178
rect 15102 45126 15154 45178
rect 24110 45126 24162 45178
rect 24174 45126 24226 45178
rect 24238 45126 24290 45178
rect 24302 45126 24354 45178
rect 24366 45126 24418 45178
rect 1952 45067 2004 45076
rect 1952 45033 1961 45067
rect 1961 45033 1995 45067
rect 1995 45033 2004 45067
rect 1952 45024 2004 45033
rect 19340 45024 19392 45076
rect 20168 45067 20220 45076
rect 20168 45033 20177 45067
rect 20177 45033 20211 45067
rect 20211 45033 20220 45067
rect 20168 45024 20220 45033
rect 21916 45024 21968 45076
rect 14372 44956 14424 45008
rect 27436 44956 27488 45008
rect 12532 44931 12584 44940
rect 12532 44897 12541 44931
rect 12541 44897 12575 44931
rect 12575 44897 12584 44931
rect 12532 44888 12584 44897
rect 27528 44931 27580 44940
rect 27528 44897 27537 44931
rect 27537 44897 27571 44931
rect 27571 44897 27580 44931
rect 27528 44888 27580 44897
rect 27896 44888 27948 44940
rect 1952 44820 2004 44872
rect 19340 44820 19392 44872
rect 19524 44820 19576 44872
rect 11612 44752 11664 44804
rect 27620 44752 27672 44804
rect 10214 44582 10266 44634
rect 10278 44582 10330 44634
rect 10342 44582 10394 44634
rect 10406 44582 10458 44634
rect 10470 44582 10522 44634
rect 19478 44582 19530 44634
rect 19542 44582 19594 44634
rect 19606 44582 19658 44634
rect 19670 44582 19722 44634
rect 19734 44582 19786 44634
rect 11612 44523 11664 44532
rect 11612 44489 11621 44523
rect 11621 44489 11655 44523
rect 11655 44489 11664 44523
rect 11612 44480 11664 44489
rect 27620 44523 27672 44532
rect 27620 44489 27629 44523
rect 27629 44489 27663 44523
rect 27663 44489 27672 44523
rect 27620 44480 27672 44489
rect 11704 44387 11756 44396
rect 11704 44353 11713 44387
rect 11713 44353 11747 44387
rect 11747 44353 11756 44387
rect 11704 44344 11756 44353
rect 27436 44344 27488 44396
rect 1400 44140 1452 44192
rect 1584 44140 1636 44192
rect 2780 44183 2832 44192
rect 2780 44149 2789 44183
rect 2789 44149 2823 44183
rect 2823 44149 2832 44183
rect 2780 44140 2832 44149
rect 26332 44140 26384 44192
rect 5582 44038 5634 44090
rect 5646 44038 5698 44090
rect 5710 44038 5762 44090
rect 5774 44038 5826 44090
rect 5838 44038 5890 44090
rect 14846 44038 14898 44090
rect 14910 44038 14962 44090
rect 14974 44038 15026 44090
rect 15038 44038 15090 44090
rect 15102 44038 15154 44090
rect 24110 44038 24162 44090
rect 24174 44038 24226 44090
rect 24238 44038 24290 44090
rect 24302 44038 24354 44090
rect 24366 44038 24418 44090
rect 1400 43843 1452 43852
rect 1400 43809 1409 43843
rect 1409 43809 1443 43843
rect 1443 43809 1452 43843
rect 1400 43800 1452 43809
rect 1584 43843 1636 43852
rect 1584 43809 1593 43843
rect 1593 43809 1627 43843
rect 1627 43809 1636 43843
rect 1584 43800 1636 43809
rect 2872 43843 2924 43852
rect 2872 43809 2881 43843
rect 2881 43809 2915 43843
rect 2915 43809 2924 43843
rect 2872 43800 2924 43809
rect 27988 43843 28040 43852
rect 27988 43809 27997 43843
rect 27997 43809 28031 43843
rect 28031 43809 28040 43843
rect 27988 43800 28040 43809
rect 27068 43664 27120 43716
rect 10214 43494 10266 43546
rect 10278 43494 10330 43546
rect 10342 43494 10394 43546
rect 10406 43494 10458 43546
rect 10470 43494 10522 43546
rect 19478 43494 19530 43546
rect 19542 43494 19594 43546
rect 19606 43494 19658 43546
rect 19670 43494 19722 43546
rect 19734 43494 19786 43546
rect 27068 43435 27120 43444
rect 27068 43401 27077 43435
rect 27077 43401 27111 43435
rect 27111 43401 27120 43435
rect 27068 43392 27120 43401
rect 2780 43324 2832 43376
rect 28264 43256 28316 43308
rect 2964 43188 3016 43240
rect 3056 43231 3108 43240
rect 3056 43197 3065 43231
rect 3065 43197 3099 43231
rect 3099 43197 3108 43231
rect 3056 43188 3108 43197
rect 26516 43052 26568 43104
rect 5582 42950 5634 43002
rect 5646 42950 5698 43002
rect 5710 42950 5762 43002
rect 5774 42950 5826 43002
rect 5838 42950 5890 43002
rect 14846 42950 14898 43002
rect 14910 42950 14962 43002
rect 14974 42950 15026 43002
rect 15038 42950 15090 43002
rect 15102 42950 15154 43002
rect 24110 42950 24162 43002
rect 24174 42950 24226 43002
rect 24238 42950 24290 43002
rect 24302 42950 24354 43002
rect 24366 42950 24418 43002
rect 2964 42755 3016 42764
rect 2964 42721 2973 42755
rect 2973 42721 3007 42755
rect 3007 42721 3016 42755
rect 2964 42712 3016 42721
rect 26332 42755 26384 42764
rect 26332 42721 26341 42755
rect 26341 42721 26375 42755
rect 26375 42721 26384 42755
rect 26332 42712 26384 42721
rect 26516 42755 26568 42764
rect 26516 42721 26525 42755
rect 26525 42721 26559 42755
rect 26559 42721 26568 42755
rect 26516 42712 26568 42721
rect 28816 42712 28868 42764
rect 1768 42687 1820 42696
rect 1768 42653 1777 42687
rect 1777 42653 1811 42687
rect 1811 42653 1820 42687
rect 1768 42644 1820 42653
rect 3148 42644 3200 42696
rect 27712 42508 27764 42560
rect 10214 42406 10266 42458
rect 10278 42406 10330 42458
rect 10342 42406 10394 42458
rect 10406 42406 10458 42458
rect 10470 42406 10522 42458
rect 19478 42406 19530 42458
rect 19542 42406 19594 42458
rect 19606 42406 19658 42458
rect 19670 42406 19722 42458
rect 19734 42406 19786 42458
rect 27712 42211 27764 42220
rect 27712 42177 27721 42211
rect 27721 42177 27755 42211
rect 27755 42177 27764 42211
rect 27712 42168 27764 42177
rect 2780 42143 2832 42152
rect 2780 42109 2789 42143
rect 2789 42109 2823 42143
rect 2823 42109 2832 42143
rect 2780 42100 2832 42109
rect 3884 42100 3936 42152
rect 4620 42143 4672 42152
rect 4620 42109 4629 42143
rect 4629 42109 4663 42143
rect 4663 42109 4672 42143
rect 4620 42100 4672 42109
rect 1584 42007 1636 42016
rect 1584 41973 1593 42007
rect 1593 41973 1627 42007
rect 1627 41973 1636 42007
rect 1584 41964 1636 41973
rect 26424 42007 26476 42016
rect 26424 41973 26433 42007
rect 26433 41973 26467 42007
rect 26467 41973 26476 42007
rect 26424 41964 26476 41973
rect 27068 42007 27120 42016
rect 27068 41973 27077 42007
rect 27077 41973 27111 42007
rect 27111 41973 27120 42007
rect 27068 41964 27120 41973
rect 27804 42007 27856 42016
rect 27804 41973 27813 42007
rect 27813 41973 27847 42007
rect 27847 41973 27856 42007
rect 27804 41964 27856 41973
rect 5582 41862 5634 41914
rect 5646 41862 5698 41914
rect 5710 41862 5762 41914
rect 5774 41862 5826 41914
rect 5838 41862 5890 41914
rect 14846 41862 14898 41914
rect 14910 41862 14962 41914
rect 14974 41862 15026 41914
rect 15038 41862 15090 41914
rect 15102 41862 15154 41914
rect 24110 41862 24162 41914
rect 24174 41862 24226 41914
rect 24238 41862 24290 41914
rect 24302 41862 24354 41914
rect 24366 41862 24418 41914
rect 3884 41803 3936 41812
rect 3884 41769 3893 41803
rect 3893 41769 3927 41803
rect 3927 41769 3936 41803
rect 3884 41760 3936 41769
rect 4620 41803 4672 41812
rect 4620 41769 4629 41803
rect 4629 41769 4663 41803
rect 4663 41769 4672 41803
rect 4620 41760 4672 41769
rect 1400 41667 1452 41676
rect 1400 41633 1409 41667
rect 1409 41633 1443 41667
rect 1443 41633 1452 41667
rect 1400 41624 1452 41633
rect 1768 41624 1820 41676
rect 27068 41624 27120 41676
rect 28172 41667 28224 41676
rect 28172 41633 28181 41667
rect 28181 41633 28215 41667
rect 28215 41633 28224 41667
rect 28172 41624 28224 41633
rect 9956 41556 10008 41608
rect 10600 41556 10652 41608
rect 3056 41531 3108 41540
rect 3056 41497 3065 41531
rect 3065 41497 3099 41531
rect 3099 41497 3108 41531
rect 3056 41488 3108 41497
rect 27804 41488 27856 41540
rect 10214 41318 10266 41370
rect 10278 41318 10330 41370
rect 10342 41318 10394 41370
rect 10406 41318 10458 41370
rect 10470 41318 10522 41370
rect 19478 41318 19530 41370
rect 19542 41318 19594 41370
rect 19606 41318 19658 41370
rect 19670 41318 19722 41370
rect 19734 41318 19786 41370
rect 1584 41123 1636 41132
rect 1584 41089 1593 41123
rect 1593 41089 1627 41123
rect 1627 41089 1636 41123
rect 1584 41080 1636 41089
rect 26424 41123 26476 41132
rect 26424 41089 26433 41123
rect 26433 41089 26467 41123
rect 26467 41089 26476 41123
rect 26424 41080 26476 41089
rect 27344 41080 27396 41132
rect 2044 41012 2096 41064
rect 3240 41055 3292 41064
rect 3240 41021 3249 41055
rect 3249 41021 3283 41055
rect 3283 41021 3292 41055
rect 3240 41012 3292 41021
rect 25964 41055 26016 41064
rect 25964 41021 25973 41055
rect 25973 41021 26007 41055
rect 26007 41021 26016 41055
rect 25964 41012 26016 41021
rect 28172 40876 28224 40928
rect 5582 40774 5634 40826
rect 5646 40774 5698 40826
rect 5710 40774 5762 40826
rect 5774 40774 5826 40826
rect 5838 40774 5890 40826
rect 14846 40774 14898 40826
rect 14910 40774 14962 40826
rect 14974 40774 15026 40826
rect 15038 40774 15090 40826
rect 15102 40774 15154 40826
rect 24110 40774 24162 40826
rect 24174 40774 24226 40826
rect 24238 40774 24290 40826
rect 24302 40774 24354 40826
rect 24366 40774 24418 40826
rect 2044 40715 2096 40724
rect 2044 40681 2053 40715
rect 2053 40681 2087 40715
rect 2087 40681 2096 40715
rect 2044 40672 2096 40681
rect 3056 40672 3108 40724
rect 27528 40579 27580 40588
rect 27528 40545 27537 40579
rect 27537 40545 27571 40579
rect 27571 40545 27580 40579
rect 27528 40536 27580 40545
rect 28172 40579 28224 40588
rect 28172 40545 28181 40579
rect 28181 40545 28215 40579
rect 28215 40545 28224 40579
rect 28172 40536 28224 40545
rect 27988 40443 28040 40452
rect 27988 40409 27997 40443
rect 27997 40409 28031 40443
rect 28031 40409 28040 40443
rect 27988 40400 28040 40409
rect 27620 40332 27672 40384
rect 10214 40230 10266 40282
rect 10278 40230 10330 40282
rect 10342 40230 10394 40282
rect 10406 40230 10458 40282
rect 10470 40230 10522 40282
rect 19478 40230 19530 40282
rect 19542 40230 19594 40282
rect 19606 40230 19658 40282
rect 19670 40230 19722 40282
rect 19734 40230 19786 40282
rect 27988 40128 28040 40180
rect 19340 40060 19392 40112
rect 27344 40060 27396 40112
rect 27712 40035 27764 40044
rect 27712 40001 27721 40035
rect 27721 40001 27755 40035
rect 27755 40001 27764 40035
rect 27712 39992 27764 40001
rect 26332 39788 26384 39840
rect 5582 39686 5634 39738
rect 5646 39686 5698 39738
rect 5710 39686 5762 39738
rect 5774 39686 5826 39738
rect 5838 39686 5890 39738
rect 14846 39686 14898 39738
rect 14910 39686 14962 39738
rect 14974 39686 15026 39738
rect 15038 39686 15090 39738
rect 15102 39686 15154 39738
rect 24110 39686 24162 39738
rect 24174 39686 24226 39738
rect 24238 39686 24290 39738
rect 24302 39686 24354 39738
rect 24366 39686 24418 39738
rect 21824 39516 21876 39568
rect 26332 39491 26384 39500
rect 26332 39457 26341 39491
rect 26341 39457 26375 39491
rect 26375 39457 26384 39491
rect 26332 39448 26384 39457
rect 28172 39491 28224 39500
rect 28172 39457 28181 39491
rect 28181 39457 28215 39491
rect 28215 39457 28224 39491
rect 28172 39448 28224 39457
rect 20812 39380 20864 39432
rect 21180 39423 21232 39432
rect 21180 39389 21189 39423
rect 21189 39389 21223 39423
rect 21223 39389 21232 39423
rect 21180 39380 21232 39389
rect 21272 39380 21324 39432
rect 26516 39355 26568 39364
rect 20536 39244 20588 39296
rect 20904 39244 20956 39296
rect 26516 39321 26525 39355
rect 26525 39321 26559 39355
rect 26559 39321 26568 39355
rect 26516 39312 26568 39321
rect 10214 39142 10266 39194
rect 10278 39142 10330 39194
rect 10342 39142 10394 39194
rect 10406 39142 10458 39194
rect 10470 39142 10522 39194
rect 19478 39142 19530 39194
rect 19542 39142 19594 39194
rect 19606 39142 19658 39194
rect 19670 39142 19722 39194
rect 19734 39142 19786 39194
rect 26516 39040 26568 39092
rect 20812 38972 20864 39024
rect 19340 38904 19392 38956
rect 19892 38904 19944 38956
rect 21824 38947 21876 38956
rect 21824 38913 21833 38947
rect 21833 38913 21867 38947
rect 21867 38913 21876 38947
rect 21824 38904 21876 38913
rect 22376 38904 22428 38956
rect 27804 38904 27856 38956
rect 28264 38904 28316 38956
rect 21272 38836 21324 38888
rect 22100 38879 22152 38888
rect 22100 38845 22109 38879
rect 22109 38845 22143 38879
rect 22143 38845 22152 38879
rect 22100 38836 22152 38845
rect 20996 38768 21048 38820
rect 1676 38743 1728 38752
rect 1676 38709 1685 38743
rect 1685 38709 1719 38743
rect 1719 38709 1728 38743
rect 1676 38700 1728 38709
rect 19524 38700 19576 38752
rect 20812 38743 20864 38752
rect 20812 38709 20821 38743
rect 20821 38709 20855 38743
rect 20855 38709 20864 38743
rect 20812 38700 20864 38709
rect 21364 38700 21416 38752
rect 22284 38743 22336 38752
rect 22284 38709 22293 38743
rect 22293 38709 22327 38743
rect 22327 38709 22336 38743
rect 22284 38700 22336 38709
rect 26332 38700 26384 38752
rect 5582 38598 5634 38650
rect 5646 38598 5698 38650
rect 5710 38598 5762 38650
rect 5774 38598 5826 38650
rect 5838 38598 5890 38650
rect 14846 38598 14898 38650
rect 14910 38598 14962 38650
rect 14974 38598 15026 38650
rect 15038 38598 15090 38650
rect 15102 38598 15154 38650
rect 24110 38598 24162 38650
rect 24174 38598 24226 38650
rect 24238 38598 24290 38650
rect 24302 38598 24354 38650
rect 24366 38598 24418 38650
rect 1676 38360 1728 38412
rect 2780 38403 2832 38412
rect 2780 38369 2789 38403
rect 2789 38369 2823 38403
rect 2823 38369 2832 38403
rect 2780 38360 2832 38369
rect 20812 38360 20864 38412
rect 26332 38403 26384 38412
rect 26332 38369 26341 38403
rect 26341 38369 26375 38403
rect 26375 38369 26384 38403
rect 26332 38360 26384 38369
rect 28724 38360 28776 38412
rect 18788 38292 18840 38344
rect 19524 38335 19576 38344
rect 19524 38301 19558 38335
rect 19558 38301 19576 38335
rect 19524 38292 19576 38301
rect 20536 38292 20588 38344
rect 23756 38335 23808 38344
rect 23756 38301 23765 38335
rect 23765 38301 23799 38335
rect 23799 38301 23808 38335
rect 23756 38292 23808 38301
rect 2136 38224 2188 38276
rect 22836 38224 22888 38276
rect 27712 38224 27764 38276
rect 22560 38156 22612 38208
rect 10214 38054 10266 38106
rect 10278 38054 10330 38106
rect 10342 38054 10394 38106
rect 10406 38054 10458 38106
rect 10470 38054 10522 38106
rect 19478 38054 19530 38106
rect 19542 38054 19594 38106
rect 19606 38054 19658 38106
rect 19670 38054 19722 38106
rect 19734 38054 19786 38106
rect 2136 37995 2188 38004
rect 2136 37961 2145 37995
rect 2145 37961 2179 37995
rect 2179 37961 2188 37995
rect 2136 37952 2188 37961
rect 19340 37952 19392 38004
rect 21180 37952 21232 38004
rect 22836 37995 22888 38004
rect 22836 37961 22845 37995
rect 22845 37961 22879 37995
rect 22879 37961 22888 37995
rect 22836 37952 22888 37961
rect 27712 37995 27764 38004
rect 27712 37961 27721 37995
rect 27721 37961 27755 37995
rect 27755 37961 27764 37995
rect 27712 37952 27764 37961
rect 2228 37859 2280 37868
rect 2228 37825 2237 37859
rect 2237 37825 2271 37859
rect 2271 37825 2280 37859
rect 2228 37816 2280 37825
rect 20168 37859 20220 37868
rect 20168 37825 20177 37859
rect 20177 37825 20211 37859
rect 20211 37825 20220 37859
rect 20168 37816 20220 37825
rect 20536 37884 20588 37936
rect 21272 37927 21324 37936
rect 21272 37893 21281 37927
rect 21281 37893 21315 37927
rect 21315 37893 21324 37927
rect 21272 37884 21324 37893
rect 20076 37791 20128 37800
rect 20076 37757 20085 37791
rect 20085 37757 20119 37791
rect 20119 37757 20128 37791
rect 20076 37748 20128 37757
rect 20352 37791 20404 37800
rect 20352 37757 20361 37791
rect 20361 37757 20395 37791
rect 20395 37757 20404 37791
rect 20352 37748 20404 37757
rect 20536 37680 20588 37732
rect 3240 37612 3292 37664
rect 20812 37612 20864 37664
rect 22284 37816 22336 37868
rect 22376 37680 22428 37732
rect 22560 37859 22612 37868
rect 22560 37825 22569 37859
rect 22569 37825 22603 37859
rect 22603 37825 22612 37859
rect 22560 37816 22612 37825
rect 27712 37816 27764 37868
rect 22744 37612 22796 37664
rect 5582 37510 5634 37562
rect 5646 37510 5698 37562
rect 5710 37510 5762 37562
rect 5774 37510 5826 37562
rect 5838 37510 5890 37562
rect 14846 37510 14898 37562
rect 14910 37510 14962 37562
rect 14974 37510 15026 37562
rect 15038 37510 15090 37562
rect 15102 37510 15154 37562
rect 24110 37510 24162 37562
rect 24174 37510 24226 37562
rect 24238 37510 24290 37562
rect 24302 37510 24354 37562
rect 24366 37510 24418 37562
rect 19892 37451 19944 37460
rect 19892 37417 19901 37451
rect 19901 37417 19935 37451
rect 19935 37417 19944 37451
rect 19892 37408 19944 37417
rect 22100 37408 22152 37460
rect 27896 37272 27948 37324
rect 28172 37272 28224 37324
rect 1400 37247 1452 37256
rect 1400 37213 1409 37247
rect 1409 37213 1443 37247
rect 1443 37213 1452 37247
rect 1400 37204 1452 37213
rect 3240 37247 3292 37256
rect 3240 37213 3249 37247
rect 3249 37213 3283 37247
rect 3283 37213 3292 37247
rect 20168 37247 20220 37256
rect 3240 37204 3292 37213
rect 20168 37213 20177 37247
rect 20177 37213 20211 37247
rect 20211 37213 20220 37247
rect 20168 37204 20220 37213
rect 20904 37247 20956 37256
rect 20904 37213 20913 37247
rect 20913 37213 20947 37247
rect 20947 37213 20956 37247
rect 20904 37204 20956 37213
rect 22560 37204 22612 37256
rect 26792 37247 26844 37256
rect 26792 37213 26801 37247
rect 26801 37213 26835 37247
rect 26835 37213 26844 37247
rect 26792 37204 26844 37213
rect 2780 37136 2832 37188
rect 20536 37136 20588 37188
rect 20260 37068 20312 37120
rect 22376 37136 22428 37188
rect 20996 37111 21048 37120
rect 20996 37077 21005 37111
rect 21005 37077 21039 37111
rect 21039 37077 21048 37111
rect 20996 37068 21048 37077
rect 21456 37068 21508 37120
rect 26608 37111 26660 37120
rect 26608 37077 26617 37111
rect 26617 37077 26651 37111
rect 26651 37077 26660 37111
rect 26608 37068 26660 37077
rect 10214 36966 10266 37018
rect 10278 36966 10330 37018
rect 10342 36966 10394 37018
rect 10406 36966 10458 37018
rect 10470 36966 10522 37018
rect 19478 36966 19530 37018
rect 19542 36966 19594 37018
rect 19606 36966 19658 37018
rect 19670 36966 19722 37018
rect 19734 36966 19786 37018
rect 2780 36907 2832 36916
rect 2780 36873 2789 36907
rect 2789 36873 2823 36907
rect 2823 36873 2832 36907
rect 2780 36864 2832 36873
rect 1860 36771 1912 36780
rect 1860 36737 1869 36771
rect 1869 36737 1903 36771
rect 1903 36737 1912 36771
rect 1860 36728 1912 36737
rect 2044 36728 2096 36780
rect 17960 36771 18012 36780
rect 17960 36737 17969 36771
rect 17969 36737 18003 36771
rect 18003 36737 18012 36771
rect 17960 36728 18012 36737
rect 22652 36771 22704 36780
rect 22652 36737 22661 36771
rect 22661 36737 22695 36771
rect 22695 36737 22704 36771
rect 22652 36728 22704 36737
rect 27620 36728 27672 36780
rect 18420 36660 18472 36712
rect 23296 36660 23348 36712
rect 2320 36524 2372 36576
rect 16948 36524 17000 36576
rect 22468 36524 22520 36576
rect 27988 36524 28040 36576
rect 5582 36422 5634 36474
rect 5646 36422 5698 36474
rect 5710 36422 5762 36474
rect 5774 36422 5826 36474
rect 5838 36422 5890 36474
rect 14846 36422 14898 36474
rect 14910 36422 14962 36474
rect 14974 36422 15026 36474
rect 15038 36422 15090 36474
rect 15102 36422 15154 36474
rect 24110 36422 24162 36474
rect 24174 36422 24226 36474
rect 24238 36422 24290 36474
rect 24302 36422 24354 36474
rect 24366 36422 24418 36474
rect 20076 36363 20128 36372
rect 20076 36329 20085 36363
rect 20085 36329 20119 36363
rect 20119 36329 20128 36363
rect 20076 36320 20128 36329
rect 22468 36252 22520 36304
rect 17960 36116 18012 36168
rect 20720 36116 20772 36168
rect 18328 36048 18380 36100
rect 19340 36048 19392 36100
rect 19892 36048 19944 36100
rect 20904 36116 20956 36168
rect 22376 36184 22428 36236
rect 22192 36159 22244 36168
rect 22192 36125 22201 36159
rect 22201 36125 22235 36159
rect 22235 36125 22244 36159
rect 22192 36116 22244 36125
rect 22744 36116 22796 36168
rect 27896 36252 27948 36304
rect 27528 36227 27580 36236
rect 27528 36193 27537 36227
rect 27537 36193 27571 36227
rect 27571 36193 27580 36227
rect 27528 36184 27580 36193
rect 27988 36227 28040 36236
rect 27988 36193 27997 36227
rect 27997 36193 28031 36227
rect 28031 36193 28040 36227
rect 27988 36184 28040 36193
rect 25228 36159 25280 36168
rect 20996 36091 21048 36100
rect 20996 36057 21005 36091
rect 21005 36057 21039 36091
rect 21039 36057 21048 36091
rect 20996 36048 21048 36057
rect 21272 35980 21324 36032
rect 22376 35980 22428 36032
rect 25228 36125 25237 36159
rect 25237 36125 25271 36159
rect 25271 36125 25280 36159
rect 25228 36116 25280 36125
rect 26792 36116 26844 36168
rect 25596 36048 25648 36100
rect 24400 35980 24452 36032
rect 10214 35878 10266 35930
rect 10278 35878 10330 35930
rect 10342 35878 10394 35930
rect 10406 35878 10458 35930
rect 10470 35878 10522 35930
rect 19478 35878 19530 35930
rect 19542 35878 19594 35930
rect 19606 35878 19658 35930
rect 19670 35878 19722 35930
rect 19734 35878 19786 35930
rect 16948 35751 17000 35760
rect 16948 35717 16957 35751
rect 16957 35717 16991 35751
rect 16991 35717 17000 35751
rect 16948 35708 17000 35717
rect 18236 35751 18288 35760
rect 18236 35717 18245 35751
rect 18245 35717 18279 35751
rect 18279 35717 18288 35751
rect 18236 35708 18288 35717
rect 18696 35708 18748 35760
rect 17960 35640 18012 35692
rect 18788 35683 18840 35692
rect 18788 35649 18797 35683
rect 18797 35649 18831 35683
rect 18831 35649 18840 35683
rect 18788 35640 18840 35649
rect 19340 35640 19392 35692
rect 20996 35776 21048 35828
rect 20720 35708 20772 35760
rect 25228 35776 25280 35828
rect 21548 35708 21600 35760
rect 21088 35683 21140 35692
rect 21088 35649 21099 35683
rect 21099 35649 21140 35683
rect 21088 35640 21140 35649
rect 22468 35683 22520 35692
rect 22468 35649 22477 35683
rect 22477 35649 22511 35683
rect 22511 35649 22520 35683
rect 22468 35640 22520 35649
rect 24400 35751 24452 35760
rect 24400 35717 24418 35751
rect 24418 35717 24452 35751
rect 24400 35708 24452 35717
rect 25596 35683 25648 35692
rect 22284 35572 22336 35624
rect 25596 35649 25605 35683
rect 25605 35649 25639 35683
rect 25639 35649 25648 35683
rect 25596 35640 25648 35649
rect 27252 35640 27304 35692
rect 22652 35504 22704 35556
rect 25872 35572 25924 35624
rect 27712 35572 27764 35624
rect 1400 35436 1452 35488
rect 3608 35436 3660 35488
rect 11704 35436 11756 35488
rect 21548 35436 21600 35488
rect 23112 35436 23164 35488
rect 23296 35479 23348 35488
rect 23296 35445 23305 35479
rect 23305 35445 23339 35479
rect 23339 35445 23348 35479
rect 23296 35436 23348 35445
rect 23480 35436 23532 35488
rect 23756 35436 23808 35488
rect 24676 35436 24728 35488
rect 26332 35436 26384 35488
rect 5582 35334 5634 35386
rect 5646 35334 5698 35386
rect 5710 35334 5762 35386
rect 5774 35334 5826 35386
rect 5838 35334 5890 35386
rect 14846 35334 14898 35386
rect 14910 35334 14962 35386
rect 14974 35334 15026 35386
rect 15038 35334 15090 35386
rect 15102 35334 15154 35386
rect 24110 35334 24162 35386
rect 24174 35334 24226 35386
rect 24238 35334 24290 35386
rect 24302 35334 24354 35386
rect 24366 35334 24418 35386
rect 20720 35232 20772 35284
rect 21180 35232 21232 35284
rect 22192 35232 22244 35284
rect 27252 35275 27304 35284
rect 27252 35241 27261 35275
rect 27261 35241 27295 35275
rect 27295 35241 27304 35275
rect 27252 35232 27304 35241
rect 1400 35139 1452 35148
rect 1400 35105 1409 35139
rect 1409 35105 1443 35139
rect 1443 35105 1452 35139
rect 1400 35096 1452 35105
rect 2780 35139 2832 35148
rect 2780 35105 2789 35139
rect 2789 35105 2823 35139
rect 2823 35105 2832 35139
rect 2780 35096 2832 35105
rect 18328 35139 18380 35148
rect 18328 35105 18337 35139
rect 18337 35105 18371 35139
rect 18371 35105 18380 35139
rect 18328 35096 18380 35105
rect 17960 35028 18012 35080
rect 20996 35096 21048 35148
rect 23572 35164 23624 35216
rect 22560 35096 22612 35148
rect 23664 35096 23716 35148
rect 24676 35096 24728 35148
rect 23112 35071 23164 35080
rect 1492 34892 1544 34944
rect 19892 34892 19944 34944
rect 21088 34935 21140 34944
rect 21088 34901 21097 34935
rect 21097 34901 21131 34935
rect 21131 34901 21140 34935
rect 21088 34892 21140 34901
rect 21272 35003 21324 35012
rect 21272 34969 21281 35003
rect 21281 34969 21315 35003
rect 21315 34969 21324 35003
rect 21272 34960 21324 34969
rect 22100 34892 22152 34944
rect 23112 35037 23121 35071
rect 23121 35037 23155 35071
rect 23155 35037 23164 35071
rect 23112 35028 23164 35037
rect 26608 35028 26660 35080
rect 27712 35071 27764 35080
rect 27712 35037 27721 35071
rect 27721 35037 27755 35071
rect 27755 35037 27764 35071
rect 27712 35028 27764 35037
rect 24860 34892 24912 34944
rect 25596 34960 25648 35012
rect 27804 34960 27856 35012
rect 28816 34960 28868 35012
rect 27436 34892 27488 34944
rect 10214 34790 10266 34842
rect 10278 34790 10330 34842
rect 10342 34790 10394 34842
rect 10406 34790 10458 34842
rect 10470 34790 10522 34842
rect 19478 34790 19530 34842
rect 19542 34790 19594 34842
rect 19606 34790 19658 34842
rect 19670 34790 19722 34842
rect 19734 34790 19786 34842
rect 2228 34688 2280 34740
rect 1768 34663 1820 34672
rect 1768 34629 1777 34663
rect 1777 34629 1811 34663
rect 1811 34629 1820 34663
rect 1768 34620 1820 34629
rect 1952 34620 2004 34672
rect 20444 34620 20496 34672
rect 20996 34663 21048 34672
rect 20996 34629 21005 34663
rect 21005 34629 21039 34663
rect 21039 34629 21048 34663
rect 20996 34620 21048 34629
rect 21088 34663 21140 34672
rect 21088 34629 21123 34663
rect 21123 34629 21140 34663
rect 21088 34620 21140 34629
rect 21272 34620 21324 34672
rect 3608 34595 3660 34604
rect 3608 34561 3617 34595
rect 3617 34561 3651 34595
rect 3651 34561 3660 34595
rect 3608 34552 3660 34561
rect 17960 34552 18012 34604
rect 19892 34552 19944 34604
rect 3424 34527 3476 34536
rect 3424 34493 3433 34527
rect 3433 34493 3467 34527
rect 3467 34493 3476 34527
rect 3424 34484 3476 34493
rect 20628 34527 20680 34536
rect 20628 34493 20637 34527
rect 20637 34493 20671 34527
rect 20671 34493 20680 34527
rect 20628 34484 20680 34493
rect 20904 34595 20956 34604
rect 20904 34561 20913 34595
rect 20913 34561 20947 34595
rect 20947 34561 20956 34595
rect 24676 34620 24728 34672
rect 27436 34663 27488 34672
rect 20904 34552 20956 34561
rect 22192 34595 22244 34604
rect 22192 34561 22201 34595
rect 22201 34561 22235 34595
rect 22235 34561 22244 34595
rect 22192 34552 22244 34561
rect 26332 34552 26384 34604
rect 27436 34629 27445 34663
rect 27445 34629 27479 34663
rect 27479 34629 27488 34663
rect 27436 34620 27488 34629
rect 27712 34552 27764 34604
rect 23296 34348 23348 34400
rect 25044 34391 25096 34400
rect 25044 34357 25053 34391
rect 25053 34357 25087 34391
rect 25087 34357 25096 34391
rect 25044 34348 25096 34357
rect 5582 34246 5634 34298
rect 5646 34246 5698 34298
rect 5710 34246 5762 34298
rect 5774 34246 5826 34298
rect 5838 34246 5890 34298
rect 14846 34246 14898 34298
rect 14910 34246 14962 34298
rect 14974 34246 15026 34298
rect 15038 34246 15090 34298
rect 15102 34246 15154 34298
rect 24110 34246 24162 34298
rect 24174 34246 24226 34298
rect 24238 34246 24290 34298
rect 24302 34246 24354 34298
rect 24366 34246 24418 34298
rect 3424 34144 3476 34196
rect 20168 34187 20220 34196
rect 20168 34153 20177 34187
rect 20177 34153 20211 34187
rect 20211 34153 20220 34187
rect 20168 34144 20220 34153
rect 2688 33983 2740 33992
rect 2688 33949 2697 33983
rect 2697 33949 2731 33983
rect 2731 33949 2740 33983
rect 2688 33940 2740 33949
rect 20444 34076 20496 34128
rect 19892 33872 19944 33924
rect 20168 33804 20220 33856
rect 20536 33915 20588 33924
rect 20536 33881 20545 33915
rect 20545 33881 20579 33915
rect 20579 33881 20588 33915
rect 20536 33872 20588 33881
rect 20904 34144 20956 34196
rect 23572 34144 23624 34196
rect 23296 34076 23348 34128
rect 21088 34008 21140 34060
rect 21272 34051 21324 34060
rect 21272 34017 21281 34051
rect 21281 34017 21315 34051
rect 21315 34017 21324 34051
rect 21272 34008 21324 34017
rect 22192 34008 22244 34060
rect 22652 34008 22704 34060
rect 27528 34051 27580 34060
rect 27528 34017 27537 34051
rect 27537 34017 27571 34051
rect 27571 34017 27580 34051
rect 27528 34008 27580 34017
rect 28172 34051 28224 34060
rect 28172 34017 28181 34051
rect 28181 34017 28215 34051
rect 28215 34017 28224 34051
rect 28172 34008 28224 34017
rect 20720 33983 20772 33992
rect 20720 33949 20729 33983
rect 20729 33949 20763 33983
rect 20763 33949 20772 33983
rect 20720 33940 20772 33949
rect 21824 33940 21876 33992
rect 22468 33940 22520 33992
rect 23388 33940 23440 33992
rect 25044 33940 25096 33992
rect 23848 33915 23900 33924
rect 23848 33881 23857 33915
rect 23857 33881 23891 33915
rect 23891 33881 23900 33915
rect 23848 33872 23900 33881
rect 24584 33915 24636 33924
rect 20904 33804 20956 33856
rect 24584 33881 24593 33915
rect 24593 33881 24627 33915
rect 24627 33881 24636 33915
rect 24584 33872 24636 33881
rect 27160 33872 27212 33924
rect 25136 33847 25188 33856
rect 25136 33813 25145 33847
rect 25145 33813 25179 33847
rect 25179 33813 25188 33847
rect 25136 33804 25188 33813
rect 10214 33702 10266 33754
rect 10278 33702 10330 33754
rect 10342 33702 10394 33754
rect 10406 33702 10458 33754
rect 10470 33702 10522 33754
rect 19478 33702 19530 33754
rect 19542 33702 19594 33754
rect 19606 33702 19658 33754
rect 19670 33702 19722 33754
rect 19734 33702 19786 33754
rect 24584 33643 24636 33652
rect 18328 33532 18380 33584
rect 18788 33532 18840 33584
rect 24584 33609 24593 33643
rect 24593 33609 24627 33643
rect 24627 33609 24636 33643
rect 24584 33600 24636 33609
rect 27160 33643 27212 33652
rect 27160 33609 27169 33643
rect 27169 33609 27203 33643
rect 27203 33609 27212 33643
rect 27160 33600 27212 33609
rect 22652 33575 22704 33584
rect 19892 33464 19944 33516
rect 22652 33541 22661 33575
rect 22661 33541 22695 33575
rect 22695 33541 22704 33575
rect 22652 33532 22704 33541
rect 23572 33532 23624 33584
rect 27620 33532 27672 33584
rect 27896 33532 27948 33584
rect 20168 33507 20220 33516
rect 20168 33473 20177 33507
rect 20177 33473 20211 33507
rect 20211 33473 20220 33507
rect 20168 33464 20220 33473
rect 25136 33464 25188 33516
rect 26976 33464 27028 33516
rect 27712 33507 27764 33516
rect 27712 33473 27721 33507
rect 27721 33473 27755 33507
rect 27755 33473 27764 33507
rect 27712 33464 27764 33473
rect 20536 33328 20588 33380
rect 19984 33260 20036 33312
rect 22744 33260 22796 33312
rect 23480 33260 23532 33312
rect 26240 33260 26292 33312
rect 26332 33260 26384 33312
rect 5582 33158 5634 33210
rect 5646 33158 5698 33210
rect 5710 33158 5762 33210
rect 5774 33158 5826 33210
rect 5838 33158 5890 33210
rect 14846 33158 14898 33210
rect 14910 33158 14962 33210
rect 14974 33158 15026 33210
rect 15038 33158 15090 33210
rect 15102 33158 15154 33210
rect 24110 33158 24162 33210
rect 24174 33158 24226 33210
rect 24238 33158 24290 33210
rect 24302 33158 24354 33210
rect 24366 33158 24418 33210
rect 19340 33056 19392 33108
rect 23572 33056 23624 33108
rect 19984 33031 20036 33040
rect 19984 32997 19993 33031
rect 19993 32997 20027 33031
rect 20027 32997 20036 33031
rect 19984 32988 20036 32997
rect 20628 32988 20680 33040
rect 22376 32988 22428 33040
rect 20168 32895 20220 32904
rect 20168 32861 20177 32895
rect 20177 32861 20211 32895
rect 20211 32861 20220 32895
rect 20168 32852 20220 32861
rect 21732 32852 21784 32904
rect 22376 32895 22428 32904
rect 22376 32861 22385 32895
rect 22385 32861 22419 32895
rect 22419 32861 22428 32895
rect 22376 32852 22428 32861
rect 22560 32895 22612 32904
rect 22560 32861 22569 32895
rect 22569 32861 22603 32895
rect 22603 32861 22612 32895
rect 22560 32852 22612 32861
rect 23664 32988 23716 33040
rect 22744 32895 22796 32904
rect 22744 32861 22753 32895
rect 22753 32861 22787 32895
rect 22787 32861 22796 32895
rect 26976 32988 27028 33040
rect 26332 32963 26384 32972
rect 26332 32929 26341 32963
rect 26341 32929 26375 32963
rect 26375 32929 26384 32963
rect 26332 32920 26384 32929
rect 28080 32963 28132 32972
rect 28080 32929 28089 32963
rect 28089 32929 28123 32963
rect 28123 32929 28132 32963
rect 28080 32920 28132 32929
rect 22744 32852 22796 32861
rect 20720 32784 20772 32836
rect 23388 32784 23440 32836
rect 23664 32759 23716 32768
rect 23664 32725 23673 32759
rect 23673 32725 23707 32759
rect 23707 32725 23716 32759
rect 23664 32716 23716 32725
rect 10214 32614 10266 32666
rect 10278 32614 10330 32666
rect 10342 32614 10394 32666
rect 10406 32614 10458 32666
rect 10470 32614 10522 32666
rect 19478 32614 19530 32666
rect 19542 32614 19594 32666
rect 19606 32614 19658 32666
rect 19670 32614 19722 32666
rect 19734 32614 19786 32666
rect 20168 32512 20220 32564
rect 18328 32444 18380 32496
rect 20260 32444 20312 32496
rect 16764 32376 16816 32428
rect 20076 32376 20128 32428
rect 21088 32376 21140 32428
rect 21180 32419 21232 32428
rect 21180 32385 21189 32419
rect 21189 32385 21223 32419
rect 21223 32385 21232 32419
rect 21180 32376 21232 32385
rect 21548 32376 21600 32428
rect 23664 32376 23716 32428
rect 26976 32419 27028 32428
rect 26976 32385 26985 32419
rect 26985 32385 27019 32419
rect 27019 32385 27028 32419
rect 26976 32376 27028 32385
rect 28448 32376 28500 32428
rect 20720 32308 20772 32360
rect 21272 32308 21324 32360
rect 22468 32308 22520 32360
rect 22744 32308 22796 32360
rect 25964 32351 26016 32360
rect 25964 32317 25973 32351
rect 25973 32317 26007 32351
rect 26007 32317 26016 32351
rect 25964 32308 26016 32317
rect 26240 32308 26292 32360
rect 1400 32172 1452 32224
rect 17684 32172 17736 32224
rect 19616 32172 19668 32224
rect 21732 32172 21784 32224
rect 22284 32215 22336 32224
rect 22284 32181 22293 32215
rect 22293 32181 22327 32215
rect 22327 32181 22336 32215
rect 22284 32172 22336 32181
rect 27252 32172 27304 32224
rect 5582 32070 5634 32122
rect 5646 32070 5698 32122
rect 5710 32070 5762 32122
rect 5774 32070 5826 32122
rect 5838 32070 5890 32122
rect 14846 32070 14898 32122
rect 14910 32070 14962 32122
rect 14974 32070 15026 32122
rect 15038 32070 15090 32122
rect 15102 32070 15154 32122
rect 24110 32070 24162 32122
rect 24174 32070 24226 32122
rect 24238 32070 24290 32122
rect 24302 32070 24354 32122
rect 24366 32070 24418 32122
rect 3332 31968 3384 32020
rect 16764 31900 16816 31952
rect 20536 31900 20588 31952
rect 22560 31968 22612 32020
rect 23664 31968 23716 32020
rect 1400 31875 1452 31884
rect 1400 31841 1409 31875
rect 1409 31841 1443 31875
rect 1443 31841 1452 31875
rect 1400 31832 1452 31841
rect 1860 31875 1912 31884
rect 1860 31841 1869 31875
rect 1869 31841 1903 31875
rect 1903 31841 1912 31875
rect 1860 31832 1912 31841
rect 17592 31875 17644 31884
rect 17592 31841 17601 31875
rect 17601 31841 17635 31875
rect 17635 31841 17644 31875
rect 17592 31832 17644 31841
rect 17868 31832 17920 31884
rect 16856 31764 16908 31816
rect 20720 31832 20772 31884
rect 22652 31832 22704 31884
rect 23112 31832 23164 31884
rect 27252 31875 27304 31884
rect 27252 31841 27261 31875
rect 27261 31841 27295 31875
rect 27295 31841 27304 31875
rect 27252 31832 27304 31841
rect 19616 31807 19668 31816
rect 19616 31773 19625 31807
rect 19625 31773 19659 31807
rect 19659 31773 19668 31807
rect 19616 31764 19668 31773
rect 20076 31807 20128 31816
rect 20076 31773 20085 31807
rect 20085 31773 20119 31807
rect 20119 31773 20128 31807
rect 20076 31764 20128 31773
rect 20444 31764 20496 31816
rect 21180 31764 21232 31816
rect 22100 31807 22152 31816
rect 22100 31773 22109 31807
rect 22109 31773 22143 31807
rect 22143 31773 22152 31807
rect 22100 31764 22152 31773
rect 22468 31807 22520 31816
rect 22468 31773 22477 31807
rect 22477 31773 22511 31807
rect 22511 31773 22520 31807
rect 22468 31764 22520 31773
rect 23848 31764 23900 31816
rect 27436 31807 27488 31816
rect 27436 31773 27445 31807
rect 27445 31773 27479 31807
rect 27479 31773 27488 31807
rect 27436 31764 27488 31773
rect 28172 31764 28224 31816
rect 1584 31739 1636 31748
rect 1584 31705 1593 31739
rect 1593 31705 1627 31739
rect 1627 31705 1636 31739
rect 1584 31696 1636 31705
rect 22192 31696 22244 31748
rect 17132 31671 17184 31680
rect 17132 31637 17141 31671
rect 17141 31637 17175 31671
rect 17175 31637 17184 31671
rect 17132 31628 17184 31637
rect 17592 31628 17644 31680
rect 18512 31671 18564 31680
rect 18512 31637 18521 31671
rect 18521 31637 18555 31671
rect 18555 31637 18564 31671
rect 18512 31628 18564 31637
rect 10214 31526 10266 31578
rect 10278 31526 10330 31578
rect 10342 31526 10394 31578
rect 10406 31526 10458 31578
rect 10470 31526 10522 31578
rect 19478 31526 19530 31578
rect 19542 31526 19594 31578
rect 19606 31526 19658 31578
rect 19670 31526 19722 31578
rect 19734 31526 19786 31578
rect 1584 31424 1636 31476
rect 16856 31467 16908 31476
rect 16856 31433 16865 31467
rect 16865 31433 16899 31467
rect 16899 31433 16908 31467
rect 16856 31424 16908 31433
rect 23848 31424 23900 31476
rect 17132 31356 17184 31408
rect 18512 31399 18564 31408
rect 18512 31365 18546 31399
rect 18546 31365 18564 31399
rect 18512 31356 18564 31365
rect 2228 31288 2280 31340
rect 18328 31288 18380 31340
rect 20168 31288 20220 31340
rect 22100 31288 22152 31340
rect 22468 31288 22520 31340
rect 27804 31331 27856 31340
rect 27804 31297 27813 31331
rect 27813 31297 27847 31331
rect 27847 31297 27856 31331
rect 27804 31288 27856 31297
rect 17224 31220 17276 31272
rect 19248 31084 19300 31136
rect 20076 31084 20128 31136
rect 21916 31084 21968 31136
rect 23480 31084 23532 31136
rect 27988 31084 28040 31136
rect 5582 30982 5634 31034
rect 5646 30982 5698 31034
rect 5710 30982 5762 31034
rect 5774 30982 5826 31034
rect 5838 30982 5890 31034
rect 14846 30982 14898 31034
rect 14910 30982 14962 31034
rect 14974 30982 15026 31034
rect 15038 30982 15090 31034
rect 15102 30982 15154 31034
rect 24110 30982 24162 31034
rect 24174 30982 24226 31034
rect 24238 30982 24290 31034
rect 24302 30982 24354 31034
rect 24366 30982 24418 31034
rect 21364 30880 21416 30932
rect 19340 30812 19392 30864
rect 20904 30812 20956 30864
rect 22100 30812 22152 30864
rect 14372 30676 14424 30728
rect 17224 30676 17276 30728
rect 21916 30744 21968 30796
rect 27528 30787 27580 30796
rect 27528 30753 27537 30787
rect 27537 30753 27571 30787
rect 27571 30753 27580 30787
rect 27528 30744 27580 30753
rect 27988 30787 28040 30796
rect 27988 30753 27997 30787
rect 27997 30753 28031 30787
rect 28031 30753 28040 30787
rect 27988 30744 28040 30753
rect 28172 30787 28224 30796
rect 28172 30753 28181 30787
rect 28181 30753 28215 30787
rect 28215 30753 28224 30787
rect 28172 30744 28224 30753
rect 20812 30676 20864 30728
rect 24860 30676 24912 30728
rect 26148 30676 26200 30728
rect 14648 30651 14700 30660
rect 14648 30617 14657 30651
rect 14657 30617 14691 30651
rect 14691 30617 14700 30651
rect 14648 30608 14700 30617
rect 17316 30651 17368 30660
rect 17316 30617 17325 30651
rect 17325 30617 17359 30651
rect 17359 30617 17368 30651
rect 17316 30608 17368 30617
rect 19248 30651 19300 30660
rect 19248 30617 19257 30651
rect 19257 30617 19291 30651
rect 19291 30617 19300 30651
rect 19248 30608 19300 30617
rect 19984 30608 20036 30660
rect 20260 30608 20312 30660
rect 21640 30608 21692 30660
rect 15476 30583 15528 30592
rect 15476 30549 15485 30583
rect 15485 30549 15519 30583
rect 15519 30549 15528 30583
rect 15476 30540 15528 30549
rect 16672 30540 16724 30592
rect 25136 30540 25188 30592
rect 10214 30438 10266 30490
rect 10278 30438 10330 30490
rect 10342 30438 10394 30490
rect 10406 30438 10458 30490
rect 10470 30438 10522 30490
rect 19478 30438 19530 30490
rect 19542 30438 19594 30490
rect 19606 30438 19658 30490
rect 19670 30438 19722 30490
rect 19734 30438 19786 30490
rect 17316 30379 17368 30388
rect 17316 30345 17325 30379
rect 17325 30345 17359 30379
rect 17359 30345 17368 30379
rect 17316 30336 17368 30345
rect 19984 30336 20036 30388
rect 22468 30379 22520 30388
rect 15476 30268 15528 30320
rect 17776 30268 17828 30320
rect 22468 30345 22477 30379
rect 22477 30345 22511 30379
rect 22511 30345 22520 30379
rect 22468 30336 22520 30345
rect 1400 30243 1452 30252
rect 1400 30209 1409 30243
rect 1409 30209 1443 30243
rect 1443 30209 1452 30243
rect 1400 30200 1452 30209
rect 16672 30243 16724 30252
rect 16672 30209 16681 30243
rect 16681 30209 16715 30243
rect 16715 30209 16724 30243
rect 16672 30200 16724 30209
rect 19340 30200 19392 30252
rect 14004 30132 14056 30184
rect 17868 30175 17920 30184
rect 17868 30141 17877 30175
rect 17877 30141 17911 30175
rect 17911 30141 17920 30175
rect 18972 30175 19024 30184
rect 17868 30132 17920 30141
rect 18972 30141 18981 30175
rect 18981 30141 19015 30175
rect 19015 30141 19024 30175
rect 18972 30132 19024 30141
rect 19800 30243 19852 30252
rect 19800 30209 19809 30243
rect 19809 30209 19843 30243
rect 19843 30209 19852 30243
rect 19800 30200 19852 30209
rect 20168 30200 20220 30252
rect 20260 30200 20312 30252
rect 20812 30243 20864 30252
rect 20812 30209 20818 30243
rect 20818 30209 20852 30243
rect 20852 30209 20864 30243
rect 20812 30200 20864 30209
rect 21824 30243 21876 30252
rect 21364 30132 21416 30184
rect 19064 30064 19116 30116
rect 20812 30064 20864 30116
rect 14556 29996 14608 30048
rect 16120 29996 16172 30048
rect 16948 29996 17000 30048
rect 19340 29996 19392 30048
rect 21824 30209 21833 30243
rect 21833 30209 21867 30243
rect 21867 30209 21876 30243
rect 21824 30200 21876 30209
rect 22008 30243 22060 30252
rect 22008 30209 22017 30243
rect 22017 30209 22051 30243
rect 22051 30209 22060 30243
rect 22008 30200 22060 30209
rect 25136 30243 25188 30252
rect 25136 30209 25170 30243
rect 25170 30209 25188 30243
rect 21916 30132 21968 30184
rect 21732 30064 21784 30116
rect 25136 30200 25188 30209
rect 26976 30200 27028 30252
rect 27620 30200 27672 30252
rect 27804 30200 27856 30252
rect 23480 30064 23532 30116
rect 24032 30064 24084 30116
rect 26148 29996 26200 30048
rect 26516 29996 26568 30048
rect 28540 29996 28592 30048
rect 5582 29894 5634 29946
rect 5646 29894 5698 29946
rect 5710 29894 5762 29946
rect 5774 29894 5826 29946
rect 5838 29894 5890 29946
rect 14846 29894 14898 29946
rect 14910 29894 14962 29946
rect 14974 29894 15026 29946
rect 15038 29894 15090 29946
rect 15102 29894 15154 29946
rect 24110 29894 24162 29946
rect 24174 29894 24226 29946
rect 24238 29894 24290 29946
rect 24302 29894 24354 29946
rect 24366 29894 24418 29946
rect 14648 29792 14700 29844
rect 16580 29792 16632 29844
rect 17868 29792 17920 29844
rect 20168 29792 20220 29844
rect 22008 29792 22060 29844
rect 14464 29724 14516 29776
rect 14556 29656 14608 29708
rect 20812 29724 20864 29776
rect 21456 29724 21508 29776
rect 20996 29656 21048 29708
rect 21824 29699 21876 29708
rect 21824 29665 21833 29699
rect 21833 29665 21867 29699
rect 21867 29665 21876 29699
rect 21824 29656 21876 29665
rect 23020 29656 23072 29708
rect 14004 29520 14056 29572
rect 16948 29588 17000 29640
rect 19248 29631 19300 29640
rect 16120 29452 16172 29504
rect 19248 29597 19257 29631
rect 19257 29597 19291 29631
rect 19291 29597 19300 29631
rect 19248 29588 19300 29597
rect 19340 29588 19392 29640
rect 19800 29588 19852 29640
rect 20444 29588 20496 29640
rect 21456 29588 21508 29640
rect 21732 29588 21784 29640
rect 22560 29631 22612 29640
rect 22560 29597 22569 29631
rect 22569 29597 22603 29631
rect 22603 29597 22612 29631
rect 22560 29588 22612 29597
rect 23112 29588 23164 29640
rect 23664 29656 23716 29708
rect 26516 29699 26568 29708
rect 26516 29665 26525 29699
rect 26525 29665 26559 29699
rect 26559 29665 26568 29699
rect 26516 29656 26568 29665
rect 28724 29656 28776 29708
rect 17776 29452 17828 29504
rect 20168 29452 20220 29504
rect 23572 29631 23624 29640
rect 23572 29597 23581 29631
rect 23581 29597 23615 29631
rect 23615 29597 23624 29631
rect 23572 29588 23624 29597
rect 24032 29588 24084 29640
rect 25688 29520 25740 29572
rect 26148 29520 26200 29572
rect 10214 29350 10266 29402
rect 10278 29350 10330 29402
rect 10342 29350 10394 29402
rect 10406 29350 10458 29402
rect 10470 29350 10522 29402
rect 19478 29350 19530 29402
rect 19542 29350 19594 29402
rect 19606 29350 19658 29402
rect 19670 29350 19722 29402
rect 19734 29350 19786 29402
rect 19064 29248 19116 29300
rect 27344 29155 27396 29164
rect 27344 29121 27353 29155
rect 27353 29121 27387 29155
rect 27387 29121 27396 29155
rect 27344 29112 27396 29121
rect 13360 28976 13412 29028
rect 16580 28976 16632 29028
rect 27988 28951 28040 28960
rect 27988 28917 27997 28951
rect 27997 28917 28031 28951
rect 28031 28917 28040 28951
rect 27988 28908 28040 28917
rect 5582 28806 5634 28858
rect 5646 28806 5698 28858
rect 5710 28806 5762 28858
rect 5774 28806 5826 28858
rect 5838 28806 5890 28858
rect 14846 28806 14898 28858
rect 14910 28806 14962 28858
rect 14974 28806 15026 28858
rect 15038 28806 15090 28858
rect 15102 28806 15154 28858
rect 24110 28806 24162 28858
rect 24174 28806 24226 28858
rect 24238 28806 24290 28858
rect 24302 28806 24354 28858
rect 24366 28806 24418 28858
rect 21824 28747 21876 28756
rect 21824 28713 21833 28747
rect 21833 28713 21867 28747
rect 21867 28713 21876 28747
rect 21824 28704 21876 28713
rect 23664 28704 23716 28756
rect 17868 28636 17920 28688
rect 27528 28611 27580 28620
rect 27528 28577 27537 28611
rect 27537 28577 27571 28611
rect 27571 28577 27580 28611
rect 27528 28568 27580 28577
rect 27988 28568 28040 28620
rect 21456 28500 21508 28552
rect 22100 28500 22152 28552
rect 22744 28500 22796 28552
rect 23296 28500 23348 28552
rect 14188 28475 14240 28484
rect 14188 28441 14197 28475
rect 14197 28441 14231 28475
rect 14231 28441 14240 28475
rect 14188 28432 14240 28441
rect 14372 28475 14424 28484
rect 14372 28441 14381 28475
rect 14381 28441 14415 28475
rect 14415 28441 14424 28475
rect 14372 28432 14424 28441
rect 17592 28432 17644 28484
rect 27344 28432 27396 28484
rect 13820 28364 13872 28416
rect 18512 28364 18564 28416
rect 22560 28407 22612 28416
rect 22560 28373 22569 28407
rect 22569 28373 22603 28407
rect 22603 28373 22612 28407
rect 22560 28364 22612 28373
rect 22652 28364 22704 28416
rect 23296 28364 23348 28416
rect 10214 28262 10266 28314
rect 10278 28262 10330 28314
rect 10342 28262 10394 28314
rect 10406 28262 10458 28314
rect 10470 28262 10522 28314
rect 19478 28262 19530 28314
rect 19542 28262 19594 28314
rect 19606 28262 19658 28314
rect 19670 28262 19722 28314
rect 19734 28262 19786 28314
rect 20720 28203 20772 28212
rect 1400 28067 1452 28076
rect 1400 28033 1409 28067
rect 1409 28033 1443 28067
rect 1443 28033 1452 28067
rect 1400 28024 1452 28033
rect 14648 28092 14700 28144
rect 15752 28135 15804 28144
rect 15752 28101 15761 28135
rect 15761 28101 15795 28135
rect 15795 28101 15804 28135
rect 15752 28092 15804 28101
rect 13636 28067 13688 28076
rect 13636 28033 13670 28067
rect 13670 28033 13688 28067
rect 13636 28024 13688 28033
rect 20720 28169 20729 28203
rect 20729 28169 20763 28203
rect 20763 28169 20772 28203
rect 20720 28160 20772 28169
rect 22100 28203 22152 28212
rect 22100 28169 22109 28203
rect 22109 28169 22143 28203
rect 22143 28169 22152 28203
rect 22100 28160 22152 28169
rect 18052 28024 18104 28076
rect 18512 28067 18564 28076
rect 18512 28033 18521 28067
rect 18521 28033 18555 28067
rect 18555 28033 18564 28067
rect 18512 28024 18564 28033
rect 18604 28067 18656 28076
rect 18604 28033 18613 28067
rect 18613 28033 18647 28067
rect 18647 28033 18656 28067
rect 21824 28092 21876 28144
rect 27344 28203 27396 28212
rect 27344 28169 27353 28203
rect 27353 28169 27387 28203
rect 27387 28169 27396 28203
rect 27344 28160 27396 28169
rect 22560 28092 22612 28144
rect 18604 28024 18656 28033
rect 20168 28067 20220 28076
rect 20168 28033 20177 28067
rect 20177 28033 20211 28067
rect 20211 28033 20220 28067
rect 20168 28024 20220 28033
rect 20536 28067 20588 28076
rect 20536 28033 20545 28067
rect 20545 28033 20579 28067
rect 20579 28033 20588 28067
rect 20536 28024 20588 28033
rect 16764 27956 16816 28008
rect 17776 27956 17828 28008
rect 20812 28024 20864 28076
rect 22376 28067 22428 28076
rect 22376 28033 22385 28067
rect 22385 28033 22419 28067
rect 22419 28033 22428 28067
rect 22376 28024 22428 28033
rect 23020 28067 23072 28076
rect 23020 28033 23029 28067
rect 23029 28033 23063 28067
rect 23063 28033 23072 28067
rect 23020 28024 23072 28033
rect 23204 28067 23256 28076
rect 23204 28033 23213 28067
rect 23213 28033 23247 28067
rect 23247 28033 23256 28067
rect 23204 28024 23256 28033
rect 23572 28024 23624 28076
rect 27252 28067 27304 28076
rect 27252 28033 27261 28067
rect 27261 28033 27295 28067
rect 27295 28033 27304 28067
rect 27252 28024 27304 28033
rect 21824 27956 21876 28008
rect 24032 27956 24084 28008
rect 17684 27931 17736 27940
rect 17684 27897 17693 27931
rect 17693 27897 17727 27931
rect 17727 27897 17736 27931
rect 17684 27888 17736 27897
rect 14004 27820 14056 27872
rect 14740 27863 14792 27872
rect 14740 27829 14749 27863
rect 14749 27829 14783 27863
rect 14783 27829 14792 27863
rect 14740 27820 14792 27829
rect 15936 27863 15988 27872
rect 15936 27829 15945 27863
rect 15945 27829 15979 27863
rect 15979 27829 15988 27863
rect 15936 27820 15988 27829
rect 16672 27863 16724 27872
rect 16672 27829 16681 27863
rect 16681 27829 16715 27863
rect 16715 27829 16724 27863
rect 16672 27820 16724 27829
rect 18052 27820 18104 27872
rect 18328 27863 18380 27872
rect 18328 27829 18337 27863
rect 18337 27829 18371 27863
rect 18371 27829 18380 27863
rect 18328 27820 18380 27829
rect 18788 27863 18840 27872
rect 18788 27829 18797 27863
rect 18797 27829 18831 27863
rect 18831 27829 18840 27863
rect 18788 27820 18840 27829
rect 19248 27863 19300 27872
rect 19248 27829 19257 27863
rect 19257 27829 19291 27863
rect 19291 27829 19300 27863
rect 19248 27820 19300 27829
rect 22560 27820 22612 27872
rect 28172 27820 28224 27872
rect 5582 27718 5634 27770
rect 5646 27718 5698 27770
rect 5710 27718 5762 27770
rect 5774 27718 5826 27770
rect 5838 27718 5890 27770
rect 14846 27718 14898 27770
rect 14910 27718 14962 27770
rect 14974 27718 15026 27770
rect 15038 27718 15090 27770
rect 15102 27718 15154 27770
rect 24110 27718 24162 27770
rect 24174 27718 24226 27770
rect 24238 27718 24290 27770
rect 24302 27718 24354 27770
rect 24366 27718 24418 27770
rect 13636 27616 13688 27668
rect 14188 27659 14240 27668
rect 14188 27625 14197 27659
rect 14197 27625 14231 27659
rect 14231 27625 14240 27659
rect 14188 27616 14240 27625
rect 23204 27616 23256 27668
rect 13912 27548 13964 27600
rect 14464 27548 14516 27600
rect 14648 27523 14700 27532
rect 14648 27489 14657 27523
rect 14657 27489 14691 27523
rect 14691 27489 14700 27523
rect 14648 27480 14700 27489
rect 17316 27548 17368 27600
rect 20076 27548 20128 27600
rect 21364 27548 21416 27600
rect 21640 27591 21692 27600
rect 21640 27557 21649 27591
rect 21649 27557 21683 27591
rect 21683 27557 21692 27591
rect 21640 27548 21692 27557
rect 23112 27548 23164 27600
rect 17868 27480 17920 27532
rect 20536 27480 20588 27532
rect 13820 27412 13872 27464
rect 14004 27412 14056 27464
rect 15108 27412 15160 27464
rect 16672 27412 16724 27464
rect 20168 27412 20220 27464
rect 20444 27455 20496 27464
rect 20444 27421 20453 27455
rect 20453 27421 20487 27455
rect 20487 27421 20496 27455
rect 20444 27412 20496 27421
rect 20720 27480 20772 27532
rect 27528 27523 27580 27532
rect 27528 27489 27537 27523
rect 27537 27489 27571 27523
rect 27571 27489 27580 27523
rect 27528 27480 27580 27489
rect 28172 27523 28224 27532
rect 28172 27489 28181 27523
rect 28181 27489 28215 27523
rect 28215 27489 28224 27523
rect 28172 27480 28224 27489
rect 22376 27412 22428 27464
rect 22652 27412 22704 27464
rect 23388 27412 23440 27464
rect 23848 27412 23900 27464
rect 14372 27344 14424 27396
rect 14096 27276 14148 27328
rect 14740 27276 14792 27328
rect 21364 27344 21416 27396
rect 21640 27344 21692 27396
rect 27712 27344 27764 27396
rect 20352 27276 20404 27328
rect 21548 27276 21600 27328
rect 23296 27276 23348 27328
rect 10214 27174 10266 27226
rect 10278 27174 10330 27226
rect 10342 27174 10394 27226
rect 10406 27174 10458 27226
rect 10470 27174 10522 27226
rect 19478 27174 19530 27226
rect 19542 27174 19594 27226
rect 19606 27174 19658 27226
rect 19670 27174 19722 27226
rect 19734 27174 19786 27226
rect 15936 27072 15988 27124
rect 16764 27115 16816 27124
rect 16764 27081 16773 27115
rect 16773 27081 16807 27115
rect 16807 27081 16816 27115
rect 16764 27072 16816 27081
rect 18696 27072 18748 27124
rect 15108 27004 15160 27056
rect 15936 26979 15988 26988
rect 15936 26945 15945 26979
rect 15945 26945 15979 26979
rect 15979 26945 15988 26979
rect 15936 26936 15988 26945
rect 17316 26979 17368 26988
rect 15660 26868 15712 26920
rect 17316 26945 17325 26979
rect 17325 26945 17359 26979
rect 17359 26945 17368 26979
rect 17316 26936 17368 26945
rect 17868 26936 17920 26988
rect 18328 26936 18380 26988
rect 15936 26800 15988 26852
rect 18604 26936 18656 26988
rect 19156 26979 19208 26988
rect 19156 26945 19190 26979
rect 19190 26945 19208 26979
rect 20168 27072 20220 27124
rect 27712 27115 27764 27124
rect 21456 27004 21508 27056
rect 19156 26936 19208 26945
rect 22836 27004 22888 27056
rect 27712 27081 27721 27115
rect 27721 27081 27755 27115
rect 27755 27081 27764 27115
rect 27712 27072 27764 27081
rect 22192 26936 22244 26988
rect 22928 26979 22980 26988
rect 22928 26945 22937 26979
rect 22937 26945 22971 26979
rect 22971 26945 22980 26979
rect 22928 26936 22980 26945
rect 27896 26936 27948 26988
rect 17592 26843 17644 26852
rect 17592 26809 17601 26843
rect 17601 26809 17635 26843
rect 17635 26809 17644 26843
rect 17592 26800 17644 26809
rect 22744 26800 22796 26852
rect 18144 26732 18196 26784
rect 21916 26775 21968 26784
rect 21916 26741 21925 26775
rect 21925 26741 21959 26775
rect 21959 26741 21968 26775
rect 21916 26732 21968 26741
rect 23388 26732 23440 26784
rect 5582 26630 5634 26682
rect 5646 26630 5698 26682
rect 5710 26630 5762 26682
rect 5774 26630 5826 26682
rect 5838 26630 5890 26682
rect 14846 26630 14898 26682
rect 14910 26630 14962 26682
rect 14974 26630 15026 26682
rect 15038 26630 15090 26682
rect 15102 26630 15154 26682
rect 24110 26630 24162 26682
rect 24174 26630 24226 26682
rect 24238 26630 24290 26682
rect 24302 26630 24354 26682
rect 24366 26630 24418 26682
rect 18328 26528 18380 26580
rect 21548 26528 21600 26580
rect 23204 26528 23256 26580
rect 23848 26528 23900 26580
rect 17776 26503 17828 26512
rect 17776 26469 17785 26503
rect 17785 26469 17819 26503
rect 17819 26469 17828 26503
rect 17776 26460 17828 26469
rect 19064 26460 19116 26512
rect 23756 26460 23808 26512
rect 16488 26392 16540 26444
rect 17684 26392 17736 26444
rect 21548 26435 21600 26444
rect 14740 26367 14792 26376
rect 14740 26333 14749 26367
rect 14749 26333 14783 26367
rect 14783 26333 14792 26367
rect 14740 26324 14792 26333
rect 15568 26367 15620 26376
rect 15568 26333 15577 26367
rect 15577 26333 15611 26367
rect 15611 26333 15620 26367
rect 15568 26324 15620 26333
rect 15660 26324 15712 26376
rect 16580 26324 16632 26376
rect 19248 26367 19300 26376
rect 19248 26333 19257 26367
rect 19257 26333 19291 26367
rect 19291 26333 19300 26367
rect 19248 26324 19300 26333
rect 21548 26401 21557 26435
rect 21557 26401 21591 26435
rect 21591 26401 21600 26435
rect 21548 26392 21600 26401
rect 21916 26392 21968 26444
rect 15936 26256 15988 26308
rect 18512 26256 18564 26308
rect 19892 26324 19944 26376
rect 20352 26324 20404 26376
rect 21364 26367 21416 26376
rect 21364 26333 21373 26367
rect 21373 26333 21407 26367
rect 21407 26333 21416 26367
rect 21364 26324 21416 26333
rect 22744 26367 22796 26376
rect 20444 26256 20496 26308
rect 22744 26333 22753 26367
rect 22753 26333 22787 26367
rect 22787 26333 22796 26367
rect 22744 26324 22796 26333
rect 23204 26367 23256 26376
rect 23204 26333 23213 26367
rect 23213 26333 23247 26367
rect 23247 26333 23256 26367
rect 23204 26324 23256 26333
rect 23296 26367 23348 26376
rect 23296 26333 23305 26367
rect 23305 26333 23339 26367
rect 23339 26333 23348 26367
rect 23480 26367 23532 26376
rect 23296 26324 23348 26333
rect 23480 26333 23489 26367
rect 23489 26333 23523 26367
rect 23523 26333 23532 26367
rect 23480 26324 23532 26333
rect 24032 26324 24084 26376
rect 26424 26324 26476 26376
rect 28172 26324 28224 26376
rect 22836 26256 22888 26308
rect 14556 26231 14608 26240
rect 14556 26197 14565 26231
rect 14565 26197 14599 26231
rect 14599 26197 14608 26231
rect 14556 26188 14608 26197
rect 15384 26231 15436 26240
rect 15384 26197 15393 26231
rect 15393 26197 15427 26231
rect 15427 26197 15436 26231
rect 15384 26188 15436 26197
rect 22008 26188 22060 26240
rect 23296 26188 23348 26240
rect 23664 26231 23716 26240
rect 23664 26197 23673 26231
rect 23673 26197 23707 26231
rect 23707 26197 23716 26231
rect 23664 26188 23716 26197
rect 24492 26256 24544 26308
rect 25136 26188 25188 26240
rect 10214 26086 10266 26138
rect 10278 26086 10330 26138
rect 10342 26086 10394 26138
rect 10406 26086 10458 26138
rect 10470 26086 10522 26138
rect 19478 26086 19530 26138
rect 19542 26086 19594 26138
rect 19606 26086 19658 26138
rect 19670 26086 19722 26138
rect 19734 26086 19786 26138
rect 15568 25984 15620 26036
rect 19156 26027 19208 26036
rect 19156 25993 19165 26027
rect 19165 25993 19199 26027
rect 19199 25993 19208 26027
rect 19156 25984 19208 25993
rect 22744 25984 22796 26036
rect 14556 25916 14608 25968
rect 12532 25891 12584 25900
rect 12532 25857 12541 25891
rect 12541 25857 12575 25891
rect 12575 25857 12584 25891
rect 12532 25848 12584 25857
rect 12716 25891 12768 25900
rect 12716 25857 12725 25891
rect 12725 25857 12759 25891
rect 12759 25857 12768 25891
rect 12716 25848 12768 25857
rect 18788 25916 18840 25968
rect 18972 25916 19024 25968
rect 17868 25891 17920 25900
rect 17868 25857 17877 25891
rect 17877 25857 17911 25891
rect 17911 25857 17920 25891
rect 18144 25891 18196 25900
rect 17868 25848 17920 25857
rect 18144 25857 18153 25891
rect 18153 25857 18187 25891
rect 18187 25857 18196 25891
rect 18144 25848 18196 25857
rect 19064 25891 19116 25900
rect 19064 25857 19073 25891
rect 19073 25857 19107 25891
rect 19107 25857 19116 25891
rect 19064 25848 19116 25857
rect 19340 25848 19392 25900
rect 22560 25848 22612 25900
rect 23020 25848 23072 25900
rect 23664 25916 23716 25968
rect 23756 25916 23808 25968
rect 24952 25916 25004 25968
rect 26884 25916 26936 25968
rect 23388 25891 23440 25900
rect 23388 25857 23397 25891
rect 23397 25857 23431 25891
rect 23431 25857 23440 25891
rect 23388 25848 23440 25857
rect 23572 25848 23624 25900
rect 25136 25891 25188 25900
rect 14004 25823 14056 25832
rect 14004 25789 14013 25823
rect 14013 25789 14047 25823
rect 14047 25789 14056 25823
rect 14004 25780 14056 25789
rect 18052 25823 18104 25832
rect 18052 25789 18061 25823
rect 18061 25789 18095 25823
rect 18095 25789 18104 25823
rect 18052 25780 18104 25789
rect 22652 25780 22704 25832
rect 23204 25780 23256 25832
rect 25136 25857 25145 25891
rect 25145 25857 25179 25891
rect 25179 25857 25188 25891
rect 25136 25848 25188 25857
rect 24492 25755 24544 25764
rect 24492 25721 24501 25755
rect 24501 25721 24535 25755
rect 24535 25721 24544 25755
rect 24492 25712 24544 25721
rect 24676 25712 24728 25764
rect 1400 25644 1452 25696
rect 13268 25644 13320 25696
rect 17776 25644 17828 25696
rect 24952 25644 25004 25696
rect 27988 25644 28040 25696
rect 5582 25542 5634 25594
rect 5646 25542 5698 25594
rect 5710 25542 5762 25594
rect 5774 25542 5826 25594
rect 5838 25542 5890 25594
rect 14846 25542 14898 25594
rect 14910 25542 14962 25594
rect 14974 25542 15026 25594
rect 15038 25542 15090 25594
rect 15102 25542 15154 25594
rect 24110 25542 24162 25594
rect 24174 25542 24226 25594
rect 24238 25542 24290 25594
rect 24302 25542 24354 25594
rect 24366 25542 24418 25594
rect 14740 25440 14792 25492
rect 15384 25440 15436 25492
rect 22192 25483 22244 25492
rect 22192 25449 22201 25483
rect 22201 25449 22235 25483
rect 22235 25449 22244 25483
rect 22192 25440 22244 25449
rect 22928 25440 22980 25492
rect 23572 25440 23624 25492
rect 16488 25415 16540 25424
rect 16488 25381 16497 25415
rect 16497 25381 16531 25415
rect 16531 25381 16540 25415
rect 16488 25372 16540 25381
rect 1400 25347 1452 25356
rect 1400 25313 1409 25347
rect 1409 25313 1443 25347
rect 1443 25313 1452 25347
rect 1400 25304 1452 25313
rect 2780 25347 2832 25356
rect 2780 25313 2789 25347
rect 2789 25313 2823 25347
rect 2823 25313 2832 25347
rect 2780 25304 2832 25313
rect 14004 25304 14056 25356
rect 5540 25279 5592 25288
rect 5540 25245 5549 25279
rect 5549 25245 5583 25279
rect 5583 25245 5592 25279
rect 5540 25236 5592 25245
rect 13268 25279 13320 25288
rect 13268 25245 13286 25279
rect 13286 25245 13320 25279
rect 13268 25236 13320 25245
rect 15936 25236 15988 25288
rect 22744 25304 22796 25356
rect 22928 25347 22980 25356
rect 22928 25313 22937 25347
rect 22937 25313 22971 25347
rect 22971 25313 22980 25347
rect 23112 25347 23164 25356
rect 22928 25304 22980 25313
rect 23112 25313 23121 25347
rect 23121 25313 23155 25347
rect 23155 25313 23164 25347
rect 23112 25304 23164 25313
rect 23296 25304 23348 25356
rect 27528 25347 27580 25356
rect 1584 25211 1636 25220
rect 1584 25177 1593 25211
rect 1593 25177 1627 25211
rect 1627 25177 1636 25211
rect 1584 25168 1636 25177
rect 4712 25168 4764 25220
rect 4988 25211 5040 25220
rect 4988 25177 4997 25211
rect 4997 25177 5031 25211
rect 5031 25177 5040 25211
rect 4988 25168 5040 25177
rect 15752 25168 15804 25220
rect 16028 25168 16080 25220
rect 23756 25236 23808 25288
rect 27528 25313 27537 25347
rect 27537 25313 27571 25347
rect 27571 25313 27580 25347
rect 27528 25304 27580 25313
rect 27988 25347 28040 25356
rect 27988 25313 27997 25347
rect 27997 25313 28031 25347
rect 28031 25313 28040 25347
rect 27988 25304 28040 25313
rect 28172 25347 28224 25356
rect 28172 25313 28181 25347
rect 28181 25313 28215 25347
rect 28215 25313 28224 25347
rect 28172 25304 28224 25313
rect 24032 25236 24084 25288
rect 23480 25168 23532 25220
rect 24952 25168 25004 25220
rect 12164 25143 12216 25152
rect 12164 25109 12173 25143
rect 12173 25109 12207 25143
rect 12207 25109 12216 25143
rect 12164 25100 12216 25109
rect 15200 25100 15252 25152
rect 15476 25100 15528 25152
rect 16212 25143 16264 25152
rect 16212 25109 16221 25143
rect 16221 25109 16255 25143
rect 16255 25109 16264 25143
rect 16212 25100 16264 25109
rect 23940 25100 23992 25152
rect 10214 24998 10266 25050
rect 10278 24998 10330 25050
rect 10342 24998 10394 25050
rect 10406 24998 10458 25050
rect 10470 24998 10522 25050
rect 19478 24998 19530 25050
rect 19542 24998 19594 25050
rect 19606 24998 19658 25050
rect 19670 24998 19722 25050
rect 19734 24998 19786 25050
rect 1584 24896 1636 24948
rect 12532 24896 12584 24948
rect 15200 24896 15252 24948
rect 17868 24896 17920 24948
rect 12164 24828 12216 24880
rect 1768 24760 1820 24812
rect 5540 24760 5592 24812
rect 5908 24760 5960 24812
rect 15476 24803 15528 24812
rect 2044 24692 2096 24744
rect 4068 24735 4120 24744
rect 4068 24701 4077 24735
rect 4077 24701 4111 24735
rect 4111 24701 4120 24735
rect 4068 24692 4120 24701
rect 13176 24735 13228 24744
rect 3148 24624 3200 24676
rect 13176 24701 13185 24735
rect 13185 24701 13219 24735
rect 13219 24701 13228 24735
rect 13176 24692 13228 24701
rect 13360 24735 13412 24744
rect 13360 24701 13369 24735
rect 13369 24701 13403 24735
rect 13403 24701 13412 24735
rect 13360 24692 13412 24701
rect 15476 24769 15485 24803
rect 15485 24769 15519 24803
rect 15519 24769 15528 24803
rect 15476 24760 15528 24769
rect 16672 24803 16724 24812
rect 16672 24769 16681 24803
rect 16681 24769 16715 24803
rect 16715 24769 16724 24803
rect 16672 24760 16724 24769
rect 17408 24760 17460 24812
rect 17684 24803 17736 24812
rect 17684 24769 17693 24803
rect 17693 24769 17727 24803
rect 17727 24769 17736 24803
rect 17684 24760 17736 24769
rect 17868 24760 17920 24812
rect 25044 24760 25096 24812
rect 26424 24803 26476 24812
rect 26424 24769 26433 24803
rect 26433 24769 26467 24803
rect 26467 24769 26476 24803
rect 26424 24760 26476 24769
rect 26792 24760 26844 24812
rect 16580 24692 16632 24744
rect 16948 24692 17000 24744
rect 17316 24692 17368 24744
rect 21824 24735 21876 24744
rect 21824 24701 21833 24735
rect 21833 24701 21867 24735
rect 21867 24701 21876 24735
rect 21824 24692 21876 24701
rect 22100 24735 22152 24744
rect 22100 24701 22109 24735
rect 22109 24701 22143 24735
rect 22143 24701 22152 24735
rect 25964 24735 26016 24744
rect 22100 24692 22152 24701
rect 25964 24701 25973 24735
rect 25973 24701 26007 24735
rect 26007 24701 26016 24735
rect 25964 24692 26016 24701
rect 1768 24556 1820 24608
rect 28264 24624 28316 24676
rect 16580 24556 16632 24608
rect 17316 24556 17368 24608
rect 18880 24556 18932 24608
rect 19984 24599 20036 24608
rect 19984 24565 19993 24599
rect 19993 24565 20027 24599
rect 20027 24565 20036 24599
rect 19984 24556 20036 24565
rect 27436 24556 27488 24608
rect 5582 24454 5634 24506
rect 5646 24454 5698 24506
rect 5710 24454 5762 24506
rect 5774 24454 5826 24506
rect 5838 24454 5890 24506
rect 14846 24454 14898 24506
rect 14910 24454 14962 24506
rect 14974 24454 15026 24506
rect 15038 24454 15090 24506
rect 15102 24454 15154 24506
rect 24110 24454 24162 24506
rect 24174 24454 24226 24506
rect 24238 24454 24290 24506
rect 24302 24454 24354 24506
rect 24366 24454 24418 24506
rect 16672 24395 16724 24404
rect 16672 24361 16681 24395
rect 16681 24361 16715 24395
rect 16715 24361 16724 24395
rect 16672 24352 16724 24361
rect 16212 24284 16264 24336
rect 19892 24352 19944 24404
rect 23020 24352 23072 24404
rect 24032 24216 24084 24268
rect 27528 24259 27580 24268
rect 27528 24225 27537 24259
rect 27537 24225 27571 24259
rect 27571 24225 27580 24259
rect 27528 24216 27580 24225
rect 1400 24191 1452 24200
rect 1400 24157 1409 24191
rect 1409 24157 1443 24191
rect 1443 24157 1452 24191
rect 1400 24148 1452 24157
rect 5908 24148 5960 24200
rect 12900 24148 12952 24200
rect 15292 24191 15344 24200
rect 15292 24157 15301 24191
rect 15301 24157 15335 24191
rect 15335 24157 15344 24191
rect 15292 24148 15344 24157
rect 16580 24191 16632 24200
rect 16580 24157 16589 24191
rect 16589 24157 16623 24191
rect 16623 24157 16632 24191
rect 16580 24148 16632 24157
rect 5448 24123 5500 24132
rect 5448 24089 5457 24123
rect 5457 24089 5491 24123
rect 5491 24089 5500 24123
rect 5448 24080 5500 24089
rect 16856 24080 16908 24132
rect 19064 24148 19116 24200
rect 21824 24148 21876 24200
rect 20260 24080 20312 24132
rect 22376 24123 22428 24132
rect 22376 24089 22385 24123
rect 22385 24089 22419 24123
rect 22419 24089 22428 24123
rect 22376 24080 22428 24089
rect 25044 24123 25096 24132
rect 25044 24089 25053 24123
rect 25053 24089 25087 24123
rect 25087 24089 25096 24123
rect 25044 24080 25096 24089
rect 25596 24080 25648 24132
rect 28172 24191 28224 24200
rect 28172 24157 28181 24191
rect 28181 24157 28215 24191
rect 28215 24157 28224 24191
rect 28172 24148 28224 24157
rect 27436 24080 27488 24132
rect 27988 24123 28040 24132
rect 27988 24089 27997 24123
rect 27997 24089 28031 24123
rect 28031 24089 28040 24123
rect 27988 24080 28040 24089
rect 1584 24055 1636 24064
rect 1584 24021 1593 24055
rect 1593 24021 1627 24055
rect 1627 24021 1636 24055
rect 1584 24012 1636 24021
rect 12440 24012 12492 24064
rect 15108 24055 15160 24064
rect 15108 24021 15117 24055
rect 15117 24021 15151 24055
rect 15151 24021 15160 24055
rect 15108 24012 15160 24021
rect 15660 24012 15712 24064
rect 16028 24012 16080 24064
rect 16764 24012 16816 24064
rect 17408 24012 17460 24064
rect 21456 24055 21508 24064
rect 21456 24021 21465 24055
rect 21465 24021 21499 24055
rect 21499 24021 21508 24055
rect 21456 24012 21508 24021
rect 10214 23910 10266 23962
rect 10278 23910 10330 23962
rect 10342 23910 10394 23962
rect 10406 23910 10458 23962
rect 10470 23910 10522 23962
rect 19478 23910 19530 23962
rect 19542 23910 19594 23962
rect 19606 23910 19658 23962
rect 19670 23910 19722 23962
rect 19734 23910 19786 23962
rect 1584 23808 1636 23860
rect 13176 23808 13228 23860
rect 17684 23808 17736 23860
rect 17868 23808 17920 23860
rect 21364 23808 21416 23860
rect 22376 23808 22428 23860
rect 2320 23740 2372 23792
rect 15108 23740 15160 23792
rect 5908 23672 5960 23724
rect 13544 23672 13596 23724
rect 9496 23604 9548 23656
rect 12808 23604 12860 23656
rect 13360 23604 13412 23656
rect 14740 23647 14792 23656
rect 14740 23613 14749 23647
rect 14749 23613 14783 23647
rect 14783 23613 14792 23647
rect 14740 23604 14792 23613
rect 3148 23468 3200 23520
rect 4160 23468 4212 23520
rect 12532 23468 12584 23520
rect 16580 23468 16632 23520
rect 16764 23672 16816 23724
rect 17132 23715 17184 23724
rect 17132 23681 17141 23715
rect 17141 23681 17175 23715
rect 17175 23681 17184 23715
rect 21732 23740 21784 23792
rect 21916 23740 21968 23792
rect 27620 23808 27672 23860
rect 27436 23783 27488 23792
rect 27436 23749 27445 23783
rect 27445 23749 27479 23783
rect 27479 23749 27488 23783
rect 27436 23740 27488 23749
rect 17132 23672 17184 23681
rect 19800 23672 19852 23724
rect 20812 23715 20864 23724
rect 20812 23681 20821 23715
rect 20821 23681 20855 23715
rect 20855 23681 20864 23715
rect 20812 23672 20864 23681
rect 21456 23672 21508 23724
rect 25596 23715 25648 23724
rect 25596 23681 25605 23715
rect 25605 23681 25639 23715
rect 25639 23681 25648 23715
rect 25596 23672 25648 23681
rect 20720 23604 20772 23656
rect 22008 23604 22060 23656
rect 20536 23536 20588 23588
rect 21824 23536 21876 23588
rect 25412 23604 25464 23656
rect 27068 23604 27120 23656
rect 18144 23468 18196 23520
rect 20076 23468 20128 23520
rect 21548 23468 21600 23520
rect 21640 23468 21692 23520
rect 22100 23468 22152 23520
rect 5582 23366 5634 23418
rect 5646 23366 5698 23418
rect 5710 23366 5762 23418
rect 5774 23366 5826 23418
rect 5838 23366 5890 23418
rect 14846 23366 14898 23418
rect 14910 23366 14962 23418
rect 14974 23366 15026 23418
rect 15038 23366 15090 23418
rect 15102 23366 15154 23418
rect 24110 23366 24162 23418
rect 24174 23366 24226 23418
rect 24238 23366 24290 23418
rect 24302 23366 24354 23418
rect 24366 23366 24418 23418
rect 13544 23307 13596 23316
rect 13544 23273 13553 23307
rect 13553 23273 13587 23307
rect 13587 23273 13596 23307
rect 13544 23264 13596 23273
rect 15292 23264 15344 23316
rect 16672 23264 16724 23316
rect 17684 23264 17736 23316
rect 19800 23264 19852 23316
rect 21088 23264 21140 23316
rect 21272 23264 21324 23316
rect 15660 23196 15712 23248
rect 18420 23239 18472 23248
rect 18420 23205 18429 23239
rect 18429 23205 18463 23239
rect 18463 23205 18472 23239
rect 18420 23196 18472 23205
rect 26976 23264 27028 23316
rect 27988 23307 28040 23316
rect 27988 23273 27997 23307
rect 27997 23273 28031 23307
rect 28031 23273 28040 23307
rect 27988 23264 28040 23273
rect 12164 23103 12216 23112
rect 12164 23069 12173 23103
rect 12173 23069 12207 23103
rect 12207 23069 12216 23103
rect 12164 23060 12216 23069
rect 12440 23103 12492 23112
rect 12440 23069 12474 23103
rect 12474 23069 12492 23103
rect 12440 23060 12492 23069
rect 14740 22992 14792 23044
rect 12624 22924 12676 22976
rect 16580 23103 16632 23112
rect 16580 23069 16589 23103
rect 16589 23069 16623 23103
rect 16623 23069 16632 23103
rect 16580 23060 16632 23069
rect 17132 23060 17184 23112
rect 18144 23103 18196 23112
rect 18144 23069 18153 23103
rect 18153 23069 18187 23103
rect 18187 23069 18196 23103
rect 18144 23060 18196 23069
rect 18972 23060 19024 23112
rect 20536 23128 20588 23180
rect 16764 23035 16816 23044
rect 16764 23001 16773 23035
rect 16773 23001 16807 23035
rect 16807 23001 16816 23035
rect 16764 22992 16816 23001
rect 16948 22992 17000 23044
rect 17316 23035 17368 23044
rect 17316 23001 17325 23035
rect 17325 23001 17359 23035
rect 17359 23001 17368 23035
rect 17316 22992 17368 23001
rect 17408 22992 17460 23044
rect 18788 22992 18840 23044
rect 18880 22992 18932 23044
rect 20444 23060 20496 23112
rect 20812 23128 20864 23180
rect 21456 23128 21508 23180
rect 21824 23128 21876 23180
rect 21456 23035 21508 23044
rect 21456 23001 21465 23035
rect 21465 23001 21499 23035
rect 21499 23001 21508 23035
rect 25228 23196 25280 23248
rect 27712 23196 27764 23248
rect 28448 23196 28500 23248
rect 23664 23171 23716 23180
rect 23664 23137 23673 23171
rect 23673 23137 23707 23171
rect 23707 23137 23716 23171
rect 23664 23128 23716 23137
rect 23388 23060 23440 23112
rect 25872 23128 25924 23180
rect 21456 22992 21508 23001
rect 21916 22992 21968 23044
rect 22560 22992 22612 23044
rect 24676 23103 24728 23112
rect 24676 23069 24685 23103
rect 24685 23069 24719 23103
rect 24719 23069 24728 23103
rect 24860 23103 24912 23112
rect 24676 23060 24728 23069
rect 24860 23069 24869 23103
rect 24869 23069 24903 23103
rect 24903 23069 24912 23103
rect 24860 23060 24912 23069
rect 25596 23103 25648 23112
rect 25596 23069 25605 23103
rect 25605 23069 25639 23103
rect 25639 23069 25648 23103
rect 25596 23060 25648 23069
rect 26976 23060 27028 23112
rect 27344 23060 27396 23112
rect 28356 23060 28408 23112
rect 27712 22992 27764 23044
rect 17684 22967 17736 22976
rect 17684 22933 17693 22967
rect 17693 22933 17727 22967
rect 17727 22933 17736 22967
rect 17684 22924 17736 22933
rect 21088 22924 21140 22976
rect 21824 22967 21876 22976
rect 21824 22933 21833 22967
rect 21833 22933 21867 22967
rect 21867 22933 21876 22967
rect 21824 22924 21876 22933
rect 22744 22924 22796 22976
rect 23480 22967 23532 22976
rect 23480 22933 23489 22967
rect 23489 22933 23523 22967
rect 23523 22933 23532 22967
rect 23480 22924 23532 22933
rect 25136 22924 25188 22976
rect 10214 22822 10266 22874
rect 10278 22822 10330 22874
rect 10342 22822 10394 22874
rect 10406 22822 10458 22874
rect 10470 22822 10522 22874
rect 19478 22822 19530 22874
rect 19542 22822 19594 22874
rect 19606 22822 19658 22874
rect 19670 22822 19722 22874
rect 19734 22822 19786 22874
rect 2688 22720 2740 22772
rect 12624 22720 12676 22772
rect 12900 22763 12952 22772
rect 12900 22729 12909 22763
rect 12909 22729 12943 22763
rect 12943 22729 12952 22763
rect 12900 22720 12952 22729
rect 18972 22763 19024 22772
rect 18972 22729 18981 22763
rect 18981 22729 19015 22763
rect 19015 22729 19024 22763
rect 18972 22720 19024 22729
rect 20260 22763 20312 22772
rect 20260 22729 20269 22763
rect 20269 22729 20303 22763
rect 20303 22729 20312 22763
rect 20260 22720 20312 22729
rect 4712 22652 4764 22704
rect 12532 22695 12584 22704
rect 12532 22661 12541 22695
rect 12541 22661 12575 22695
rect 12575 22661 12584 22695
rect 12532 22652 12584 22661
rect 12716 22695 12768 22704
rect 12716 22661 12725 22695
rect 12725 22661 12759 22695
rect 12759 22661 12768 22695
rect 12716 22652 12768 22661
rect 23388 22720 23440 22772
rect 23480 22720 23532 22772
rect 24676 22720 24728 22772
rect 25136 22720 25188 22772
rect 21456 22652 21508 22704
rect 21916 22652 21968 22704
rect 14464 22627 14516 22636
rect 14464 22593 14482 22627
rect 14482 22593 14516 22627
rect 14464 22584 14516 22593
rect 14740 22627 14792 22636
rect 14740 22593 14749 22627
rect 14749 22593 14783 22627
rect 14783 22593 14792 22627
rect 14740 22584 14792 22593
rect 18880 22627 18932 22636
rect 18880 22593 18889 22627
rect 18889 22593 18923 22627
rect 18923 22593 18932 22627
rect 18880 22584 18932 22593
rect 18972 22584 19024 22636
rect 20076 22627 20128 22636
rect 20076 22593 20085 22627
rect 20085 22593 20119 22627
rect 20119 22593 20128 22627
rect 20076 22584 20128 22593
rect 20720 22516 20772 22568
rect 22928 22584 22980 22636
rect 25044 22584 25096 22636
rect 27712 22627 27764 22636
rect 27712 22593 27721 22627
rect 27721 22593 27755 22627
rect 27755 22593 27764 22627
rect 27712 22584 27764 22593
rect 25964 22448 26016 22500
rect 13360 22423 13412 22432
rect 13360 22389 13369 22423
rect 13369 22389 13403 22423
rect 13403 22389 13412 22423
rect 13360 22380 13412 22389
rect 22008 22423 22060 22432
rect 22008 22389 22017 22423
rect 22017 22389 22051 22423
rect 22051 22389 22060 22423
rect 22008 22380 22060 22389
rect 22192 22423 22244 22432
rect 22192 22389 22201 22423
rect 22201 22389 22235 22423
rect 22235 22389 22244 22423
rect 22192 22380 22244 22389
rect 26240 22380 26292 22432
rect 26516 22380 26568 22432
rect 5582 22278 5634 22330
rect 5646 22278 5698 22330
rect 5710 22278 5762 22330
rect 5774 22278 5826 22330
rect 5838 22278 5890 22330
rect 14846 22278 14898 22330
rect 14910 22278 14962 22330
rect 14974 22278 15026 22330
rect 15038 22278 15090 22330
rect 15102 22278 15154 22330
rect 24110 22278 24162 22330
rect 24174 22278 24226 22330
rect 24238 22278 24290 22330
rect 24302 22278 24354 22330
rect 24366 22278 24418 22330
rect 14464 22176 14516 22228
rect 22928 22219 22980 22228
rect 22928 22185 22937 22219
rect 22937 22185 22971 22219
rect 22971 22185 22980 22219
rect 22928 22176 22980 22185
rect 25044 22219 25096 22228
rect 25044 22185 25053 22219
rect 25053 22185 25087 22219
rect 25087 22185 25096 22219
rect 25044 22176 25096 22185
rect 25504 22108 25556 22160
rect 12716 22040 12768 22092
rect 17224 22040 17276 22092
rect 23664 22040 23716 22092
rect 26240 22108 26292 22160
rect 26516 22083 26568 22092
rect 26516 22049 26525 22083
rect 26525 22049 26559 22083
rect 26559 22049 26568 22083
rect 26516 22040 26568 22049
rect 28632 22040 28684 22092
rect 1584 22015 1636 22024
rect 1584 21981 1593 22015
rect 1593 21981 1627 22015
rect 1627 21981 1636 22015
rect 1584 21972 1636 21981
rect 14096 22015 14148 22024
rect 14096 21981 14105 22015
rect 14105 21981 14139 22015
rect 14139 21981 14148 22015
rect 14096 21972 14148 21981
rect 20168 21972 20220 22024
rect 20904 21972 20956 22024
rect 21640 21972 21692 22024
rect 22744 22015 22796 22024
rect 22744 21981 22753 22015
rect 22753 21981 22787 22015
rect 22787 21981 22796 22015
rect 22744 21972 22796 21981
rect 24584 22015 24636 22024
rect 24584 21981 24593 22015
rect 24593 21981 24627 22015
rect 24627 21981 24636 22015
rect 24584 21972 24636 21981
rect 25228 22015 25280 22024
rect 25228 21981 25237 22015
rect 25237 21981 25271 22015
rect 25271 21981 25280 22015
rect 25228 21972 25280 21981
rect 25320 21972 25372 22024
rect 21364 21904 21416 21956
rect 20812 21879 20864 21888
rect 20812 21845 20821 21879
rect 20821 21845 20855 21879
rect 20855 21845 20864 21879
rect 20812 21836 20864 21845
rect 10214 21734 10266 21786
rect 10278 21734 10330 21786
rect 10342 21734 10394 21786
rect 10406 21734 10458 21786
rect 10470 21734 10522 21786
rect 19478 21734 19530 21786
rect 19542 21734 19594 21786
rect 19606 21734 19658 21786
rect 19670 21734 19722 21786
rect 19734 21734 19786 21786
rect 17224 21675 17276 21684
rect 17224 21641 17233 21675
rect 17233 21641 17267 21675
rect 17267 21641 17276 21675
rect 17224 21632 17276 21641
rect 18144 21632 18196 21684
rect 18420 21632 18472 21684
rect 19340 21632 19392 21684
rect 16764 21564 16816 21616
rect 17684 21564 17736 21616
rect 19064 21607 19116 21616
rect 19064 21573 19073 21607
rect 19073 21573 19107 21607
rect 19107 21573 19116 21607
rect 19064 21564 19116 21573
rect 4712 21496 4764 21548
rect 13360 21496 13412 21548
rect 15384 21496 15436 21548
rect 15568 21539 15620 21548
rect 15568 21505 15577 21539
rect 15577 21505 15611 21539
rect 15611 21505 15620 21539
rect 15568 21496 15620 21505
rect 17316 21539 17368 21548
rect 17316 21505 17325 21539
rect 17325 21505 17359 21539
rect 17359 21505 17368 21539
rect 17316 21496 17368 21505
rect 18052 21496 18104 21548
rect 2044 21335 2096 21344
rect 2044 21301 2053 21335
rect 2053 21301 2087 21335
rect 2087 21301 2096 21335
rect 2044 21292 2096 21301
rect 14740 21292 14792 21344
rect 18512 21292 18564 21344
rect 18972 21335 19024 21344
rect 18972 21301 18981 21335
rect 18981 21301 19015 21335
rect 19015 21301 19024 21335
rect 18972 21292 19024 21301
rect 20168 21496 20220 21548
rect 21364 21632 21416 21684
rect 23664 21632 23716 21684
rect 20812 21564 20864 21616
rect 25964 21564 26016 21616
rect 20444 21539 20496 21548
rect 20444 21505 20453 21539
rect 20453 21505 20487 21539
rect 20487 21505 20496 21539
rect 20444 21496 20496 21505
rect 22008 21539 22060 21548
rect 22008 21505 22017 21539
rect 22017 21505 22051 21539
rect 22051 21505 22060 21539
rect 22008 21496 22060 21505
rect 22192 21539 22244 21548
rect 22192 21505 22201 21539
rect 22201 21505 22235 21539
rect 22235 21505 22244 21539
rect 22192 21496 22244 21505
rect 27712 21539 27764 21548
rect 27712 21505 27721 21539
rect 27721 21505 27755 21539
rect 27755 21505 27764 21539
rect 27712 21496 27764 21505
rect 22284 21471 22336 21480
rect 22284 21437 22293 21471
rect 22293 21437 22327 21471
rect 22327 21437 22336 21471
rect 22284 21428 22336 21437
rect 26148 21471 26200 21480
rect 26148 21437 26157 21471
rect 26157 21437 26191 21471
rect 26191 21437 26200 21471
rect 26148 21428 26200 21437
rect 24860 21360 24912 21412
rect 20812 21292 20864 21344
rect 21732 21292 21784 21344
rect 26516 21292 26568 21344
rect 5582 21190 5634 21242
rect 5646 21190 5698 21242
rect 5710 21190 5762 21242
rect 5774 21190 5826 21242
rect 5838 21190 5890 21242
rect 14846 21190 14898 21242
rect 14910 21190 14962 21242
rect 14974 21190 15026 21242
rect 15038 21190 15090 21242
rect 15102 21190 15154 21242
rect 24110 21190 24162 21242
rect 24174 21190 24226 21242
rect 24238 21190 24290 21242
rect 24302 21190 24354 21242
rect 24366 21190 24418 21242
rect 14740 21088 14792 21140
rect 16764 21088 16816 21140
rect 19064 21088 19116 21140
rect 14096 21020 14148 21072
rect 1584 20952 1636 21004
rect 14280 20927 14332 20936
rect 14280 20893 14289 20927
rect 14289 20893 14323 20927
rect 14323 20893 14332 20927
rect 14280 20884 14332 20893
rect 18512 20952 18564 21004
rect 16028 20884 16080 20936
rect 16856 20884 16908 20936
rect 17776 20884 17828 20936
rect 18052 20927 18104 20936
rect 18052 20893 18061 20927
rect 18061 20893 18095 20927
rect 18095 20893 18104 20927
rect 18052 20884 18104 20893
rect 18144 20927 18196 20936
rect 18144 20893 18153 20927
rect 18153 20893 18187 20927
rect 18187 20893 18196 20927
rect 18144 20884 18196 20893
rect 18788 20884 18840 20936
rect 23204 20952 23256 21004
rect 25320 20995 25372 21004
rect 25320 20961 25329 20995
rect 25329 20961 25363 20995
rect 25363 20961 25372 20995
rect 25320 20952 25372 20961
rect 25504 20952 25556 21004
rect 26516 20995 26568 21004
rect 26516 20961 26525 20995
rect 26525 20961 26559 20995
rect 26559 20961 26568 20995
rect 26516 20952 26568 20961
rect 28172 20995 28224 21004
rect 28172 20961 28181 20995
rect 28181 20961 28215 20995
rect 28215 20961 28224 20995
rect 28172 20952 28224 20961
rect 2044 20816 2096 20868
rect 3700 20816 3752 20868
rect 12072 20859 12124 20868
rect 12072 20825 12081 20859
rect 12081 20825 12115 20859
rect 12115 20825 12124 20859
rect 12072 20816 12124 20825
rect 12716 20816 12768 20868
rect 15476 20816 15528 20868
rect 15752 20816 15804 20868
rect 18696 20816 18748 20868
rect 20444 20884 20496 20936
rect 21088 20884 21140 20936
rect 21456 20927 21508 20936
rect 21456 20893 21465 20927
rect 21465 20893 21499 20927
rect 21499 20893 21508 20927
rect 21456 20884 21508 20893
rect 21732 20927 21784 20936
rect 21732 20893 21766 20927
rect 21766 20893 21784 20927
rect 21732 20884 21784 20893
rect 23572 20884 23624 20936
rect 12624 20748 12676 20800
rect 14096 20791 14148 20800
rect 14096 20757 14105 20791
rect 14105 20757 14139 20791
rect 14139 20757 14148 20791
rect 14096 20748 14148 20757
rect 14740 20748 14792 20800
rect 15292 20748 15344 20800
rect 17316 20748 17368 20800
rect 20168 20748 20220 20800
rect 22468 20748 22520 20800
rect 22836 20791 22888 20800
rect 22836 20757 22845 20791
rect 22845 20757 22879 20791
rect 22879 20757 22888 20791
rect 22836 20748 22888 20757
rect 23756 20748 23808 20800
rect 24492 20748 24544 20800
rect 25136 20791 25188 20800
rect 25136 20757 25145 20791
rect 25145 20757 25179 20791
rect 25179 20757 25188 20791
rect 25136 20748 25188 20757
rect 10214 20646 10266 20698
rect 10278 20646 10330 20698
rect 10342 20646 10394 20698
rect 10406 20646 10458 20698
rect 10470 20646 10522 20698
rect 19478 20646 19530 20698
rect 19542 20646 19594 20698
rect 19606 20646 19658 20698
rect 19670 20646 19722 20698
rect 19734 20646 19786 20698
rect 18420 20544 18472 20596
rect 18696 20587 18748 20596
rect 18696 20553 18705 20587
rect 18705 20553 18739 20587
rect 18739 20553 18748 20587
rect 18696 20544 18748 20553
rect 21088 20587 21140 20596
rect 21088 20553 21097 20587
rect 21097 20553 21131 20587
rect 21131 20553 21140 20587
rect 21088 20544 21140 20553
rect 22836 20544 22888 20596
rect 26148 20544 26200 20596
rect 2320 20383 2372 20392
rect 2320 20349 2329 20383
rect 2329 20349 2363 20383
rect 2363 20349 2372 20383
rect 2320 20340 2372 20349
rect 2872 20340 2924 20392
rect 2964 20383 3016 20392
rect 2964 20349 2973 20383
rect 2973 20349 3007 20383
rect 3007 20349 3016 20383
rect 2964 20340 3016 20349
rect 11888 20340 11940 20392
rect 12164 20476 12216 20528
rect 14096 20519 14148 20528
rect 12624 20408 12676 20460
rect 14096 20485 14130 20519
rect 14130 20485 14148 20519
rect 14096 20476 14148 20485
rect 15568 20408 15620 20460
rect 16856 20476 16908 20528
rect 20812 20476 20864 20528
rect 20996 20476 21048 20528
rect 21456 20476 21508 20528
rect 23756 20519 23808 20528
rect 23756 20485 23790 20519
rect 23790 20485 23808 20519
rect 23756 20476 23808 20485
rect 15936 20408 15988 20460
rect 18512 20451 18564 20460
rect 18512 20417 18521 20451
rect 18521 20417 18555 20451
rect 18555 20417 18564 20451
rect 18512 20408 18564 20417
rect 18788 20451 18840 20460
rect 18788 20417 18797 20451
rect 18797 20417 18831 20451
rect 18831 20417 18840 20451
rect 18788 20408 18840 20417
rect 23480 20451 23532 20460
rect 22468 20383 22520 20392
rect 14096 20204 14148 20256
rect 15200 20247 15252 20256
rect 15200 20213 15209 20247
rect 15209 20213 15243 20247
rect 15243 20213 15252 20247
rect 15200 20204 15252 20213
rect 15384 20204 15436 20256
rect 15752 20204 15804 20256
rect 16028 20247 16080 20256
rect 16028 20213 16037 20247
rect 16037 20213 16071 20247
rect 16071 20213 16080 20247
rect 16028 20204 16080 20213
rect 17684 20204 17736 20256
rect 22468 20349 22477 20383
rect 22477 20349 22511 20383
rect 22511 20349 22520 20383
rect 22468 20340 22520 20349
rect 23480 20417 23489 20451
rect 23489 20417 23523 20451
rect 23523 20417 23532 20451
rect 23480 20408 23532 20417
rect 20720 20204 20772 20256
rect 20996 20204 21048 20256
rect 23388 20204 23440 20256
rect 27344 20451 27396 20460
rect 27344 20417 27353 20451
rect 27353 20417 27387 20451
rect 27387 20417 27396 20451
rect 27344 20408 27396 20417
rect 28080 20451 28132 20460
rect 28080 20417 28089 20451
rect 28089 20417 28123 20451
rect 28123 20417 28132 20451
rect 28080 20408 28132 20417
rect 24952 20340 25004 20392
rect 25688 20340 25740 20392
rect 25412 20247 25464 20256
rect 25412 20213 25421 20247
rect 25421 20213 25455 20247
rect 25455 20213 25464 20247
rect 25412 20204 25464 20213
rect 26516 20204 26568 20256
rect 5582 20102 5634 20154
rect 5646 20102 5698 20154
rect 5710 20102 5762 20154
rect 5774 20102 5826 20154
rect 5838 20102 5890 20154
rect 14846 20102 14898 20154
rect 14910 20102 14962 20154
rect 14974 20102 15026 20154
rect 15038 20102 15090 20154
rect 15102 20102 15154 20154
rect 24110 20102 24162 20154
rect 24174 20102 24226 20154
rect 24238 20102 24290 20154
rect 24302 20102 24354 20154
rect 24366 20102 24418 20154
rect 2320 20043 2372 20052
rect 2320 20009 2329 20043
rect 2329 20009 2363 20043
rect 2363 20009 2372 20043
rect 2320 20000 2372 20009
rect 2872 20043 2924 20052
rect 2872 20009 2881 20043
rect 2881 20009 2915 20043
rect 2915 20009 2924 20043
rect 2872 20000 2924 20009
rect 12072 20000 12124 20052
rect 14280 20000 14332 20052
rect 15292 20000 15344 20052
rect 21364 20043 21416 20052
rect 21364 20009 21373 20043
rect 21373 20009 21407 20043
rect 21407 20009 21416 20043
rect 21364 20000 21416 20009
rect 22284 20043 22336 20052
rect 22284 20009 22293 20043
rect 22293 20009 22327 20043
rect 22327 20009 22336 20043
rect 22284 20000 22336 20009
rect 23572 20043 23624 20052
rect 23572 20009 23581 20043
rect 23581 20009 23615 20043
rect 23615 20009 23624 20043
rect 23572 20000 23624 20009
rect 25136 20000 25188 20052
rect 16672 19932 16724 19984
rect 18972 19932 19024 19984
rect 22192 19932 22244 19984
rect 12808 19907 12860 19916
rect 12808 19873 12817 19907
rect 12817 19873 12851 19907
rect 12851 19873 12860 19907
rect 12808 19864 12860 19873
rect 1400 19796 1452 19848
rect 4160 19796 4212 19848
rect 14188 19839 14240 19848
rect 14188 19805 14197 19839
rect 14197 19805 14231 19839
rect 14231 19805 14240 19839
rect 14188 19796 14240 19805
rect 14740 19796 14792 19848
rect 14096 19728 14148 19780
rect 2964 19660 3016 19712
rect 12716 19703 12768 19712
rect 12716 19669 12725 19703
rect 12725 19669 12759 19703
rect 12759 19669 12768 19703
rect 15476 19864 15528 19916
rect 15844 19864 15896 19916
rect 15384 19728 15436 19780
rect 15752 19839 15804 19848
rect 15752 19805 15761 19839
rect 15761 19805 15795 19839
rect 15795 19805 15804 19839
rect 15936 19839 15988 19848
rect 15752 19796 15804 19805
rect 15936 19805 15945 19839
rect 15945 19805 15979 19839
rect 15979 19805 15988 19839
rect 15936 19796 15988 19805
rect 17408 19796 17460 19848
rect 18328 19796 18380 19848
rect 20904 19796 20956 19848
rect 21088 19796 21140 19848
rect 22836 19864 22888 19916
rect 23480 19864 23532 19916
rect 26516 19907 26568 19916
rect 26516 19873 26525 19907
rect 26525 19873 26559 19907
rect 26559 19873 26568 19907
rect 26516 19864 26568 19873
rect 28172 19907 28224 19916
rect 28172 19873 28181 19907
rect 28181 19873 28215 19907
rect 28215 19873 28224 19907
rect 28172 19864 28224 19873
rect 22744 19796 22796 19848
rect 23388 19839 23440 19848
rect 12716 19660 12768 19669
rect 17316 19728 17368 19780
rect 17684 19771 17736 19780
rect 17684 19737 17693 19771
rect 17693 19737 17727 19771
rect 17727 19737 17736 19771
rect 17684 19728 17736 19737
rect 22192 19728 22244 19780
rect 22836 19728 22888 19780
rect 23388 19805 23397 19839
rect 23397 19805 23431 19839
rect 23431 19805 23440 19839
rect 23388 19796 23440 19805
rect 26332 19839 26384 19848
rect 26332 19805 26341 19839
rect 26341 19805 26375 19839
rect 26375 19805 26384 19839
rect 26332 19796 26384 19805
rect 24032 19728 24084 19780
rect 25136 19728 25188 19780
rect 22468 19660 22520 19712
rect 23664 19660 23716 19712
rect 10214 19558 10266 19610
rect 10278 19558 10330 19610
rect 10342 19558 10394 19610
rect 10406 19558 10458 19610
rect 10470 19558 10522 19610
rect 19478 19558 19530 19610
rect 19542 19558 19594 19610
rect 19606 19558 19658 19610
rect 19670 19558 19722 19610
rect 19734 19558 19786 19610
rect 25136 19499 25188 19508
rect 25136 19465 25145 19499
rect 25145 19465 25179 19499
rect 25179 19465 25188 19499
rect 25136 19456 25188 19465
rect 16856 19388 16908 19440
rect 17408 19388 17460 19440
rect 19984 19388 20036 19440
rect 1400 19363 1452 19372
rect 1400 19329 1409 19363
rect 1409 19329 1443 19363
rect 1443 19329 1452 19363
rect 1400 19320 1452 19329
rect 14280 19320 14332 19372
rect 15200 19320 15252 19372
rect 24492 19363 24544 19372
rect 24492 19329 24501 19363
rect 24501 19329 24535 19363
rect 24535 19329 24544 19363
rect 24492 19320 24544 19329
rect 26332 19320 26384 19372
rect 1584 19295 1636 19304
rect 1584 19261 1593 19295
rect 1593 19261 1627 19295
rect 1627 19261 1636 19295
rect 1584 19252 1636 19261
rect 1860 19295 1912 19304
rect 1860 19261 1869 19295
rect 1869 19261 1903 19295
rect 1903 19261 1912 19295
rect 1860 19252 1912 19261
rect 24032 19252 24084 19304
rect 16488 19116 16540 19168
rect 19340 19184 19392 19236
rect 17316 19159 17368 19168
rect 17316 19125 17325 19159
rect 17325 19125 17359 19159
rect 17359 19125 17368 19159
rect 17316 19116 17368 19125
rect 17868 19159 17920 19168
rect 17868 19125 17877 19159
rect 17877 19125 17911 19159
rect 17911 19125 17920 19159
rect 17868 19116 17920 19125
rect 20996 19116 21048 19168
rect 27436 19159 27488 19168
rect 27436 19125 27445 19159
rect 27445 19125 27479 19159
rect 27479 19125 27488 19159
rect 27436 19116 27488 19125
rect 28172 19116 28224 19168
rect 5582 19014 5634 19066
rect 5646 19014 5698 19066
rect 5710 19014 5762 19066
rect 5774 19014 5826 19066
rect 5838 19014 5890 19066
rect 14846 19014 14898 19066
rect 14910 19014 14962 19066
rect 14974 19014 15026 19066
rect 15038 19014 15090 19066
rect 15102 19014 15154 19066
rect 24110 19014 24162 19066
rect 24174 19014 24226 19066
rect 24238 19014 24290 19066
rect 24302 19014 24354 19066
rect 24366 19014 24418 19066
rect 1584 18912 1636 18964
rect 17500 18955 17552 18964
rect 17500 18921 17509 18955
rect 17509 18921 17543 18955
rect 17543 18921 17552 18955
rect 17500 18912 17552 18921
rect 21824 18912 21876 18964
rect 24860 18844 24912 18896
rect 17316 18776 17368 18828
rect 17776 18776 17828 18828
rect 27344 18819 27396 18828
rect 27344 18785 27353 18819
rect 27353 18785 27387 18819
rect 27387 18785 27396 18819
rect 27344 18776 27396 18785
rect 27436 18776 27488 18828
rect 2228 18708 2280 18760
rect 2412 18751 2464 18760
rect 2412 18717 2421 18751
rect 2421 18717 2455 18751
rect 2455 18717 2464 18751
rect 2412 18708 2464 18717
rect 16488 18751 16540 18760
rect 16488 18717 16497 18751
rect 16497 18717 16531 18751
rect 16531 18717 16540 18751
rect 16488 18708 16540 18717
rect 16304 18683 16356 18692
rect 16304 18649 16313 18683
rect 16313 18649 16347 18683
rect 16347 18649 16356 18683
rect 16304 18640 16356 18649
rect 12716 18572 12768 18624
rect 21272 18708 21324 18760
rect 21916 18751 21968 18760
rect 21916 18717 21925 18751
rect 21925 18717 21959 18751
rect 21959 18717 21968 18751
rect 21916 18708 21968 18717
rect 22008 18708 22060 18760
rect 27804 18640 27856 18692
rect 18328 18615 18380 18624
rect 18328 18581 18337 18615
rect 18337 18581 18371 18615
rect 18371 18581 18380 18615
rect 18328 18572 18380 18581
rect 22376 18615 22428 18624
rect 22376 18581 22385 18615
rect 22385 18581 22419 18615
rect 22419 18581 22428 18615
rect 22376 18572 22428 18581
rect 10214 18470 10266 18522
rect 10278 18470 10330 18522
rect 10342 18470 10394 18522
rect 10406 18470 10458 18522
rect 10470 18470 10522 18522
rect 19478 18470 19530 18522
rect 19542 18470 19594 18522
rect 19606 18470 19658 18522
rect 19670 18470 19722 18522
rect 19734 18470 19786 18522
rect 16304 18368 16356 18420
rect 20812 18368 20864 18420
rect 21916 18368 21968 18420
rect 25228 18368 25280 18420
rect 27804 18411 27856 18420
rect 27804 18377 27813 18411
rect 27813 18377 27847 18411
rect 27847 18377 27856 18411
rect 27804 18368 27856 18377
rect 18328 18343 18380 18352
rect 18328 18309 18362 18343
rect 18362 18309 18380 18343
rect 18328 18300 18380 18309
rect 12348 18275 12400 18284
rect 12348 18241 12357 18275
rect 12357 18241 12391 18275
rect 12391 18241 12400 18275
rect 12348 18232 12400 18241
rect 12440 18275 12492 18284
rect 12440 18241 12449 18275
rect 12449 18241 12483 18275
rect 12483 18241 12492 18275
rect 12440 18232 12492 18241
rect 13360 18232 13412 18284
rect 14372 18275 14424 18284
rect 14372 18241 14381 18275
rect 14381 18241 14415 18275
rect 14415 18241 14424 18275
rect 14372 18232 14424 18241
rect 14556 18232 14608 18284
rect 14832 18275 14884 18284
rect 14832 18241 14841 18275
rect 14841 18241 14875 18275
rect 14875 18241 14884 18275
rect 14832 18232 14884 18241
rect 14740 18164 14792 18216
rect 16948 18275 17000 18284
rect 16948 18241 16957 18275
rect 16957 18241 16991 18275
rect 16991 18241 17000 18275
rect 16948 18232 17000 18241
rect 17868 18232 17920 18284
rect 22100 18300 22152 18352
rect 22836 18343 22888 18352
rect 21180 18232 21232 18284
rect 22008 18275 22060 18284
rect 22008 18241 22017 18275
rect 22017 18241 22051 18275
rect 22051 18241 22060 18275
rect 22008 18232 22060 18241
rect 22836 18309 22845 18343
rect 22845 18309 22879 18343
rect 22879 18309 22888 18343
rect 22836 18300 22888 18309
rect 22744 18275 22796 18284
rect 22744 18241 22753 18275
rect 22753 18241 22787 18275
rect 22787 18241 22796 18275
rect 22744 18232 22796 18241
rect 23848 18275 23900 18284
rect 23848 18241 23857 18275
rect 23857 18241 23891 18275
rect 23891 18241 23900 18275
rect 23848 18232 23900 18241
rect 25596 18232 25648 18284
rect 27252 18232 27304 18284
rect 27620 18232 27672 18284
rect 28448 18232 28500 18284
rect 28724 18232 28776 18284
rect 17408 18164 17460 18216
rect 21088 18207 21140 18216
rect 21088 18173 21097 18207
rect 21097 18173 21131 18207
rect 21131 18173 21140 18207
rect 21088 18164 21140 18173
rect 22100 18164 22152 18216
rect 23204 18207 23256 18216
rect 23204 18173 23213 18207
rect 23213 18173 23247 18207
rect 23247 18173 23256 18207
rect 23204 18164 23256 18173
rect 23480 18164 23532 18216
rect 24032 18207 24084 18216
rect 24032 18173 24041 18207
rect 24041 18173 24075 18207
rect 24075 18173 24084 18207
rect 24032 18164 24084 18173
rect 24952 18164 25004 18216
rect 14556 18139 14608 18148
rect 14556 18105 14565 18139
rect 14565 18105 14599 18139
rect 14599 18105 14608 18139
rect 14556 18096 14608 18105
rect 1400 18071 1452 18080
rect 1400 18037 1409 18071
rect 1409 18037 1443 18071
rect 1443 18037 1452 18071
rect 1400 18028 1452 18037
rect 11244 18028 11296 18080
rect 13268 18028 13320 18080
rect 14096 18028 14148 18080
rect 18328 18028 18380 18080
rect 19340 18028 19392 18080
rect 20628 18071 20680 18080
rect 20628 18037 20637 18071
rect 20637 18037 20671 18071
rect 20671 18037 20680 18071
rect 20628 18028 20680 18037
rect 21272 18028 21324 18080
rect 23572 18028 23624 18080
rect 25504 18028 25556 18080
rect 26516 18028 26568 18080
rect 5582 17926 5634 17978
rect 5646 17926 5698 17978
rect 5710 17926 5762 17978
rect 5774 17926 5826 17978
rect 5838 17926 5890 17978
rect 14846 17926 14898 17978
rect 14910 17926 14962 17978
rect 14974 17926 15026 17978
rect 15038 17926 15090 17978
rect 15102 17926 15154 17978
rect 24110 17926 24162 17978
rect 24174 17926 24226 17978
rect 24238 17926 24290 17978
rect 24302 17926 24354 17978
rect 24366 17926 24418 17978
rect 16672 17824 16724 17876
rect 18788 17824 18840 17876
rect 23204 17824 23256 17876
rect 16304 17756 16356 17808
rect 26056 17756 26108 17808
rect 1400 17731 1452 17740
rect 1400 17697 1409 17731
rect 1409 17697 1443 17731
rect 1443 17697 1452 17731
rect 1400 17688 1452 17697
rect 2780 17731 2832 17740
rect 2780 17697 2789 17731
rect 2789 17697 2823 17731
rect 2823 17697 2832 17731
rect 2780 17688 2832 17697
rect 14740 17688 14792 17740
rect 26516 17731 26568 17740
rect 11244 17663 11296 17672
rect 11244 17629 11253 17663
rect 11253 17629 11287 17663
rect 11287 17629 11296 17663
rect 11244 17620 11296 17629
rect 11888 17663 11940 17672
rect 11888 17629 11897 17663
rect 11897 17629 11931 17663
rect 11931 17629 11940 17663
rect 11888 17620 11940 17629
rect 14188 17620 14240 17672
rect 14372 17663 14424 17672
rect 14372 17629 14381 17663
rect 14381 17629 14415 17663
rect 14415 17629 14424 17663
rect 14372 17620 14424 17629
rect 18328 17663 18380 17672
rect 1676 17552 1728 17604
rect 13912 17552 13964 17604
rect 18328 17629 18337 17663
rect 18337 17629 18371 17663
rect 18371 17629 18380 17663
rect 18328 17620 18380 17629
rect 20996 17620 21048 17672
rect 26516 17697 26525 17731
rect 26525 17697 26559 17731
rect 26559 17697 26568 17731
rect 26516 17688 26568 17697
rect 26332 17663 26384 17672
rect 26332 17629 26341 17663
rect 26341 17629 26375 17663
rect 26375 17629 26384 17663
rect 26332 17620 26384 17629
rect 13268 17527 13320 17536
rect 13268 17493 13277 17527
rect 13277 17493 13311 17527
rect 13311 17493 13320 17527
rect 13268 17484 13320 17493
rect 14280 17484 14332 17536
rect 14648 17484 14700 17536
rect 19892 17552 19944 17604
rect 20628 17552 20680 17604
rect 22376 17552 22428 17604
rect 23756 17552 23808 17604
rect 24860 17552 24912 17604
rect 27528 17552 27580 17604
rect 16120 17527 16172 17536
rect 16120 17493 16129 17527
rect 16129 17493 16163 17527
rect 16163 17493 16172 17527
rect 16120 17484 16172 17493
rect 17316 17484 17368 17536
rect 18052 17484 18104 17536
rect 21364 17484 21416 17536
rect 25596 17484 25648 17536
rect 10214 17382 10266 17434
rect 10278 17382 10330 17434
rect 10342 17382 10394 17434
rect 10406 17382 10458 17434
rect 10470 17382 10522 17434
rect 19478 17382 19530 17434
rect 19542 17382 19594 17434
rect 19606 17382 19658 17434
rect 19670 17382 19722 17434
rect 19734 17382 19786 17434
rect 1676 17323 1728 17332
rect 1676 17289 1685 17323
rect 1685 17289 1719 17323
rect 1719 17289 1728 17323
rect 1676 17280 1728 17289
rect 12348 17280 12400 17332
rect 13268 17280 13320 17332
rect 13912 17323 13964 17332
rect 13912 17289 13921 17323
rect 13921 17289 13955 17323
rect 13955 17289 13964 17323
rect 13912 17280 13964 17289
rect 14556 17280 14608 17332
rect 14740 17280 14792 17332
rect 21088 17280 21140 17332
rect 22192 17280 22244 17332
rect 22836 17280 22888 17332
rect 23848 17280 23900 17332
rect 26332 17280 26384 17332
rect 13360 17212 13412 17264
rect 14096 17212 14148 17264
rect 1768 17187 1820 17196
rect 1768 17153 1777 17187
rect 1777 17153 1811 17187
rect 1811 17153 1820 17187
rect 1768 17144 1820 17153
rect 14648 17144 14700 17196
rect 6552 17076 6604 17128
rect 12900 17119 12952 17128
rect 12900 17085 12909 17119
rect 12909 17085 12943 17119
rect 12943 17085 12952 17119
rect 12900 17076 12952 17085
rect 14464 17076 14516 17128
rect 15568 17144 15620 17196
rect 16856 17187 16908 17196
rect 16856 17153 16865 17187
rect 16865 17153 16899 17187
rect 16899 17153 16908 17187
rect 16856 17144 16908 17153
rect 20168 17187 20220 17196
rect 20168 17153 20177 17187
rect 20177 17153 20211 17187
rect 20211 17153 20220 17187
rect 20168 17144 20220 17153
rect 20628 17144 20680 17196
rect 22744 17212 22796 17264
rect 23204 17212 23256 17264
rect 27160 17212 27212 17264
rect 15476 17076 15528 17128
rect 18144 17076 18196 17128
rect 21364 17076 21416 17128
rect 22100 17187 22152 17196
rect 22100 17153 22109 17187
rect 22109 17153 22143 17187
rect 22143 17153 22152 17187
rect 22100 17144 22152 17153
rect 25596 17144 25648 17196
rect 22192 17076 22244 17128
rect 22836 17076 22888 17128
rect 23664 17076 23716 17128
rect 13268 17008 13320 17060
rect 14004 17008 14056 17060
rect 15568 17051 15620 17060
rect 15568 17017 15577 17051
rect 15577 17017 15611 17051
rect 15611 17017 15620 17051
rect 15568 17008 15620 17017
rect 17960 16940 18012 16992
rect 20260 16983 20312 16992
rect 20260 16949 20269 16983
rect 20269 16949 20303 16983
rect 20303 16949 20312 16983
rect 20260 16940 20312 16949
rect 25872 17144 25924 17196
rect 26240 17144 26292 17196
rect 27068 17187 27120 17196
rect 27068 17153 27077 17187
rect 27077 17153 27111 17187
rect 27111 17153 27120 17187
rect 27436 17212 27488 17264
rect 27068 17144 27120 17153
rect 26332 17076 26384 17128
rect 27620 17144 27672 17196
rect 27344 17008 27396 17060
rect 26332 16940 26384 16992
rect 27988 16940 28040 16992
rect 5582 16838 5634 16890
rect 5646 16838 5698 16890
rect 5710 16838 5762 16890
rect 5774 16838 5826 16890
rect 5838 16838 5890 16890
rect 14846 16838 14898 16890
rect 14910 16838 14962 16890
rect 14974 16838 15026 16890
rect 15038 16838 15090 16890
rect 15102 16838 15154 16890
rect 24110 16838 24162 16890
rect 24174 16838 24226 16890
rect 24238 16838 24290 16890
rect 24302 16838 24354 16890
rect 24366 16838 24418 16890
rect 14188 16736 14240 16788
rect 14188 16643 14240 16652
rect 14188 16609 14197 16643
rect 14197 16609 14231 16643
rect 14231 16609 14240 16643
rect 14188 16600 14240 16609
rect 14280 16600 14332 16652
rect 14096 16575 14148 16584
rect 14096 16541 14105 16575
rect 14105 16541 14139 16575
rect 14139 16541 14148 16575
rect 14096 16532 14148 16541
rect 14556 16736 14608 16788
rect 16120 16736 16172 16788
rect 17408 16736 17460 16788
rect 18144 16736 18196 16788
rect 23756 16779 23808 16788
rect 23756 16745 23765 16779
rect 23765 16745 23799 16779
rect 23799 16745 23808 16779
rect 23756 16736 23808 16745
rect 21180 16668 21232 16720
rect 15476 16643 15528 16652
rect 15476 16609 15485 16643
rect 15485 16609 15519 16643
rect 15519 16609 15528 16643
rect 15476 16600 15528 16609
rect 17592 16643 17644 16652
rect 17592 16609 17601 16643
rect 17601 16609 17635 16643
rect 17635 16609 17644 16643
rect 17592 16600 17644 16609
rect 17868 16600 17920 16652
rect 15384 16575 15436 16584
rect 15384 16541 15393 16575
rect 15393 16541 15427 16575
rect 15427 16541 15436 16575
rect 15384 16532 15436 16541
rect 17316 16575 17368 16584
rect 19340 16600 19392 16652
rect 19984 16600 20036 16652
rect 20812 16600 20864 16652
rect 26976 16736 27028 16788
rect 26332 16668 26384 16720
rect 27988 16643 28040 16652
rect 17316 16541 17334 16575
rect 17334 16541 17368 16575
rect 17316 16532 17368 16541
rect 20260 16532 20312 16584
rect 23572 16575 23624 16584
rect 23572 16541 23581 16575
rect 23581 16541 23615 16575
rect 23615 16541 23624 16575
rect 23572 16532 23624 16541
rect 27988 16609 27997 16643
rect 27997 16609 28031 16643
rect 28031 16609 28040 16643
rect 27988 16600 28040 16609
rect 28172 16643 28224 16652
rect 28172 16609 28181 16643
rect 28181 16609 28215 16643
rect 28215 16609 28224 16643
rect 28172 16600 28224 16609
rect 25504 16575 25556 16584
rect 25504 16541 25513 16575
rect 25513 16541 25547 16575
rect 25547 16541 25556 16575
rect 25504 16532 25556 16541
rect 25688 16575 25740 16584
rect 25688 16541 25697 16575
rect 25697 16541 25731 16575
rect 25731 16541 25740 16575
rect 25688 16532 25740 16541
rect 25780 16532 25832 16584
rect 15660 16464 15712 16516
rect 16212 16439 16264 16448
rect 16212 16405 16221 16439
rect 16221 16405 16255 16439
rect 16255 16405 16264 16439
rect 19340 16439 19392 16448
rect 16212 16396 16264 16405
rect 19340 16405 19349 16439
rect 19349 16405 19383 16439
rect 19383 16405 19392 16439
rect 19340 16396 19392 16405
rect 27068 16396 27120 16448
rect 10214 16294 10266 16346
rect 10278 16294 10330 16346
rect 10342 16294 10394 16346
rect 10406 16294 10458 16346
rect 10470 16294 10522 16346
rect 19478 16294 19530 16346
rect 19542 16294 19594 16346
rect 19606 16294 19658 16346
rect 19670 16294 19722 16346
rect 19734 16294 19786 16346
rect 7288 16192 7340 16244
rect 15660 16235 15712 16244
rect 15660 16201 15669 16235
rect 15669 16201 15703 16235
rect 15703 16201 15712 16235
rect 15660 16192 15712 16201
rect 18052 16235 18104 16244
rect 18052 16201 18061 16235
rect 18061 16201 18095 16235
rect 18095 16201 18104 16235
rect 18052 16192 18104 16201
rect 19892 16192 19944 16244
rect 19248 16124 19300 16176
rect 27344 16192 27396 16244
rect 13360 16056 13412 16108
rect 16028 16056 16080 16108
rect 16212 16056 16264 16108
rect 12900 15988 12952 16040
rect 14556 15988 14608 16040
rect 18696 16031 18748 16040
rect 16488 15920 16540 15972
rect 18696 15997 18705 16031
rect 18705 15997 18739 16031
rect 18739 15997 18748 16031
rect 18696 15988 18748 15997
rect 20720 16056 20772 16108
rect 25872 16124 25924 16176
rect 25780 16099 25832 16108
rect 25780 16065 25789 16099
rect 25789 16065 25823 16099
rect 25823 16065 25832 16099
rect 28080 16167 28132 16176
rect 28080 16133 28089 16167
rect 28089 16133 28123 16167
rect 28123 16133 28132 16167
rect 28080 16124 28132 16133
rect 25780 16056 25832 16065
rect 26240 16056 26292 16108
rect 19892 15988 19944 16040
rect 25872 15988 25924 16040
rect 26976 16031 27028 16040
rect 26976 15997 26985 16031
rect 26985 15997 27019 16031
rect 27019 15997 27028 16031
rect 26976 15988 27028 15997
rect 26056 15920 26108 15972
rect 4344 15852 4396 15904
rect 12164 15852 12216 15904
rect 17684 15852 17736 15904
rect 26148 15852 26200 15904
rect 26608 15852 26660 15904
rect 27988 15895 28040 15904
rect 27988 15861 27997 15895
rect 27997 15861 28031 15895
rect 28031 15861 28040 15895
rect 27988 15852 28040 15861
rect 5582 15750 5634 15802
rect 5646 15750 5698 15802
rect 5710 15750 5762 15802
rect 5774 15750 5826 15802
rect 5838 15750 5890 15802
rect 14846 15750 14898 15802
rect 14910 15750 14962 15802
rect 14974 15750 15026 15802
rect 15038 15750 15090 15802
rect 15102 15750 15154 15802
rect 24110 15750 24162 15802
rect 24174 15750 24226 15802
rect 24238 15750 24290 15802
rect 24302 15750 24354 15802
rect 24366 15750 24418 15802
rect 14096 15648 14148 15700
rect 18696 15648 18748 15700
rect 19248 15691 19300 15700
rect 19248 15657 19257 15691
rect 19257 15657 19291 15691
rect 19291 15657 19300 15691
rect 19248 15648 19300 15657
rect 13360 15580 13412 15632
rect 14188 15623 14240 15632
rect 14188 15589 14197 15623
rect 14197 15589 14231 15623
rect 14231 15589 14240 15623
rect 14188 15580 14240 15589
rect 15016 15580 15068 15632
rect 17684 15580 17736 15632
rect 12440 15512 12492 15564
rect 14372 15512 14424 15564
rect 16212 15512 16264 15564
rect 19156 15580 19208 15632
rect 20720 15691 20772 15700
rect 20720 15657 20729 15691
rect 20729 15657 20763 15691
rect 20763 15657 20772 15691
rect 20720 15648 20772 15657
rect 24584 15648 24636 15700
rect 20628 15580 20680 15632
rect 27988 15648 28040 15700
rect 1400 15444 1452 15496
rect 3976 15487 4028 15496
rect 3976 15453 3985 15487
rect 3985 15453 4019 15487
rect 4019 15453 4028 15487
rect 3976 15444 4028 15453
rect 12164 15487 12216 15496
rect 12164 15453 12173 15487
rect 12173 15453 12207 15487
rect 12207 15453 12216 15487
rect 12164 15444 12216 15453
rect 15384 15444 15436 15496
rect 15752 15444 15804 15496
rect 18328 15487 18380 15496
rect 18328 15453 18337 15487
rect 18337 15453 18371 15487
rect 18371 15453 18380 15487
rect 18328 15444 18380 15453
rect 18420 15487 18472 15496
rect 18420 15453 18429 15487
rect 18429 15453 18463 15487
rect 18463 15453 18472 15487
rect 18420 15444 18472 15453
rect 14556 15419 14608 15428
rect 14556 15385 14565 15419
rect 14565 15385 14599 15419
rect 14599 15385 14608 15419
rect 14556 15376 14608 15385
rect 16304 15376 16356 15428
rect 19432 15487 19484 15496
rect 19432 15453 19441 15487
rect 19441 15453 19475 15487
rect 19475 15453 19484 15487
rect 19432 15444 19484 15453
rect 19524 15487 19576 15496
rect 19524 15453 19533 15487
rect 19533 15453 19567 15487
rect 19567 15453 19576 15487
rect 22836 15555 22888 15564
rect 19524 15444 19576 15453
rect 4160 15308 4212 15360
rect 12808 15351 12860 15360
rect 12808 15317 12817 15351
rect 12817 15317 12851 15351
rect 12851 15317 12860 15351
rect 12808 15308 12860 15317
rect 15476 15308 15528 15360
rect 18696 15308 18748 15360
rect 19156 15308 19208 15360
rect 22836 15521 22845 15555
rect 22845 15521 22879 15555
rect 22879 15521 22888 15555
rect 22836 15512 22888 15521
rect 25688 15512 25740 15564
rect 26056 15512 26108 15564
rect 28172 15555 28224 15564
rect 28172 15521 28181 15555
rect 28181 15521 28215 15555
rect 28215 15521 28224 15555
rect 28172 15512 28224 15521
rect 23572 15444 23624 15496
rect 24860 15444 24912 15496
rect 24124 15376 24176 15428
rect 25320 15376 25372 15428
rect 23020 15308 23072 15360
rect 23664 15308 23716 15360
rect 25872 15308 25924 15360
rect 26332 15376 26384 15428
rect 26516 15419 26568 15428
rect 26516 15385 26525 15419
rect 26525 15385 26559 15419
rect 26559 15385 26568 15419
rect 26516 15376 26568 15385
rect 26424 15308 26476 15360
rect 10214 15206 10266 15258
rect 10278 15206 10330 15258
rect 10342 15206 10394 15258
rect 10406 15206 10458 15258
rect 10470 15206 10522 15258
rect 19478 15206 19530 15258
rect 19542 15206 19594 15258
rect 19606 15206 19658 15258
rect 19670 15206 19722 15258
rect 19734 15206 19786 15258
rect 4068 15104 4120 15156
rect 13360 15147 13412 15156
rect 13360 15113 13369 15147
rect 13369 15113 13403 15147
rect 13403 15113 13412 15147
rect 13360 15104 13412 15113
rect 18328 15104 18380 15156
rect 23664 15104 23716 15156
rect 24124 15147 24176 15156
rect 24124 15113 24133 15147
rect 24133 15113 24167 15147
rect 24167 15113 24176 15147
rect 24124 15104 24176 15113
rect 24768 15104 24820 15156
rect 26240 15104 26292 15156
rect 26516 15104 26568 15156
rect 4160 15079 4212 15088
rect 4160 15045 4169 15079
rect 4169 15045 4203 15079
rect 4203 15045 4212 15079
rect 4160 15036 4212 15045
rect 12808 15036 12860 15088
rect 19984 15036 20036 15088
rect 22284 15036 22336 15088
rect 25320 15036 25372 15088
rect 25596 15036 25648 15088
rect 2136 14968 2188 15020
rect 4344 15011 4396 15020
rect 4344 14977 4353 15011
rect 4353 14977 4387 15011
rect 4387 14977 4396 15011
rect 4344 14968 4396 14977
rect 11888 14968 11940 15020
rect 15016 15011 15068 15020
rect 15016 14977 15025 15011
rect 15025 14977 15059 15011
rect 15059 14977 15068 15011
rect 15016 14968 15068 14977
rect 15292 14968 15344 15020
rect 20536 15011 20588 15020
rect 20536 14977 20545 15011
rect 20545 14977 20579 15011
rect 20579 14977 20588 15011
rect 20536 14968 20588 14977
rect 22100 15011 22152 15020
rect 22100 14977 22109 15011
rect 22109 14977 22143 15011
rect 22143 14977 22152 15011
rect 22100 14968 22152 14977
rect 26424 15011 26476 15020
rect 2780 14943 2832 14952
rect 2780 14909 2789 14943
rect 2789 14909 2823 14943
rect 2823 14909 2832 14943
rect 2780 14900 2832 14909
rect 16488 14900 16540 14952
rect 20260 14900 20312 14952
rect 21824 14900 21876 14952
rect 25136 14900 25188 14952
rect 25780 14900 25832 14952
rect 26424 14977 26433 15011
rect 26433 14977 26467 15011
rect 26467 14977 26476 15011
rect 26424 14968 26476 14977
rect 20536 14832 20588 14884
rect 22284 14875 22336 14884
rect 22284 14841 22293 14875
rect 22293 14841 22327 14875
rect 22327 14841 22336 14875
rect 22284 14832 22336 14841
rect 26332 14900 26384 14952
rect 27252 14943 27304 14952
rect 27252 14909 27261 14943
rect 27261 14909 27295 14943
rect 27295 14909 27304 14943
rect 27252 14900 27304 14909
rect 27436 14943 27488 14952
rect 27436 14909 27445 14943
rect 27445 14909 27479 14943
rect 27479 14909 27488 14943
rect 27436 14900 27488 14909
rect 26884 14832 26936 14884
rect 27528 14832 27580 14884
rect 1584 14764 1636 14816
rect 15200 14764 15252 14816
rect 19340 14764 19392 14816
rect 19984 14764 20036 14816
rect 24860 14764 24912 14816
rect 25228 14764 25280 14816
rect 26516 14764 26568 14816
rect 27344 14764 27396 14816
rect 5582 14662 5634 14714
rect 5646 14662 5698 14714
rect 5710 14662 5762 14714
rect 5774 14662 5826 14714
rect 5838 14662 5890 14714
rect 14846 14662 14898 14714
rect 14910 14662 14962 14714
rect 14974 14662 15026 14714
rect 15038 14662 15090 14714
rect 15102 14662 15154 14714
rect 24110 14662 24162 14714
rect 24174 14662 24226 14714
rect 24238 14662 24290 14714
rect 24302 14662 24354 14714
rect 24366 14662 24418 14714
rect 15476 14560 15528 14612
rect 16856 14560 16908 14612
rect 22100 14560 22152 14612
rect 25136 14603 25188 14612
rect 25136 14569 25145 14603
rect 25145 14569 25179 14603
rect 25179 14569 25188 14603
rect 25136 14560 25188 14569
rect 27436 14560 27488 14612
rect 22744 14492 22796 14544
rect 24952 14492 25004 14544
rect 1400 14467 1452 14476
rect 1400 14433 1409 14467
rect 1409 14433 1443 14467
rect 1443 14433 1452 14467
rect 1400 14424 1452 14433
rect 1584 14467 1636 14476
rect 1584 14433 1593 14467
rect 1593 14433 1627 14467
rect 1627 14433 1636 14467
rect 1584 14424 1636 14433
rect 1860 14467 1912 14476
rect 1860 14433 1869 14467
rect 1869 14433 1903 14467
rect 1903 14433 1912 14467
rect 1860 14424 1912 14433
rect 19340 14424 19392 14476
rect 20812 14424 20864 14476
rect 24492 14467 24544 14476
rect 24492 14433 24501 14467
rect 24501 14433 24535 14467
rect 24535 14433 24544 14467
rect 24492 14424 24544 14433
rect 24676 14467 24728 14476
rect 24676 14433 24685 14467
rect 24685 14433 24719 14467
rect 24719 14433 24728 14467
rect 24676 14424 24728 14433
rect 27528 14467 27580 14476
rect 27528 14433 27537 14467
rect 27537 14433 27571 14467
rect 27571 14433 27580 14467
rect 27528 14424 27580 14433
rect 15568 14356 15620 14408
rect 16120 14356 16172 14408
rect 19984 14399 20036 14408
rect 19984 14365 19993 14399
rect 19993 14365 20027 14399
rect 20027 14365 20036 14399
rect 19984 14356 20036 14365
rect 20996 14399 21048 14408
rect 20996 14365 21005 14399
rect 21005 14365 21039 14399
rect 21039 14365 21048 14399
rect 20996 14356 21048 14365
rect 21824 14356 21876 14408
rect 23020 14399 23072 14408
rect 23020 14365 23029 14399
rect 23029 14365 23063 14399
rect 23063 14365 23072 14399
rect 23020 14356 23072 14365
rect 23388 14356 23440 14408
rect 24768 14399 24820 14408
rect 24768 14365 24777 14399
rect 24777 14365 24811 14399
rect 24811 14365 24820 14399
rect 24768 14356 24820 14365
rect 25596 14399 25648 14408
rect 25596 14365 25605 14399
rect 25605 14365 25639 14399
rect 25639 14365 25648 14399
rect 25596 14356 25648 14365
rect 25872 14399 25924 14408
rect 25872 14365 25881 14399
rect 25881 14365 25915 14399
rect 25915 14365 25924 14399
rect 25872 14356 25924 14365
rect 28172 14399 28224 14408
rect 28172 14365 28181 14399
rect 28181 14365 28215 14399
rect 28215 14365 28224 14399
rect 28172 14356 28224 14365
rect 15200 14288 15252 14340
rect 15384 14288 15436 14340
rect 16672 14288 16724 14340
rect 21272 14331 21324 14340
rect 21272 14297 21306 14331
rect 21306 14297 21324 14331
rect 21272 14288 21324 14297
rect 27896 14288 27948 14340
rect 14280 14220 14332 14272
rect 20076 14220 20128 14272
rect 25780 14220 25832 14272
rect 26608 14220 26660 14272
rect 10214 14118 10266 14170
rect 10278 14118 10330 14170
rect 10342 14118 10394 14170
rect 10406 14118 10458 14170
rect 10470 14118 10522 14170
rect 19478 14118 19530 14170
rect 19542 14118 19594 14170
rect 19606 14118 19658 14170
rect 19670 14118 19722 14170
rect 19734 14118 19786 14170
rect 16672 14016 16724 14068
rect 11888 13880 11940 13932
rect 14740 13948 14792 14000
rect 16856 13948 16908 14000
rect 17868 14016 17920 14068
rect 18696 14059 18748 14068
rect 18696 14025 18705 14059
rect 18705 14025 18739 14059
rect 18739 14025 18748 14059
rect 18696 14016 18748 14025
rect 20536 14016 20588 14068
rect 25136 14016 25188 14068
rect 25596 14016 25648 14068
rect 27896 14059 27948 14068
rect 27896 14025 27905 14059
rect 27905 14025 27939 14059
rect 27939 14025 27948 14059
rect 27896 14016 27948 14025
rect 14096 13880 14148 13932
rect 15476 13880 15528 13932
rect 17776 13880 17828 13932
rect 18328 13880 18380 13932
rect 20996 13948 21048 14000
rect 25872 13948 25924 14000
rect 27252 13948 27304 14000
rect 19800 13923 19852 13932
rect 19800 13889 19834 13923
rect 19834 13889 19852 13923
rect 23296 13923 23348 13932
rect 19800 13880 19852 13889
rect 23296 13889 23305 13923
rect 23305 13889 23339 13923
rect 23339 13889 23348 13923
rect 23296 13880 23348 13889
rect 23388 13923 23440 13932
rect 23388 13889 23397 13923
rect 23397 13889 23431 13923
rect 23431 13889 23440 13923
rect 23388 13880 23440 13889
rect 1492 13855 1544 13864
rect 1492 13821 1501 13855
rect 1501 13821 1535 13855
rect 1535 13821 1544 13855
rect 1492 13812 1544 13821
rect 1676 13855 1728 13864
rect 1676 13821 1685 13855
rect 1685 13821 1719 13855
rect 1719 13821 1728 13855
rect 1676 13812 1728 13821
rect 1952 13855 2004 13864
rect 1952 13821 1961 13855
rect 1961 13821 1995 13855
rect 1995 13821 2004 13855
rect 1952 13812 2004 13821
rect 14556 13812 14608 13864
rect 23020 13812 23072 13864
rect 25412 13880 25464 13932
rect 27804 13923 27856 13932
rect 25504 13812 25556 13864
rect 27804 13889 27813 13923
rect 27813 13889 27847 13923
rect 27847 13889 27856 13923
rect 27804 13880 27856 13889
rect 25688 13744 25740 13796
rect 27252 13812 27304 13864
rect 15568 13676 15620 13728
rect 17132 13676 17184 13728
rect 17408 13719 17460 13728
rect 17408 13685 17417 13719
rect 17417 13685 17451 13719
rect 17451 13685 17460 13719
rect 17408 13676 17460 13685
rect 25964 13719 26016 13728
rect 25964 13685 25973 13719
rect 25973 13685 26007 13719
rect 26007 13685 26016 13719
rect 25964 13676 26016 13685
rect 5582 13574 5634 13626
rect 5646 13574 5698 13626
rect 5710 13574 5762 13626
rect 5774 13574 5826 13626
rect 5838 13574 5890 13626
rect 14846 13574 14898 13626
rect 14910 13574 14962 13626
rect 14974 13574 15026 13626
rect 15038 13574 15090 13626
rect 15102 13574 15154 13626
rect 24110 13574 24162 13626
rect 24174 13574 24226 13626
rect 24238 13574 24290 13626
rect 24302 13574 24354 13626
rect 24366 13574 24418 13626
rect 1676 13472 1728 13524
rect 14096 13515 14148 13524
rect 14096 13481 14105 13515
rect 14105 13481 14139 13515
rect 14139 13481 14148 13515
rect 14096 13472 14148 13481
rect 19800 13472 19852 13524
rect 25688 13515 25740 13524
rect 21180 13404 21232 13456
rect 21364 13336 21416 13388
rect 2136 13268 2188 13320
rect 2780 13268 2832 13320
rect 14280 13311 14332 13320
rect 14280 13277 14289 13311
rect 14289 13277 14323 13311
rect 14323 13277 14332 13311
rect 14280 13268 14332 13277
rect 15476 13268 15528 13320
rect 16856 13268 16908 13320
rect 17592 13268 17644 13320
rect 20076 13311 20128 13320
rect 20076 13277 20085 13311
rect 20085 13277 20119 13311
rect 20119 13277 20128 13311
rect 20076 13268 20128 13277
rect 15384 13243 15436 13252
rect 15384 13209 15393 13243
rect 15393 13209 15427 13243
rect 15427 13209 15436 13243
rect 15384 13200 15436 13209
rect 17224 13243 17276 13252
rect 17224 13209 17258 13243
rect 17258 13209 17276 13243
rect 17224 13200 17276 13209
rect 17316 13200 17368 13252
rect 22008 13268 22060 13320
rect 23388 13268 23440 13320
rect 24676 13268 24728 13320
rect 25688 13481 25697 13515
rect 25697 13481 25731 13515
rect 25731 13481 25740 13515
rect 25688 13472 25740 13481
rect 25780 13472 25832 13524
rect 26976 13404 27028 13456
rect 25964 13336 26016 13388
rect 27528 13379 27580 13388
rect 27528 13345 27537 13379
rect 27537 13345 27571 13379
rect 27571 13345 27580 13379
rect 27528 13336 27580 13345
rect 25228 13268 25280 13320
rect 25504 13268 25556 13320
rect 26240 13268 26292 13320
rect 15568 13175 15620 13184
rect 15568 13141 15593 13175
rect 15593 13141 15620 13175
rect 15752 13175 15804 13184
rect 15568 13132 15620 13141
rect 15752 13141 15761 13175
rect 15761 13141 15795 13175
rect 15795 13141 15804 13175
rect 15752 13132 15804 13141
rect 18328 13175 18380 13184
rect 18328 13141 18337 13175
rect 18337 13141 18371 13175
rect 18371 13141 18380 13175
rect 18328 13132 18380 13141
rect 20996 13132 21048 13184
rect 23572 13200 23624 13252
rect 24032 13200 24084 13252
rect 28080 13200 28132 13252
rect 23204 13132 23256 13184
rect 10214 13030 10266 13082
rect 10278 13030 10330 13082
rect 10342 13030 10394 13082
rect 10406 13030 10458 13082
rect 10470 13030 10522 13082
rect 19478 13030 19530 13082
rect 19542 13030 19594 13082
rect 19606 13030 19658 13082
rect 19670 13030 19722 13082
rect 19734 13030 19786 13082
rect 16120 12971 16172 12980
rect 16120 12937 16129 12971
rect 16129 12937 16163 12971
rect 16163 12937 16172 12971
rect 16120 12928 16172 12937
rect 23204 12971 23256 12980
rect 23204 12937 23213 12971
rect 23213 12937 23247 12971
rect 23247 12937 23256 12971
rect 23204 12928 23256 12937
rect 24676 12971 24728 12980
rect 24676 12937 24685 12971
rect 24685 12937 24719 12971
rect 24719 12937 24728 12971
rect 24676 12928 24728 12937
rect 28080 12971 28132 12980
rect 28080 12937 28089 12971
rect 28089 12937 28123 12971
rect 28123 12937 28132 12971
rect 28080 12928 28132 12937
rect 1492 12792 1544 12844
rect 14740 12835 14792 12844
rect 14740 12801 14749 12835
rect 14749 12801 14783 12835
rect 14783 12801 14792 12835
rect 17316 12860 17368 12912
rect 18328 12860 18380 12912
rect 14740 12792 14792 12801
rect 15568 12792 15620 12844
rect 17776 12792 17828 12844
rect 20812 12835 20864 12844
rect 20812 12801 20821 12835
rect 20821 12801 20855 12835
rect 20855 12801 20864 12835
rect 20812 12792 20864 12801
rect 20996 12835 21048 12844
rect 20996 12801 21005 12835
rect 21005 12801 21039 12835
rect 21039 12801 21048 12835
rect 20996 12792 21048 12801
rect 22100 12835 22152 12844
rect 22100 12801 22134 12835
rect 22134 12801 22152 12835
rect 22100 12792 22152 12801
rect 23848 12792 23900 12844
rect 25412 12792 25464 12844
rect 25688 12792 25740 12844
rect 25872 12835 25924 12844
rect 25872 12801 25881 12835
rect 25881 12801 25915 12835
rect 25915 12801 25924 12835
rect 25872 12792 25924 12801
rect 27712 12792 27764 12844
rect 27988 12835 28040 12844
rect 27988 12801 27997 12835
rect 27997 12801 28031 12835
rect 28031 12801 28040 12835
rect 27988 12792 28040 12801
rect 17132 12724 17184 12776
rect 21824 12767 21876 12776
rect 21824 12733 21833 12767
rect 21833 12733 21867 12767
rect 21867 12733 21876 12767
rect 21824 12724 21876 12733
rect 24492 12724 24544 12776
rect 25964 12724 26016 12776
rect 26884 12656 26936 12708
rect 21088 12588 21140 12640
rect 26976 12631 27028 12640
rect 26976 12597 26985 12631
rect 26985 12597 27019 12631
rect 27019 12597 27028 12631
rect 26976 12588 27028 12597
rect 5582 12486 5634 12538
rect 5646 12486 5698 12538
rect 5710 12486 5762 12538
rect 5774 12486 5826 12538
rect 5838 12486 5890 12538
rect 14846 12486 14898 12538
rect 14910 12486 14962 12538
rect 14974 12486 15026 12538
rect 15038 12486 15090 12538
rect 15102 12486 15154 12538
rect 24110 12486 24162 12538
rect 24174 12486 24226 12538
rect 24238 12486 24290 12538
rect 24302 12486 24354 12538
rect 24366 12486 24418 12538
rect 15568 12427 15620 12436
rect 15568 12393 15577 12427
rect 15577 12393 15611 12427
rect 15611 12393 15620 12427
rect 15568 12384 15620 12393
rect 17224 12427 17276 12436
rect 17224 12393 17233 12427
rect 17233 12393 17267 12427
rect 17267 12393 17276 12427
rect 17224 12384 17276 12393
rect 22100 12384 22152 12436
rect 23848 12427 23900 12436
rect 23848 12393 23857 12427
rect 23857 12393 23891 12427
rect 23891 12393 23900 12427
rect 23848 12384 23900 12393
rect 27712 12427 27764 12436
rect 27712 12393 27721 12427
rect 27721 12393 27755 12427
rect 27755 12393 27764 12427
rect 27712 12384 27764 12393
rect 26332 12316 26384 12368
rect 20720 12248 20772 12300
rect 21824 12248 21876 12300
rect 26148 12248 26200 12300
rect 27344 12248 27396 12300
rect 27712 12248 27764 12300
rect 1492 12223 1544 12232
rect 1492 12189 1501 12223
rect 1501 12189 1535 12223
rect 1535 12189 1544 12223
rect 1492 12180 1544 12189
rect 15752 12223 15804 12232
rect 15752 12189 15761 12223
rect 15761 12189 15795 12223
rect 15795 12189 15804 12223
rect 15752 12180 15804 12189
rect 17408 12223 17460 12232
rect 17408 12189 17417 12223
rect 17417 12189 17451 12223
rect 17451 12189 17460 12223
rect 17408 12180 17460 12189
rect 18696 12180 18748 12232
rect 21088 12223 21140 12232
rect 21088 12189 21097 12223
rect 21097 12189 21131 12223
rect 21131 12189 21140 12223
rect 21088 12180 21140 12189
rect 3332 12112 3384 12164
rect 26884 12223 26936 12232
rect 26884 12189 26893 12223
rect 26893 12189 26927 12223
rect 26927 12189 26936 12223
rect 26884 12180 26936 12189
rect 22836 12112 22888 12164
rect 24952 12112 25004 12164
rect 26424 12112 26476 12164
rect 27252 12180 27304 12232
rect 19340 12087 19392 12096
rect 19340 12053 19349 12087
rect 19349 12053 19383 12087
rect 19383 12053 19392 12087
rect 19340 12044 19392 12053
rect 25872 12044 25924 12096
rect 10214 11942 10266 11994
rect 10278 11942 10330 11994
rect 10342 11942 10394 11994
rect 10406 11942 10458 11994
rect 10470 11942 10522 11994
rect 19478 11942 19530 11994
rect 19542 11942 19594 11994
rect 19606 11942 19658 11994
rect 19670 11942 19722 11994
rect 19734 11942 19786 11994
rect 18420 11840 18472 11892
rect 19892 11840 19944 11892
rect 22836 11883 22888 11892
rect 22836 11849 22845 11883
rect 22845 11849 22879 11883
rect 22879 11849 22888 11883
rect 22836 11840 22888 11849
rect 23296 11840 23348 11892
rect 23940 11883 23992 11892
rect 23940 11849 23949 11883
rect 23949 11849 23983 11883
rect 23983 11849 23992 11883
rect 23940 11840 23992 11849
rect 24952 11883 25004 11892
rect 24952 11849 24961 11883
rect 24961 11849 24995 11883
rect 24995 11849 25004 11883
rect 24952 11840 25004 11849
rect 26424 11840 26476 11892
rect 19340 11772 19392 11824
rect 1492 11747 1544 11756
rect 1492 11713 1501 11747
rect 1501 11713 1535 11747
rect 1535 11713 1544 11747
rect 1492 11704 1544 11713
rect 15476 11704 15528 11756
rect 17868 11704 17920 11756
rect 18696 11747 18748 11756
rect 18696 11713 18705 11747
rect 18705 11713 18739 11747
rect 18739 11713 18748 11747
rect 18696 11704 18748 11713
rect 19984 11747 20036 11756
rect 19984 11713 19993 11747
rect 19993 11713 20027 11747
rect 20027 11713 20036 11747
rect 19984 11704 20036 11713
rect 22008 11772 22060 11824
rect 23848 11815 23900 11824
rect 23848 11781 23857 11815
rect 23857 11781 23891 11815
rect 23891 11781 23900 11815
rect 23848 11772 23900 11781
rect 25228 11772 25280 11824
rect 25688 11772 25740 11824
rect 20904 11704 20956 11756
rect 23020 11747 23072 11756
rect 23020 11713 23029 11747
rect 23029 11713 23063 11747
rect 23063 11713 23072 11747
rect 23020 11704 23072 11713
rect 25044 11704 25096 11756
rect 28172 11704 28224 11756
rect 1860 11636 1912 11688
rect 1952 11679 2004 11688
rect 1952 11645 1961 11679
rect 1961 11645 1995 11679
rect 1995 11645 2004 11679
rect 24032 11679 24084 11688
rect 1952 11636 2004 11645
rect 24032 11645 24041 11679
rect 24041 11645 24075 11679
rect 24075 11645 24084 11679
rect 24032 11636 24084 11645
rect 19340 11568 19392 11620
rect 17592 11500 17644 11552
rect 21364 11500 21416 11552
rect 27896 11500 27948 11552
rect 5582 11398 5634 11450
rect 5646 11398 5698 11450
rect 5710 11398 5762 11450
rect 5774 11398 5826 11450
rect 5838 11398 5890 11450
rect 14846 11398 14898 11450
rect 14910 11398 14962 11450
rect 14974 11398 15026 11450
rect 15038 11398 15090 11450
rect 15102 11398 15154 11450
rect 24110 11398 24162 11450
rect 24174 11398 24226 11450
rect 24238 11398 24290 11450
rect 24302 11398 24354 11450
rect 24366 11398 24418 11450
rect 1860 11339 1912 11348
rect 1860 11305 1869 11339
rect 1869 11305 1903 11339
rect 1903 11305 1912 11339
rect 1860 11296 1912 11305
rect 18696 11339 18748 11348
rect 18696 11305 18705 11339
rect 18705 11305 18739 11339
rect 18739 11305 18748 11339
rect 18696 11296 18748 11305
rect 26240 11296 26292 11348
rect 13820 11160 13872 11212
rect 2044 11092 2096 11144
rect 16948 11160 17000 11212
rect 17316 11203 17368 11212
rect 17316 11169 17325 11203
rect 17325 11169 17359 11203
rect 17359 11169 17368 11203
rect 17316 11160 17368 11169
rect 20720 11203 20772 11212
rect 20720 11169 20729 11203
rect 20729 11169 20763 11203
rect 20763 11169 20772 11203
rect 20720 11160 20772 11169
rect 16580 11092 16632 11144
rect 17592 11135 17644 11144
rect 17592 11101 17626 11135
rect 17626 11101 17644 11135
rect 17592 11092 17644 11101
rect 27528 11203 27580 11212
rect 27528 11169 27537 11203
rect 27537 11169 27571 11203
rect 27571 11169 27580 11203
rect 27528 11160 27580 11169
rect 27896 11160 27948 11212
rect 21364 11135 21416 11144
rect 21364 11101 21373 11135
rect 21373 11101 21407 11135
rect 21407 11101 21416 11135
rect 21364 11092 21416 11101
rect 19248 11024 19300 11076
rect 27988 11067 28040 11076
rect 27988 11033 27997 11067
rect 27997 11033 28031 11067
rect 28031 11033 28040 11067
rect 27988 11024 28040 11033
rect 15568 10999 15620 11008
rect 15568 10965 15577 10999
rect 15577 10965 15611 10999
rect 15611 10965 15620 10999
rect 15568 10956 15620 10965
rect 15936 10956 15988 11008
rect 19340 10999 19392 11008
rect 19340 10965 19349 10999
rect 19349 10965 19383 10999
rect 19383 10965 19392 10999
rect 19340 10956 19392 10965
rect 10214 10854 10266 10906
rect 10278 10854 10330 10906
rect 10342 10854 10394 10906
rect 10406 10854 10458 10906
rect 10470 10854 10522 10906
rect 19478 10854 19530 10906
rect 19542 10854 19594 10906
rect 19606 10854 19658 10906
rect 19670 10854 19722 10906
rect 19734 10854 19786 10906
rect 17684 10752 17736 10804
rect 19340 10752 19392 10804
rect 19984 10752 20036 10804
rect 20904 10795 20956 10804
rect 20904 10761 20913 10795
rect 20913 10761 20947 10795
rect 20947 10761 20956 10795
rect 20904 10752 20956 10761
rect 27988 10752 28040 10804
rect 15936 10659 15988 10668
rect 15936 10625 15945 10659
rect 15945 10625 15979 10659
rect 15979 10625 15988 10659
rect 15936 10616 15988 10625
rect 17316 10684 17368 10736
rect 27620 10616 27672 10668
rect 20260 10591 20312 10600
rect 20260 10557 20269 10591
rect 20269 10557 20303 10591
rect 20303 10557 20312 10591
rect 20260 10548 20312 10557
rect 20444 10591 20496 10600
rect 20444 10557 20453 10591
rect 20453 10557 20487 10591
rect 20487 10557 20496 10591
rect 20444 10548 20496 10557
rect 25964 10591 26016 10600
rect 25964 10557 25973 10591
rect 25973 10557 26007 10591
rect 26007 10557 26016 10591
rect 25964 10548 26016 10557
rect 26240 10591 26292 10600
rect 26240 10557 26249 10591
rect 26249 10557 26283 10591
rect 26283 10557 26292 10591
rect 26240 10548 26292 10557
rect 1400 10412 1452 10464
rect 5582 10310 5634 10362
rect 5646 10310 5698 10362
rect 5710 10310 5762 10362
rect 5774 10310 5826 10362
rect 5838 10310 5890 10362
rect 14846 10310 14898 10362
rect 14910 10310 14962 10362
rect 14974 10310 15026 10362
rect 15038 10310 15090 10362
rect 15102 10310 15154 10362
rect 24110 10310 24162 10362
rect 24174 10310 24226 10362
rect 24238 10310 24290 10362
rect 24302 10310 24354 10362
rect 24366 10310 24418 10362
rect 16580 10208 16632 10260
rect 1768 10047 1820 10056
rect 1768 10013 1777 10047
rect 1777 10013 1811 10047
rect 1811 10013 1820 10047
rect 1768 10004 1820 10013
rect 28356 10140 28408 10192
rect 15568 10072 15620 10124
rect 20260 10072 20312 10124
rect 25320 10115 25372 10124
rect 25320 10081 25329 10115
rect 25329 10081 25363 10115
rect 25363 10081 25372 10115
rect 25320 10072 25372 10081
rect 3792 10004 3844 10056
rect 17684 10004 17736 10056
rect 25044 10004 25096 10056
rect 26976 10115 27028 10124
rect 26976 10081 26985 10115
rect 26985 10081 27019 10115
rect 27019 10081 27028 10115
rect 26976 10072 27028 10081
rect 1584 9868 1636 9920
rect 3608 9868 3660 9920
rect 17500 9868 17552 9920
rect 25044 9868 25096 9920
rect 27528 9911 27580 9920
rect 27528 9877 27537 9911
rect 27537 9877 27571 9911
rect 27571 9877 27580 9911
rect 27528 9868 27580 9877
rect 10214 9766 10266 9818
rect 10278 9766 10330 9818
rect 10342 9766 10394 9818
rect 10406 9766 10458 9818
rect 10470 9766 10522 9818
rect 19478 9766 19530 9818
rect 19542 9766 19594 9818
rect 19606 9766 19658 9818
rect 19670 9766 19722 9818
rect 19734 9766 19786 9818
rect 26240 9664 26292 9716
rect 3608 9639 3660 9648
rect 3608 9605 3617 9639
rect 3617 9605 3651 9639
rect 3651 9605 3660 9639
rect 3608 9596 3660 9605
rect 3792 9571 3844 9580
rect 3792 9537 3801 9571
rect 3801 9537 3835 9571
rect 3835 9537 3844 9571
rect 3792 9528 3844 9537
rect 3240 9503 3292 9512
rect 3240 9469 3249 9503
rect 3249 9469 3283 9503
rect 3283 9469 3292 9503
rect 3240 9460 3292 9469
rect 2964 9392 3016 9444
rect 26516 9528 26568 9580
rect 24860 9503 24912 9512
rect 24860 9469 24869 9503
rect 24869 9469 24903 9503
rect 24903 9469 24912 9503
rect 24860 9460 24912 9469
rect 25228 9460 25280 9512
rect 28264 9460 28316 9512
rect 25504 9324 25556 9376
rect 5582 9222 5634 9274
rect 5646 9222 5698 9274
rect 5710 9222 5762 9274
rect 5774 9222 5826 9274
rect 5838 9222 5890 9274
rect 14846 9222 14898 9274
rect 14910 9222 14962 9274
rect 14974 9222 15026 9274
rect 15038 9222 15090 9274
rect 15102 9222 15154 9274
rect 24110 9222 24162 9274
rect 24174 9222 24226 9274
rect 24238 9222 24290 9274
rect 24302 9222 24354 9274
rect 24366 9222 24418 9274
rect 25228 9163 25280 9172
rect 25228 9129 25237 9163
rect 25237 9129 25271 9163
rect 25271 9129 25280 9163
rect 25228 9120 25280 9129
rect 1400 9027 1452 9036
rect 1400 8993 1409 9027
rect 1409 8993 1443 9027
rect 1443 8993 1452 9027
rect 1400 8984 1452 8993
rect 1584 9027 1636 9036
rect 1584 8993 1593 9027
rect 1593 8993 1627 9027
rect 1627 8993 1636 9027
rect 1584 8984 1636 8993
rect 1860 9027 1912 9036
rect 1860 8993 1869 9027
rect 1869 8993 1903 9027
rect 1903 8993 1912 9027
rect 1860 8984 1912 8993
rect 26332 9027 26384 9036
rect 26332 8993 26341 9027
rect 26341 8993 26375 9027
rect 26375 8993 26384 9027
rect 26332 8984 26384 8993
rect 27528 8984 27580 9036
rect 24584 8916 24636 8968
rect 25044 8916 25096 8968
rect 29000 8848 29052 8900
rect 10214 8678 10266 8730
rect 10278 8678 10330 8730
rect 10342 8678 10394 8730
rect 10406 8678 10458 8730
rect 10470 8678 10522 8730
rect 19478 8678 19530 8730
rect 19542 8678 19594 8730
rect 19606 8678 19658 8730
rect 19670 8678 19722 8730
rect 19734 8678 19786 8730
rect 27160 8440 27212 8492
rect 2964 8415 3016 8424
rect 2964 8381 2973 8415
rect 2973 8381 3007 8415
rect 3007 8381 3016 8415
rect 2964 8372 3016 8381
rect 3148 8415 3200 8424
rect 3148 8381 3157 8415
rect 3157 8381 3191 8415
rect 3191 8381 3200 8415
rect 3148 8372 3200 8381
rect 25964 8415 26016 8424
rect 25964 8381 25973 8415
rect 25973 8381 26007 8415
rect 26007 8381 26016 8415
rect 25964 8372 26016 8381
rect 26240 8415 26292 8424
rect 26240 8381 26249 8415
rect 26249 8381 26283 8415
rect 26283 8381 26292 8415
rect 26424 8415 26476 8424
rect 26240 8372 26292 8381
rect 26424 8381 26433 8415
rect 26433 8381 26467 8415
rect 26467 8381 26476 8415
rect 26424 8372 26476 8381
rect 27896 8304 27948 8356
rect 1492 8236 1544 8288
rect 3424 8236 3476 8288
rect 27988 8279 28040 8288
rect 27988 8245 27997 8279
rect 27997 8245 28031 8279
rect 28031 8245 28040 8279
rect 27988 8236 28040 8245
rect 5582 8134 5634 8186
rect 5646 8134 5698 8186
rect 5710 8134 5762 8186
rect 5774 8134 5826 8186
rect 5838 8134 5890 8186
rect 14846 8134 14898 8186
rect 14910 8134 14962 8186
rect 14974 8134 15026 8186
rect 15038 8134 15090 8186
rect 15102 8134 15154 8186
rect 24110 8134 24162 8186
rect 24174 8134 24226 8186
rect 24238 8134 24290 8186
rect 24302 8134 24354 8186
rect 24366 8134 24418 8186
rect 1676 8032 1728 8084
rect 2964 8075 3016 8084
rect 2964 8041 2973 8075
rect 2973 8041 3007 8075
rect 3007 8041 3016 8075
rect 2964 8032 3016 8041
rect 3148 8032 3200 8084
rect 26240 8032 26292 8084
rect 27528 7939 27580 7948
rect 27528 7905 27537 7939
rect 27537 7905 27571 7939
rect 27571 7905 27580 7939
rect 27528 7896 27580 7905
rect 27988 7896 28040 7948
rect 2044 7871 2096 7880
rect 2044 7837 2053 7871
rect 2053 7837 2087 7871
rect 2087 7837 2096 7871
rect 2044 7828 2096 7837
rect 18696 7828 18748 7880
rect 9220 7760 9272 7812
rect 27896 7760 27948 7812
rect 3976 7692 4028 7744
rect 10214 7590 10266 7642
rect 10278 7590 10330 7642
rect 10342 7590 10394 7642
rect 10406 7590 10458 7642
rect 10470 7590 10522 7642
rect 19478 7590 19530 7642
rect 19542 7590 19594 7642
rect 19606 7590 19658 7642
rect 19670 7590 19722 7642
rect 19734 7590 19786 7642
rect 3976 7463 4028 7472
rect 3976 7429 3985 7463
rect 3985 7429 4019 7463
rect 4019 7429 4028 7463
rect 3976 7420 4028 7429
rect 25504 7420 25556 7472
rect 1492 7395 1544 7404
rect 1492 7361 1501 7395
rect 1501 7361 1535 7395
rect 1535 7361 1544 7395
rect 1492 7352 1544 7361
rect 24584 7395 24636 7404
rect 24584 7361 24593 7395
rect 24593 7361 24627 7395
rect 24627 7361 24636 7395
rect 24584 7352 24636 7361
rect 26424 7352 26476 7404
rect 1676 7327 1728 7336
rect 1676 7293 1685 7327
rect 1685 7293 1719 7327
rect 1719 7293 1728 7327
rect 1676 7284 1728 7293
rect 2872 7327 2924 7336
rect 2872 7293 2881 7327
rect 2881 7293 2915 7327
rect 2915 7293 2924 7327
rect 2872 7284 2924 7293
rect 3792 7327 3844 7336
rect 3792 7293 3801 7327
rect 3801 7293 3835 7327
rect 3835 7293 3844 7327
rect 3792 7284 3844 7293
rect 4160 7284 4212 7336
rect 26148 7327 26200 7336
rect 26148 7293 26157 7327
rect 26157 7293 26191 7327
rect 26191 7293 26200 7327
rect 26148 7284 26200 7293
rect 28172 7148 28224 7200
rect 5582 7046 5634 7098
rect 5646 7046 5698 7098
rect 5710 7046 5762 7098
rect 5774 7046 5826 7098
rect 5838 7046 5890 7098
rect 14846 7046 14898 7098
rect 14910 7046 14962 7098
rect 14974 7046 15026 7098
rect 15038 7046 15090 7098
rect 15102 7046 15154 7098
rect 24110 7046 24162 7098
rect 24174 7046 24226 7098
rect 24238 7046 24290 7098
rect 24302 7046 24354 7098
rect 24366 7046 24418 7098
rect 1676 6944 1728 6996
rect 3792 6987 3844 6996
rect 3792 6953 3801 6987
rect 3801 6953 3835 6987
rect 3835 6953 3844 6987
rect 3792 6944 3844 6953
rect 3424 6808 3476 6860
rect 24860 6808 24912 6860
rect 27528 6851 27580 6860
rect 27528 6817 27537 6851
rect 27537 6817 27571 6851
rect 27571 6817 27580 6851
rect 27528 6808 27580 6817
rect 28172 6851 28224 6860
rect 28172 6817 28181 6851
rect 28181 6817 28215 6851
rect 28215 6817 28224 6851
rect 28172 6808 28224 6817
rect 2044 6783 2096 6792
rect 2044 6749 2053 6783
rect 2053 6749 2087 6783
rect 2087 6749 2096 6783
rect 2044 6740 2096 6749
rect 6184 6740 6236 6792
rect 27804 6672 27856 6724
rect 10214 6502 10266 6554
rect 10278 6502 10330 6554
rect 10342 6502 10394 6554
rect 10406 6502 10458 6554
rect 10470 6502 10522 6554
rect 19478 6502 19530 6554
rect 19542 6502 19594 6554
rect 19606 6502 19658 6554
rect 19670 6502 19722 6554
rect 19734 6502 19786 6554
rect 27804 6443 27856 6452
rect 27804 6409 27813 6443
rect 27813 6409 27847 6443
rect 27847 6409 27856 6443
rect 27804 6400 27856 6409
rect 27620 6264 27672 6316
rect 2320 6239 2372 6248
rect 2320 6205 2329 6239
rect 2329 6205 2363 6239
rect 2363 6205 2372 6239
rect 2320 6196 2372 6205
rect 2596 6239 2648 6248
rect 2596 6205 2605 6239
rect 2605 6205 2639 6239
rect 2639 6205 2648 6239
rect 2596 6196 2648 6205
rect 26332 6060 26384 6112
rect 5582 5958 5634 6010
rect 5646 5958 5698 6010
rect 5710 5958 5762 6010
rect 5774 5958 5826 6010
rect 5838 5958 5890 6010
rect 14846 5958 14898 6010
rect 14910 5958 14962 6010
rect 14974 5958 15026 6010
rect 15038 5958 15090 6010
rect 15102 5958 15154 6010
rect 24110 5958 24162 6010
rect 24174 5958 24226 6010
rect 24238 5958 24290 6010
rect 24302 5958 24354 6010
rect 24366 5958 24418 6010
rect 2320 5856 2372 5908
rect 27620 5788 27672 5840
rect 26332 5763 26384 5772
rect 26332 5729 26341 5763
rect 26341 5729 26375 5763
rect 26375 5729 26384 5763
rect 26332 5720 26384 5729
rect 18604 5652 18656 5704
rect 22744 5652 22796 5704
rect 26516 5627 26568 5636
rect 26516 5593 26525 5627
rect 26525 5593 26559 5627
rect 26559 5593 26568 5627
rect 26516 5584 26568 5593
rect 28172 5627 28224 5636
rect 28172 5593 28181 5627
rect 28181 5593 28215 5627
rect 28215 5593 28224 5627
rect 28172 5584 28224 5593
rect 2872 5559 2924 5568
rect 2872 5525 2881 5559
rect 2881 5525 2915 5559
rect 2915 5525 2924 5559
rect 2872 5516 2924 5525
rect 10214 5414 10266 5466
rect 10278 5414 10330 5466
rect 10342 5414 10394 5466
rect 10406 5414 10458 5466
rect 10470 5414 10522 5466
rect 19478 5414 19530 5466
rect 19542 5414 19594 5466
rect 19606 5414 19658 5466
rect 19670 5414 19722 5466
rect 19734 5414 19786 5466
rect 26516 5312 26568 5364
rect 2872 5244 2924 5296
rect 18604 5176 18656 5228
rect 22744 5219 22796 5228
rect 22744 5185 22753 5219
rect 22753 5185 22787 5219
rect 22787 5185 22796 5219
rect 22744 5176 22796 5185
rect 3148 5151 3200 5160
rect 3148 5117 3157 5151
rect 3157 5117 3191 5151
rect 3191 5117 3200 5151
rect 3148 5108 3200 5117
rect 19340 5108 19392 5160
rect 27896 5176 27948 5228
rect 6276 4972 6328 5024
rect 17684 5015 17736 5024
rect 17684 4981 17693 5015
rect 17693 4981 17727 5015
rect 17727 4981 17736 5015
rect 17684 4972 17736 4981
rect 22836 5015 22888 5024
rect 22836 4981 22845 5015
rect 22845 4981 22879 5015
rect 22879 4981 22888 5015
rect 22836 4972 22888 4981
rect 5582 4870 5634 4922
rect 5646 4870 5698 4922
rect 5710 4870 5762 4922
rect 5774 4870 5826 4922
rect 5838 4870 5890 4922
rect 14846 4870 14898 4922
rect 14910 4870 14962 4922
rect 14974 4870 15026 4922
rect 15038 4870 15090 4922
rect 15102 4870 15154 4922
rect 24110 4870 24162 4922
rect 24174 4870 24226 4922
rect 24238 4870 24290 4922
rect 24302 4870 24354 4922
rect 24366 4870 24418 4922
rect 2780 4632 2832 4684
rect 3332 4632 3384 4684
rect 6276 4675 6328 4684
rect 6276 4641 6285 4675
rect 6285 4641 6319 4675
rect 6319 4641 6328 4675
rect 6276 4632 6328 4641
rect 21364 4675 21416 4684
rect 21364 4641 21373 4675
rect 21373 4641 21407 4675
rect 21407 4641 21416 4675
rect 21364 4632 21416 4641
rect 27436 4675 27488 4684
rect 27436 4641 27445 4675
rect 27445 4641 27479 4675
rect 27479 4641 27488 4675
rect 27436 4632 27488 4641
rect 28540 4632 28592 4684
rect 20720 4607 20772 4616
rect 20720 4573 20729 4607
rect 20729 4573 20763 4607
rect 20763 4573 20772 4607
rect 20720 4564 20772 4573
rect 28172 4607 28224 4616
rect 28172 4573 28181 4607
rect 28181 4573 28215 4607
rect 28215 4573 28224 4607
rect 28172 4564 28224 4573
rect 1400 4539 1452 4548
rect 1400 4505 1409 4539
rect 1409 4505 1443 4539
rect 1443 4505 1452 4539
rect 1400 4496 1452 4505
rect 2964 4496 3016 4548
rect 17684 4496 17736 4548
rect 20904 4539 20956 4548
rect 20904 4505 20913 4539
rect 20913 4505 20947 4539
rect 20947 4505 20956 4539
rect 20904 4496 20956 4505
rect 10214 4326 10266 4378
rect 10278 4326 10330 4378
rect 10342 4326 10394 4378
rect 10406 4326 10458 4378
rect 10470 4326 10522 4378
rect 19478 4326 19530 4378
rect 19542 4326 19594 4378
rect 19606 4326 19658 4378
rect 19670 4326 19722 4378
rect 19734 4326 19786 4378
rect 20904 4267 20956 4276
rect 20904 4233 20913 4267
rect 20913 4233 20947 4267
rect 20947 4233 20956 4267
rect 20904 4224 20956 4233
rect 1952 4088 2004 4140
rect 2780 4088 2832 4140
rect 5264 4131 5316 4140
rect 5264 4097 5273 4131
rect 5273 4097 5307 4131
rect 5307 4097 5316 4131
rect 5264 4088 5316 4097
rect 9220 4131 9272 4140
rect 9220 4097 9229 4131
rect 9229 4097 9263 4131
rect 9263 4097 9272 4131
rect 9220 4088 9272 4097
rect 12900 4088 12952 4140
rect 20628 4088 20680 4140
rect 22744 4088 22796 4140
rect 28172 4088 28224 4140
rect 2872 4063 2924 4072
rect 2872 4029 2881 4063
rect 2881 4029 2915 4063
rect 2915 4029 2924 4063
rect 2872 4020 2924 4029
rect 3056 4063 3108 4072
rect 3056 4029 3065 4063
rect 3065 4029 3099 4063
rect 3099 4029 3108 4063
rect 3056 4020 3108 4029
rect 3240 4020 3292 4072
rect 2964 3952 3016 4004
rect 12624 4020 12676 4072
rect 13176 4063 13228 4072
rect 13176 4029 13185 4063
rect 13185 4029 13219 4063
rect 13219 4029 13228 4063
rect 13176 4020 13228 4029
rect 13544 4063 13596 4072
rect 13544 4029 13553 4063
rect 13553 4029 13587 4063
rect 13587 4029 13596 4063
rect 13544 4020 13596 4029
rect 18052 4063 18104 4072
rect 18052 4029 18061 4063
rect 18061 4029 18095 4063
rect 18095 4029 18104 4063
rect 18052 4020 18104 4029
rect 18236 4020 18288 4072
rect 19616 4020 19668 4072
rect 19892 4063 19944 4072
rect 19892 4029 19901 4063
rect 19901 4029 19935 4063
rect 19935 4029 19944 4063
rect 19892 4020 19944 4029
rect 20720 4020 20772 4072
rect 5356 3927 5408 3936
rect 5356 3893 5365 3927
rect 5365 3893 5399 3927
rect 5399 3893 5408 3927
rect 5356 3884 5408 3893
rect 6368 3927 6420 3936
rect 6368 3893 6377 3927
rect 6377 3893 6411 3927
rect 6411 3893 6420 3927
rect 6368 3884 6420 3893
rect 8668 3884 8720 3936
rect 9312 3927 9364 3936
rect 9312 3893 9321 3927
rect 9321 3893 9355 3927
rect 9355 3893 9364 3927
rect 9312 3884 9364 3893
rect 11704 3884 11756 3936
rect 12900 3884 12952 3936
rect 19984 3884 20036 3936
rect 26792 3952 26844 4004
rect 26424 3927 26476 3936
rect 26424 3893 26433 3927
rect 26433 3893 26467 3927
rect 26467 3893 26476 3927
rect 26424 3884 26476 3893
rect 26976 3927 27028 3936
rect 26976 3893 26985 3927
rect 26985 3893 27019 3927
rect 27019 3893 27028 3927
rect 26976 3884 27028 3893
rect 5582 3782 5634 3834
rect 5646 3782 5698 3834
rect 5710 3782 5762 3834
rect 5774 3782 5826 3834
rect 5838 3782 5890 3834
rect 14846 3782 14898 3834
rect 14910 3782 14962 3834
rect 14974 3782 15026 3834
rect 15038 3782 15090 3834
rect 15102 3782 15154 3834
rect 24110 3782 24162 3834
rect 24174 3782 24226 3834
rect 24238 3782 24290 3834
rect 24302 3782 24354 3834
rect 24366 3782 24418 3834
rect 3056 3680 3108 3732
rect 5448 3680 5500 3732
rect 12624 3723 12676 3732
rect 12624 3689 12633 3723
rect 12633 3689 12667 3723
rect 12667 3689 12676 3723
rect 12624 3680 12676 3689
rect 13176 3723 13228 3732
rect 13176 3689 13185 3723
rect 13185 3689 13219 3723
rect 13219 3689 13228 3723
rect 13176 3680 13228 3689
rect 19892 3680 19944 3732
rect 5356 3587 5408 3596
rect 1676 3476 1728 3528
rect 2780 3519 2832 3528
rect 2780 3485 2789 3519
rect 2789 3485 2823 3519
rect 2823 3485 2832 3519
rect 2780 3476 2832 3485
rect 5356 3553 5365 3587
rect 5365 3553 5399 3587
rect 5399 3553 5408 3587
rect 5356 3544 5408 3553
rect 5908 3587 5960 3596
rect 5908 3553 5917 3587
rect 5917 3553 5951 3587
rect 5951 3553 5960 3587
rect 5908 3544 5960 3553
rect 9312 3587 9364 3596
rect 9312 3553 9321 3587
rect 9321 3553 9355 3587
rect 9355 3553 9364 3587
rect 9312 3544 9364 3553
rect 9680 3587 9732 3596
rect 9680 3553 9689 3587
rect 9689 3553 9723 3587
rect 9723 3553 9732 3587
rect 9680 3544 9732 3553
rect 19294 3544 19346 3596
rect 5172 3519 5224 3528
rect 5172 3485 5181 3519
rect 5181 3485 5215 3519
rect 5215 3485 5224 3519
rect 5172 3476 5224 3485
rect 11520 3476 11572 3528
rect 13084 3519 13136 3528
rect 13084 3485 13093 3519
rect 13093 3485 13127 3519
rect 13127 3485 13136 3519
rect 13084 3476 13136 3485
rect 14648 3519 14700 3528
rect 14648 3485 14657 3519
rect 14657 3485 14691 3519
rect 14691 3485 14700 3519
rect 14648 3476 14700 3485
rect 16304 3519 16356 3528
rect 14280 3408 14332 3460
rect 16304 3485 16313 3519
rect 16313 3485 16347 3519
rect 16347 3485 16356 3519
rect 16304 3476 16356 3485
rect 16672 3476 16724 3528
rect 20628 3612 20680 3664
rect 21916 3587 21968 3596
rect 21916 3553 21925 3587
rect 21925 3553 21959 3587
rect 21959 3553 21968 3587
rect 21916 3544 21968 3553
rect 19616 3476 19668 3528
rect 21272 3519 21324 3528
rect 21272 3485 21281 3519
rect 21281 3485 21315 3519
rect 21315 3485 21324 3519
rect 21272 3476 21324 3485
rect 24032 3476 24084 3528
rect 28448 3612 28500 3664
rect 26976 3544 27028 3596
rect 27528 3587 27580 3596
rect 27528 3553 27537 3587
rect 27537 3553 27571 3587
rect 27571 3553 27580 3587
rect 27528 3544 27580 3553
rect 1860 3340 1912 3392
rect 4160 3340 4212 3392
rect 8852 3340 8904 3392
rect 14464 3340 14516 3392
rect 16856 3340 16908 3392
rect 19340 3340 19392 3392
rect 27068 3408 27120 3460
rect 26976 3340 27028 3392
rect 10214 3238 10266 3290
rect 10278 3238 10330 3290
rect 10342 3238 10394 3290
rect 10406 3238 10458 3290
rect 10470 3238 10522 3290
rect 19478 3238 19530 3290
rect 19542 3238 19594 3290
rect 19606 3238 19658 3290
rect 19670 3238 19722 3290
rect 19734 3238 19786 3290
rect 664 3136 716 3188
rect 2596 3136 2648 3188
rect 1860 3111 1912 3120
rect 1860 3077 1869 3111
rect 1869 3077 1903 3111
rect 1903 3077 1912 3111
rect 1860 3068 1912 3077
rect 1952 3068 2004 3120
rect 13084 3136 13136 3188
rect 19984 3136 20036 3188
rect 27068 3179 27120 3188
rect 4160 3111 4212 3120
rect 4160 3077 4169 3111
rect 4169 3077 4203 3111
rect 4203 3077 4212 3111
rect 4160 3068 4212 3077
rect 8852 3111 8904 3120
rect 8852 3077 8861 3111
rect 8861 3077 8895 3111
rect 8895 3077 8904 3111
rect 8852 3068 8904 3077
rect 11704 3111 11756 3120
rect 11704 3077 11713 3111
rect 11713 3077 11747 3111
rect 11747 3077 11756 3111
rect 11704 3068 11756 3077
rect 14464 3111 14516 3120
rect 14464 3077 14473 3111
rect 14473 3077 14507 3111
rect 14507 3077 14516 3111
rect 14464 3068 14516 3077
rect 16856 3111 16908 3120
rect 16856 3077 16865 3111
rect 16865 3077 16899 3111
rect 16899 3077 16908 3111
rect 16856 3068 16908 3077
rect 19340 3068 19392 3120
rect 27068 3145 27077 3179
rect 27077 3145 27111 3179
rect 27111 3145 27120 3179
rect 27068 3136 27120 3145
rect 28080 3068 28132 3120
rect 1676 3043 1728 3052
rect 1676 3009 1685 3043
rect 1685 3009 1719 3043
rect 1719 3009 1728 3043
rect 1676 3000 1728 3009
rect 6368 3043 6420 3052
rect 6368 3009 6377 3043
rect 6377 3009 6411 3043
rect 6411 3009 6420 3043
rect 6368 3000 6420 3009
rect 8668 3043 8720 3052
rect 8668 3009 8677 3043
rect 8677 3009 8711 3043
rect 8711 3009 8720 3043
rect 8668 3000 8720 3009
rect 11520 3043 11572 3052
rect 11520 3009 11529 3043
rect 11529 3009 11563 3043
rect 11563 3009 11572 3043
rect 11520 3000 11572 3009
rect 14280 3043 14332 3052
rect 14280 3009 14289 3043
rect 14289 3009 14323 3043
rect 14323 3009 14332 3043
rect 14280 3000 14332 3009
rect 16672 3043 16724 3052
rect 16672 3009 16681 3043
rect 16681 3009 16715 3043
rect 16715 3009 16724 3043
rect 16672 3000 16724 3009
rect 21272 3000 21324 3052
rect 2780 2975 2832 2984
rect 2780 2941 2789 2975
rect 2789 2941 2823 2975
rect 2823 2941 2832 2975
rect 2780 2932 2832 2941
rect 3976 2975 4028 2984
rect 3976 2941 3985 2975
rect 3985 2941 4019 2975
rect 4019 2941 4028 2975
rect 3976 2932 4028 2941
rect 4528 2975 4580 2984
rect 4528 2941 4537 2975
rect 4537 2941 4571 2975
rect 4571 2941 4580 2975
rect 4528 2932 4580 2941
rect 6552 2975 6604 2984
rect 6552 2941 6561 2975
rect 6561 2941 6595 2975
rect 6595 2941 6604 2975
rect 6552 2932 6604 2941
rect 6460 2864 6512 2916
rect 8392 2932 8444 2984
rect 14740 2975 14792 2984
rect 10968 2864 11020 2916
rect 14740 2941 14749 2975
rect 14749 2941 14783 2975
rect 14783 2941 14792 2975
rect 14740 2932 14792 2941
rect 19432 2975 19484 2984
rect 19432 2941 19441 2975
rect 19441 2941 19475 2975
rect 19475 2941 19484 2975
rect 19432 2932 19484 2941
rect 19984 2975 20036 2984
rect 19984 2941 19993 2975
rect 19993 2941 20027 2975
rect 20027 2941 20036 2975
rect 19984 2932 20036 2941
rect 16764 2864 16816 2916
rect 2596 2796 2648 2848
rect 3148 2796 3200 2848
rect 16028 2796 16080 2848
rect 16304 2796 16356 2848
rect 22836 3000 22888 3052
rect 24032 3043 24084 3052
rect 24032 3009 24041 3043
rect 24041 3009 24075 3043
rect 24075 3009 24084 3043
rect 24032 3000 24084 3009
rect 26976 3043 27028 3052
rect 26976 3009 26985 3043
rect 26985 3009 27019 3043
rect 27019 3009 27028 3043
rect 26976 3000 27028 3009
rect 27712 3000 27764 3052
rect 25136 2975 25188 2984
rect 25136 2941 25145 2975
rect 25145 2941 25179 2975
rect 25179 2941 25188 2975
rect 25136 2932 25188 2941
rect 26240 2796 26292 2848
rect 5582 2694 5634 2746
rect 5646 2694 5698 2746
rect 5710 2694 5762 2746
rect 5774 2694 5826 2746
rect 5838 2694 5890 2746
rect 14846 2694 14898 2746
rect 14910 2694 14962 2746
rect 14974 2694 15026 2746
rect 15038 2694 15090 2746
rect 15102 2694 15154 2746
rect 24110 2694 24162 2746
rect 24174 2694 24226 2746
rect 24238 2694 24290 2746
rect 24302 2694 24354 2746
rect 24366 2694 24418 2746
rect 2872 2635 2924 2644
rect 2872 2601 2881 2635
rect 2881 2601 2915 2635
rect 2915 2601 2924 2635
rect 2872 2592 2924 2601
rect 3976 2592 4028 2644
rect 5172 2592 5224 2644
rect 6552 2592 6604 2644
rect 9496 2635 9548 2644
rect 9496 2601 9505 2635
rect 9505 2601 9539 2635
rect 9539 2601 9548 2635
rect 9496 2592 9548 2601
rect 16856 2635 16908 2644
rect 16856 2601 16865 2635
rect 16865 2601 16899 2635
rect 16899 2601 16908 2635
rect 16856 2592 16908 2601
rect 17500 2635 17552 2644
rect 17500 2601 17509 2635
rect 17509 2601 17543 2635
rect 17543 2601 17552 2635
rect 17500 2592 17552 2601
rect 19432 2635 19484 2644
rect 19432 2601 19441 2635
rect 19441 2601 19475 2635
rect 19475 2601 19484 2635
rect 19432 2592 19484 2601
rect 20444 2592 20496 2644
rect 3424 2524 3476 2576
rect 25320 2524 25372 2576
rect 25964 2499 26016 2508
rect 25964 2465 25973 2499
rect 25973 2465 26007 2499
rect 26007 2465 26016 2499
rect 25964 2456 26016 2465
rect 26240 2499 26292 2508
rect 26240 2465 26249 2499
rect 26249 2465 26283 2499
rect 26283 2465 26292 2499
rect 26424 2499 26476 2508
rect 26240 2456 26292 2465
rect 26424 2465 26433 2499
rect 26433 2465 26467 2499
rect 26467 2465 26476 2499
rect 26424 2456 26476 2465
rect 6184 2388 6236 2440
rect 16028 2388 16080 2440
rect 16120 2388 16172 2440
rect 17408 2388 17460 2440
rect 27068 2388 27120 2440
rect 9036 2320 9088 2372
rect 10214 2150 10266 2202
rect 10278 2150 10330 2202
rect 10342 2150 10394 2202
rect 10406 2150 10458 2202
rect 10470 2150 10522 2202
rect 19478 2150 19530 2202
rect 19542 2150 19594 2202
rect 19606 2150 19658 2202
rect 19670 2150 19722 2202
rect 19734 2150 19786 2202
<< metal2 >>
rect -10 49200 102 50000
rect 634 49200 746 50000
rect 1278 49200 1390 50000
rect 1922 49314 2034 50000
rect 1922 49286 2360 49314
rect 1922 49200 2034 49286
rect 676 45554 704 49200
rect 1320 46442 1348 49200
rect 1676 47048 1728 47054
rect 1676 46990 1728 46996
rect 1688 46578 1716 46990
rect 1676 46572 1728 46578
rect 1676 46514 1728 46520
rect 2136 46504 2188 46510
rect 2136 46446 2188 46452
rect 1308 46436 1360 46442
rect 1308 46378 1360 46384
rect 2148 46170 2176 46446
rect 2332 46442 2360 49286
rect 2566 49200 2678 50000
rect 3210 49200 3322 50000
rect 4066 49736 4122 49745
rect 4066 49671 4122 49680
rect 2608 46918 2636 49200
rect 3608 47048 3660 47054
rect 3608 46990 3660 46996
rect 3792 47048 3844 47054
rect 3792 46990 3844 46996
rect 2596 46912 2648 46918
rect 2596 46854 2648 46860
rect 3056 46912 3108 46918
rect 3056 46854 3108 46860
rect 2320 46436 2372 46442
rect 2320 46378 2372 46384
rect 2136 46164 2188 46170
rect 2136 46106 2188 46112
rect 1584 45960 1636 45966
rect 1584 45902 1636 45908
rect 32 45526 704 45554
rect 32 45354 60 45526
rect 1596 45490 1624 45902
rect 1584 45484 1636 45490
rect 1584 45426 1636 45432
rect 1952 45416 2004 45422
rect 1952 45358 2004 45364
rect 20 45348 72 45354
rect 20 45290 72 45296
rect 1964 45082 1992 45358
rect 1952 45076 2004 45082
rect 1952 45018 2004 45024
rect 1952 44872 2004 44878
rect 1952 44814 2004 44820
rect 1400 44192 1452 44198
rect 1400 44134 1452 44140
rect 1584 44192 1636 44198
rect 1584 44134 1636 44140
rect 1412 43858 1440 44134
rect 1596 43858 1624 44134
rect 1400 43852 1452 43858
rect 1400 43794 1452 43800
rect 1584 43852 1636 43858
rect 1584 43794 1636 43800
rect 1768 42696 1820 42702
rect 1768 42638 1820 42644
rect 1398 42256 1454 42265
rect 1398 42191 1454 42200
rect 1412 41682 1440 42191
rect 1584 42016 1636 42022
rect 1584 41958 1636 41964
rect 1400 41676 1452 41682
rect 1400 41618 1452 41624
rect 1596 41138 1624 41958
rect 1780 41682 1808 42638
rect 1768 41676 1820 41682
rect 1768 41618 1820 41624
rect 1584 41132 1636 41138
rect 1584 41074 1636 41080
rect 1676 38752 1728 38758
rect 1676 38694 1728 38700
rect 1688 38418 1716 38694
rect 1676 38412 1728 38418
rect 1676 38354 1728 38360
rect 1964 37890 1992 44814
rect 2870 44296 2926 44305
rect 2870 44231 2926 44240
rect 2780 44192 2832 44198
rect 2780 44134 2832 44140
rect 2792 43382 2820 44134
rect 2884 43858 2912 44231
rect 2872 43852 2924 43858
rect 2872 43794 2924 43800
rect 2780 43376 2832 43382
rect 2780 43318 2832 43324
rect 3068 43246 3096 46854
rect 3620 46578 3648 46990
rect 3608 46572 3660 46578
rect 3608 46514 3660 46520
rect 3804 46034 3832 46990
rect 4080 46034 4108 49671
rect 4498 49200 4610 50000
rect 5142 49200 5254 50000
rect 5786 49314 5898 50000
rect 5786 49286 6132 49314
rect 5786 49200 5898 49286
rect 5582 47356 5890 47376
rect 5582 47354 5588 47356
rect 5644 47354 5668 47356
rect 5724 47354 5748 47356
rect 5804 47354 5828 47356
rect 5884 47354 5890 47356
rect 5644 47302 5646 47354
rect 5826 47302 5828 47354
rect 5582 47300 5588 47302
rect 5644 47300 5668 47302
rect 5724 47300 5748 47302
rect 5804 47300 5828 47302
rect 5884 47300 5890 47302
rect 5582 47280 5890 47300
rect 6104 47054 6132 49286
rect 6430 49200 6542 50000
rect 7074 49200 7186 50000
rect 7718 49200 7830 50000
rect 8362 49200 8474 50000
rect 9650 49200 9762 50000
rect 10294 49314 10406 50000
rect 10152 49286 10406 49314
rect 6092 47048 6144 47054
rect 6092 46990 6144 46996
rect 6472 47002 6500 49200
rect 7840 47048 7892 47054
rect 6472 46974 6684 47002
rect 7840 46990 7892 46996
rect 6656 46918 6684 46974
rect 6552 46912 6604 46918
rect 6552 46854 6604 46860
rect 6644 46912 6696 46918
rect 6644 46854 6696 46860
rect 7288 46912 7340 46918
rect 7288 46854 7340 46860
rect 4160 46504 4212 46510
rect 4160 46446 4212 46452
rect 4172 46170 4200 46446
rect 5582 46268 5890 46288
rect 5582 46266 5588 46268
rect 5644 46266 5668 46268
rect 5724 46266 5748 46268
rect 5804 46266 5828 46268
rect 5884 46266 5890 46268
rect 5644 46214 5646 46266
rect 5826 46214 5828 46266
rect 5582 46212 5588 46214
rect 5644 46212 5668 46214
rect 5724 46212 5748 46214
rect 5804 46212 5828 46214
rect 5884 46212 5890 46214
rect 5582 46192 5890 46212
rect 4160 46164 4212 46170
rect 4160 46106 4212 46112
rect 4988 46096 5040 46102
rect 4988 46038 5040 46044
rect 3792 46028 3844 46034
rect 3792 45970 3844 45976
rect 4068 46028 4120 46034
rect 4068 45970 4120 45976
rect 4528 45892 4580 45898
rect 4528 45834 4580 45840
rect 4540 45558 4568 45834
rect 4528 45552 4580 45558
rect 4528 45494 4580 45500
rect 3238 44976 3294 44985
rect 3238 44911 3294 44920
rect 2964 43240 3016 43246
rect 2964 43182 3016 43188
rect 3056 43240 3108 43246
rect 3056 43182 3108 43188
rect 2976 42770 3004 43182
rect 2964 42764 3016 42770
rect 2964 42706 3016 42712
rect 3148 42696 3200 42702
rect 3148 42638 3200 42644
rect 2780 42152 2832 42158
rect 2780 42094 2832 42100
rect 2792 41585 2820 42094
rect 2778 41576 2834 41585
rect 2778 41511 2834 41520
rect 3056 41540 3108 41546
rect 3056 41482 3108 41488
rect 2044 41064 2096 41070
rect 2044 41006 2096 41012
rect 2056 40730 2084 41006
rect 3068 40730 3096 41482
rect 2044 40724 2096 40730
rect 2044 40666 2096 40672
rect 3056 40724 3108 40730
rect 3056 40666 3108 40672
rect 2778 38856 2834 38865
rect 2778 38791 2834 38800
rect 2792 38418 2820 38791
rect 2780 38412 2832 38418
rect 2780 38354 2832 38360
rect 2136 38276 2188 38282
rect 2136 38218 2188 38224
rect 2148 38010 2176 38218
rect 2136 38004 2188 38010
rect 2136 37946 2188 37952
rect 1964 37862 2176 37890
rect 1398 37496 1454 37505
rect 1398 37431 1454 37440
rect 1412 37262 1440 37431
rect 1400 37256 1452 37262
rect 1400 37198 1452 37204
rect 1858 36816 1914 36825
rect 1858 36751 1860 36760
rect 1912 36751 1914 36760
rect 2044 36780 2096 36786
rect 1860 36722 1912 36728
rect 2044 36722 2096 36728
rect 2056 35894 2084 36722
rect 1964 35866 2084 35894
rect 1400 35488 1452 35494
rect 1400 35430 1452 35436
rect 1412 35154 1440 35430
rect 1400 35148 1452 35154
rect 1400 35090 1452 35096
rect 1492 34944 1544 34950
rect 1492 34886 1544 34892
rect 1400 32224 1452 32230
rect 1400 32166 1452 32172
rect 1412 31890 1440 32166
rect 1400 31884 1452 31890
rect 1400 31826 1452 31832
rect 1400 30252 1452 30258
rect 1400 30194 1452 30200
rect 1412 30025 1440 30194
rect 1398 30016 1454 30025
rect 1398 29951 1454 29960
rect 1400 28076 1452 28082
rect 1400 28018 1452 28024
rect 1412 27985 1440 28018
rect 1398 27976 1454 27985
rect 1398 27911 1454 27920
rect 1400 25696 1452 25702
rect 1400 25638 1452 25644
rect 1412 25362 1440 25638
rect 1400 25356 1452 25362
rect 1400 25298 1452 25304
rect 1398 25256 1454 25265
rect 1398 25191 1454 25200
rect 1412 24206 1440 25191
rect 1400 24200 1452 24206
rect 1400 24142 1452 24148
rect 1400 19848 1452 19854
rect 1400 19790 1452 19796
rect 1412 19378 1440 19790
rect 1400 19372 1452 19378
rect 1400 19314 1452 19320
rect 1400 18080 1452 18086
rect 1400 18022 1452 18028
rect 1412 17746 1440 18022
rect 1400 17740 1452 17746
rect 1400 17682 1452 17688
rect 1400 15496 1452 15502
rect 1400 15438 1452 15444
rect 1412 14482 1440 15438
rect 1400 14476 1452 14482
rect 1400 14418 1452 14424
rect 1504 13954 1532 34886
rect 1766 34776 1822 34785
rect 1766 34711 1822 34720
rect 1780 34678 1808 34711
rect 1964 34678 1992 35866
rect 1768 34672 1820 34678
rect 1768 34614 1820 34620
rect 1952 34672 2004 34678
rect 1952 34614 2004 34620
rect 1858 32056 1914 32065
rect 1858 31991 1914 32000
rect 1872 31890 1900 31991
rect 1860 31884 1912 31890
rect 1860 31826 1912 31832
rect 1584 31748 1636 31754
rect 1584 31690 1636 31696
rect 1596 31482 1624 31690
rect 1584 31476 1636 31482
rect 1584 31418 1636 31424
rect 1584 25220 1636 25226
rect 1584 25162 1636 25168
rect 1596 24954 1624 25162
rect 1584 24948 1636 24954
rect 1584 24890 1636 24896
rect 1768 24812 1820 24818
rect 1768 24754 1820 24760
rect 1780 24614 1808 24754
rect 1768 24608 1820 24614
rect 1768 24550 1820 24556
rect 1584 24064 1636 24070
rect 1584 24006 1636 24012
rect 1596 23866 1624 24006
rect 1584 23860 1636 23866
rect 1584 23802 1636 23808
rect 1584 22024 1636 22030
rect 1584 21966 1636 21972
rect 1596 21010 1624 21966
rect 1584 21004 1636 21010
rect 1584 20946 1636 20952
rect 1584 19304 1636 19310
rect 1584 19246 1636 19252
rect 1596 18970 1624 19246
rect 1584 18964 1636 18970
rect 1584 18906 1636 18912
rect 1676 17604 1728 17610
rect 1676 17546 1728 17552
rect 1688 17338 1716 17546
rect 1676 17332 1728 17338
rect 1676 17274 1728 17280
rect 1780 17202 1808 24550
rect 1860 19304 1912 19310
rect 1860 19246 1912 19252
rect 1872 19145 1900 19246
rect 1858 19136 1914 19145
rect 1858 19071 1914 19080
rect 1768 17196 1820 17202
rect 1768 17138 1820 17144
rect 1584 14816 1636 14822
rect 1584 14758 1636 14764
rect 1596 14482 1624 14758
rect 1584 14476 1636 14482
rect 1584 14418 1636 14424
rect 1504 13926 1624 13954
rect 1492 13864 1544 13870
rect 1492 13806 1544 13812
rect 1504 12850 1532 13806
rect 1492 12844 1544 12850
rect 1492 12786 1544 12792
rect 1492 12232 1544 12238
rect 1492 12174 1544 12180
rect 1504 11762 1532 12174
rect 1492 11756 1544 11762
rect 1492 11698 1544 11704
rect 1400 10464 1452 10470
rect 1400 10406 1452 10412
rect 1412 9042 1440 10406
rect 1596 10010 1624 13926
rect 1676 13864 1728 13870
rect 1676 13806 1728 13812
rect 1688 13530 1716 13806
rect 1676 13524 1728 13530
rect 1676 13466 1728 13472
rect 1780 10062 1808 17138
rect 1964 16574 1992 34614
rect 2148 26234 2176 37862
rect 2228 37868 2280 37874
rect 2228 37810 2280 37816
rect 2240 34746 2268 37810
rect 2780 37188 2832 37194
rect 2780 37130 2832 37136
rect 2792 36922 2820 37130
rect 2780 36916 2832 36922
rect 2780 36858 2832 36864
rect 2320 36576 2372 36582
rect 2320 36518 2372 36524
rect 2228 34740 2280 34746
rect 2228 34682 2280 34688
rect 2228 31340 2280 31346
rect 2228 31282 2280 31288
rect 2056 26206 2176 26234
rect 2056 24750 2084 26206
rect 2044 24744 2096 24750
rect 2044 24686 2096 24692
rect 2044 21344 2096 21350
rect 2044 21286 2096 21292
rect 2056 20874 2084 21286
rect 2044 20868 2096 20874
rect 2044 20810 2096 20816
rect 2240 18766 2268 31282
rect 2332 23798 2360 36518
rect 2778 36136 2834 36145
rect 2778 36071 2834 36080
rect 2792 35154 2820 36071
rect 2780 35148 2832 35154
rect 2780 35090 2832 35096
rect 2688 33992 2740 33998
rect 2688 33934 2740 33940
rect 2320 23792 2372 23798
rect 2320 23734 2372 23740
rect 2700 22778 2728 33934
rect 2778 25936 2834 25945
rect 2778 25871 2834 25880
rect 2792 25362 2820 25871
rect 2780 25356 2832 25362
rect 2780 25298 2832 25304
rect 3160 24682 3188 42638
rect 3252 41070 3280 44911
rect 3884 42152 3936 42158
rect 3884 42094 3936 42100
rect 4620 42152 4672 42158
rect 4620 42094 4672 42100
rect 3896 41818 3924 42094
rect 4632 41818 4660 42094
rect 3884 41812 3936 41818
rect 3884 41754 3936 41760
rect 4620 41812 4672 41818
rect 4620 41754 4672 41760
rect 3240 41064 3292 41070
rect 3240 41006 3292 41012
rect 3240 37664 3292 37670
rect 3240 37606 3292 37612
rect 3252 37262 3280 37606
rect 3240 37256 3292 37262
rect 3240 37198 3292 37204
rect 3608 35488 3660 35494
rect 3608 35430 3660 35436
rect 3620 34610 3648 35430
rect 3608 34604 3660 34610
rect 3608 34546 3660 34552
rect 3424 34536 3476 34542
rect 3424 34478 3476 34484
rect 3436 34202 3464 34478
rect 3424 34196 3476 34202
rect 3424 34138 3476 34144
rect 3330 33416 3386 33425
rect 3330 33351 3386 33360
rect 3344 32026 3372 33351
rect 3332 32020 3384 32026
rect 3332 31962 3384 31968
rect 5000 25226 5028 46038
rect 5448 45484 5500 45490
rect 5448 45426 5500 45432
rect 5460 45354 5488 45426
rect 5448 45348 5500 45354
rect 5448 45290 5500 45296
rect 4712 25220 4764 25226
rect 4712 25162 4764 25168
rect 4988 25220 5040 25226
rect 4988 25162 5040 25168
rect 4068 24744 4120 24750
rect 4068 24686 4120 24692
rect 3148 24676 3200 24682
rect 3148 24618 3200 24624
rect 3160 23526 3188 24618
rect 3148 23520 3200 23526
rect 3148 23462 3200 23468
rect 2688 22772 2740 22778
rect 2688 22714 2740 22720
rect 3700 20868 3752 20874
rect 3700 20810 3752 20816
rect 2320 20392 2372 20398
rect 2320 20334 2372 20340
rect 2872 20392 2924 20398
rect 2872 20334 2924 20340
rect 2964 20392 3016 20398
rect 2964 20334 3016 20340
rect 2332 20058 2360 20334
rect 2884 20058 2912 20334
rect 2320 20052 2372 20058
rect 2320 19994 2372 20000
rect 2872 20052 2924 20058
rect 2872 19994 2924 20000
rect 2976 19825 3004 20334
rect 2962 19816 3018 19825
rect 2962 19751 3018 19760
rect 2964 19712 3016 19718
rect 2964 19654 3016 19660
rect 2228 18760 2280 18766
rect 2228 18702 2280 18708
rect 2412 18760 2464 18766
rect 2412 18702 2464 18708
rect 2424 18465 2452 18702
rect 2410 18456 2466 18465
rect 2410 18391 2466 18400
rect 2778 17776 2834 17785
rect 2778 17711 2780 17720
rect 2832 17711 2834 17720
rect 2780 17682 2832 17688
rect 1964 16546 2084 16574
rect 1860 14476 1912 14482
rect 1860 14418 1912 14424
rect 1872 14385 1900 14418
rect 1858 14376 1914 14385
rect 1858 14311 1914 14320
rect 1952 13864 2004 13870
rect 1952 13806 2004 13812
rect 1964 13705 1992 13806
rect 1950 13696 2006 13705
rect 1950 13631 2006 13640
rect 1860 11688 1912 11694
rect 1952 11688 2004 11694
rect 1860 11630 1912 11636
rect 1950 11656 1952 11665
rect 2004 11656 2006 11665
rect 1872 11354 1900 11630
rect 1950 11591 2006 11600
rect 1860 11348 1912 11354
rect 1860 11290 1912 11296
rect 2056 11150 2084 16546
rect 2778 15736 2834 15745
rect 2778 15671 2834 15680
rect 2136 15020 2188 15026
rect 2136 14962 2188 14968
rect 2148 13326 2176 14962
rect 2792 14958 2820 15671
rect 2780 14952 2832 14958
rect 2780 14894 2832 14900
rect 2136 13320 2188 13326
rect 2136 13262 2188 13268
rect 2780 13320 2832 13326
rect 2780 13262 2832 13268
rect 2044 11144 2096 11150
rect 1964 11092 2044 11098
rect 1964 11086 2096 11092
rect 1964 11070 2084 11086
rect 1768 10056 1820 10062
rect 1596 9982 1716 10010
rect 1768 9998 1820 10004
rect 1584 9920 1636 9926
rect 1584 9862 1636 9868
rect 1596 9042 1624 9862
rect 1400 9036 1452 9042
rect 1400 8978 1452 8984
rect 1584 9036 1636 9042
rect 1584 8978 1636 8984
rect 1492 8288 1544 8294
rect 1492 8230 1544 8236
rect 1504 7410 1532 8230
rect 1688 8090 1716 9982
rect 1860 9036 1912 9042
rect 1860 8978 1912 8984
rect 1872 8945 1900 8978
rect 1858 8936 1914 8945
rect 1858 8871 1914 8880
rect 1676 8084 1728 8090
rect 1676 8026 1728 8032
rect 1492 7404 1544 7410
rect 1492 7346 1544 7352
rect 1676 7336 1728 7342
rect 1676 7278 1728 7284
rect 1688 7002 1716 7278
rect 1676 6996 1728 7002
rect 1676 6938 1728 6944
rect 1400 4548 1452 4554
rect 1400 4490 1452 4496
rect 1412 4185 1440 4490
rect 1398 4176 1454 4185
rect 1964 4146 1992 11070
rect 2044 7880 2096 7886
rect 2044 7822 2096 7828
rect 2056 6798 2084 7822
rect 2044 6792 2096 6798
rect 2044 6734 2096 6740
rect 2320 6248 2372 6254
rect 2320 6190 2372 6196
rect 2596 6248 2648 6254
rect 2596 6190 2648 6196
rect 2332 5914 2360 6190
rect 2320 5908 2372 5914
rect 2320 5850 2372 5856
rect 1398 4111 1454 4120
rect 1952 4140 2004 4146
rect 1952 4082 2004 4088
rect 1676 3528 1728 3534
rect 1676 3470 1728 3476
rect 664 3188 716 3194
rect 664 3130 716 3136
rect 676 800 704 3130
rect 1688 3058 1716 3470
rect 1860 3392 1912 3398
rect 1860 3334 1912 3340
rect 1872 3126 1900 3334
rect 1964 3126 1992 4082
rect 2608 3194 2636 6190
rect 2792 4842 2820 13262
rect 2976 9450 3004 19654
rect 3330 12336 3386 12345
rect 3330 12271 3386 12280
rect 3344 12170 3372 12271
rect 3332 12164 3384 12170
rect 3332 12106 3384 12112
rect 3608 9920 3660 9926
rect 3608 9862 3660 9868
rect 3620 9654 3648 9862
rect 3608 9648 3660 9654
rect 3608 9590 3660 9596
rect 3240 9512 3292 9518
rect 3240 9454 3292 9460
rect 2964 9444 3016 9450
rect 2964 9386 3016 9392
rect 2964 8424 3016 8430
rect 2964 8366 3016 8372
rect 3148 8424 3200 8430
rect 3148 8366 3200 8372
rect 2976 8090 3004 8366
rect 3160 8090 3188 8366
rect 2964 8084 3016 8090
rect 2964 8026 3016 8032
rect 3148 8084 3200 8090
rect 3148 8026 3200 8032
rect 2870 7576 2926 7585
rect 2870 7511 2926 7520
rect 2884 7342 2912 7511
rect 2872 7336 2924 7342
rect 2872 7278 2924 7284
rect 2872 5568 2924 5574
rect 2872 5510 2924 5516
rect 2884 5302 2912 5510
rect 2872 5296 2924 5302
rect 2872 5238 2924 5244
rect 3148 5160 3200 5166
rect 3148 5102 3200 5108
rect 2700 4814 2820 4842
rect 2700 4026 2728 4814
rect 2780 4684 2832 4690
rect 2780 4626 2832 4632
rect 2792 4146 2820 4626
rect 2964 4548 3016 4554
rect 2964 4490 3016 4496
rect 2780 4140 2832 4146
rect 2780 4082 2832 4088
rect 2872 4072 2924 4078
rect 2700 3998 2820 4026
rect 2872 4014 2924 4020
rect 2792 3534 2820 3998
rect 2780 3528 2832 3534
rect 2780 3470 2832 3476
rect 2596 3188 2648 3194
rect 2596 3130 2648 3136
rect 1860 3120 1912 3126
rect 1860 3062 1912 3068
rect 1952 3120 2004 3126
rect 1952 3062 2004 3068
rect 1676 3052 1728 3058
rect 1676 2994 1728 3000
rect 2780 2984 2832 2990
rect 2780 2926 2832 2932
rect 2596 2848 2648 2854
rect 2792 2825 2820 2926
rect 2596 2790 2648 2796
rect 2778 2816 2834 2825
rect 2608 800 2636 2790
rect 2778 2751 2834 2760
rect 2884 2650 2912 4014
rect 2976 4010 3004 4490
rect 3056 4072 3108 4078
rect 3056 4014 3108 4020
rect 2964 4004 3016 4010
rect 2964 3946 3016 3952
rect 3068 3738 3096 4014
rect 3056 3732 3108 3738
rect 3056 3674 3108 3680
rect 3160 2854 3188 5102
rect 3252 4162 3280 9454
rect 3424 8288 3476 8294
rect 3422 8256 3424 8265
rect 3476 8256 3478 8265
rect 3422 8191 3478 8200
rect 3424 6860 3476 6866
rect 3424 6802 3476 6808
rect 3436 6225 3464 6802
rect 3422 6216 3478 6225
rect 3422 6151 3478 6160
rect 3330 4856 3386 4865
rect 3330 4791 3386 4800
rect 3344 4690 3372 4791
rect 3332 4684 3384 4690
rect 3332 4626 3384 4632
rect 3252 4134 3372 4162
rect 3240 4072 3292 4078
rect 3240 4014 3292 4020
rect 3148 2848 3200 2854
rect 3148 2790 3200 2796
rect 2872 2644 2924 2650
rect 2872 2586 2924 2592
rect 3252 800 3280 4014
rect 3344 1465 3372 4134
rect 3712 3505 3740 20810
rect 3974 15600 4030 15609
rect 3974 15535 4030 15544
rect 3988 15502 4016 15535
rect 3976 15496 4028 15502
rect 3976 15438 4028 15444
rect 4080 15162 4108 24686
rect 4160 23520 4212 23526
rect 4160 23462 4212 23468
rect 4172 19854 4200 23462
rect 4724 22710 4752 25162
rect 5460 24138 5488 45290
rect 5582 45180 5890 45200
rect 5582 45178 5588 45180
rect 5644 45178 5668 45180
rect 5724 45178 5748 45180
rect 5804 45178 5828 45180
rect 5884 45178 5890 45180
rect 5644 45126 5646 45178
rect 5826 45126 5828 45178
rect 5582 45124 5588 45126
rect 5644 45124 5668 45126
rect 5724 45124 5748 45126
rect 5804 45124 5828 45126
rect 5884 45124 5890 45126
rect 5582 45104 5890 45124
rect 5582 44092 5890 44112
rect 5582 44090 5588 44092
rect 5644 44090 5668 44092
rect 5724 44090 5748 44092
rect 5804 44090 5828 44092
rect 5884 44090 5890 44092
rect 5644 44038 5646 44090
rect 5826 44038 5828 44090
rect 5582 44036 5588 44038
rect 5644 44036 5668 44038
rect 5724 44036 5748 44038
rect 5804 44036 5828 44038
rect 5884 44036 5890 44038
rect 5582 44016 5890 44036
rect 5582 43004 5890 43024
rect 5582 43002 5588 43004
rect 5644 43002 5668 43004
rect 5724 43002 5748 43004
rect 5804 43002 5828 43004
rect 5884 43002 5890 43004
rect 5644 42950 5646 43002
rect 5826 42950 5828 43002
rect 5582 42948 5588 42950
rect 5644 42948 5668 42950
rect 5724 42948 5748 42950
rect 5804 42948 5828 42950
rect 5884 42948 5890 42950
rect 5582 42928 5890 42948
rect 5582 41916 5890 41936
rect 5582 41914 5588 41916
rect 5644 41914 5668 41916
rect 5724 41914 5748 41916
rect 5804 41914 5828 41916
rect 5884 41914 5890 41916
rect 5644 41862 5646 41914
rect 5826 41862 5828 41914
rect 5582 41860 5588 41862
rect 5644 41860 5668 41862
rect 5724 41860 5748 41862
rect 5804 41860 5828 41862
rect 5884 41860 5890 41862
rect 5582 41840 5890 41860
rect 5582 40828 5890 40848
rect 5582 40826 5588 40828
rect 5644 40826 5668 40828
rect 5724 40826 5748 40828
rect 5804 40826 5828 40828
rect 5884 40826 5890 40828
rect 5644 40774 5646 40826
rect 5826 40774 5828 40826
rect 5582 40772 5588 40774
rect 5644 40772 5668 40774
rect 5724 40772 5748 40774
rect 5804 40772 5828 40774
rect 5884 40772 5890 40774
rect 5582 40752 5890 40772
rect 5582 39740 5890 39760
rect 5582 39738 5588 39740
rect 5644 39738 5668 39740
rect 5724 39738 5748 39740
rect 5804 39738 5828 39740
rect 5884 39738 5890 39740
rect 5644 39686 5646 39738
rect 5826 39686 5828 39738
rect 5582 39684 5588 39686
rect 5644 39684 5668 39686
rect 5724 39684 5748 39686
rect 5804 39684 5828 39686
rect 5884 39684 5890 39686
rect 5582 39664 5890 39684
rect 5582 38652 5890 38672
rect 5582 38650 5588 38652
rect 5644 38650 5668 38652
rect 5724 38650 5748 38652
rect 5804 38650 5828 38652
rect 5884 38650 5890 38652
rect 5644 38598 5646 38650
rect 5826 38598 5828 38650
rect 5582 38596 5588 38598
rect 5644 38596 5668 38598
rect 5724 38596 5748 38598
rect 5804 38596 5828 38598
rect 5884 38596 5890 38598
rect 5582 38576 5890 38596
rect 5582 37564 5890 37584
rect 5582 37562 5588 37564
rect 5644 37562 5668 37564
rect 5724 37562 5748 37564
rect 5804 37562 5828 37564
rect 5884 37562 5890 37564
rect 5644 37510 5646 37562
rect 5826 37510 5828 37562
rect 5582 37508 5588 37510
rect 5644 37508 5668 37510
rect 5724 37508 5748 37510
rect 5804 37508 5828 37510
rect 5884 37508 5890 37510
rect 5582 37488 5890 37508
rect 5582 36476 5890 36496
rect 5582 36474 5588 36476
rect 5644 36474 5668 36476
rect 5724 36474 5748 36476
rect 5804 36474 5828 36476
rect 5884 36474 5890 36476
rect 5644 36422 5646 36474
rect 5826 36422 5828 36474
rect 5582 36420 5588 36422
rect 5644 36420 5668 36422
rect 5724 36420 5748 36422
rect 5804 36420 5828 36422
rect 5884 36420 5890 36422
rect 5582 36400 5890 36420
rect 5582 35388 5890 35408
rect 5582 35386 5588 35388
rect 5644 35386 5668 35388
rect 5724 35386 5748 35388
rect 5804 35386 5828 35388
rect 5884 35386 5890 35388
rect 5644 35334 5646 35386
rect 5826 35334 5828 35386
rect 5582 35332 5588 35334
rect 5644 35332 5668 35334
rect 5724 35332 5748 35334
rect 5804 35332 5828 35334
rect 5884 35332 5890 35334
rect 5582 35312 5890 35332
rect 5582 34300 5890 34320
rect 5582 34298 5588 34300
rect 5644 34298 5668 34300
rect 5724 34298 5748 34300
rect 5804 34298 5828 34300
rect 5884 34298 5890 34300
rect 5644 34246 5646 34298
rect 5826 34246 5828 34298
rect 5582 34244 5588 34246
rect 5644 34244 5668 34246
rect 5724 34244 5748 34246
rect 5804 34244 5828 34246
rect 5884 34244 5890 34246
rect 5582 34224 5890 34244
rect 5582 33212 5890 33232
rect 5582 33210 5588 33212
rect 5644 33210 5668 33212
rect 5724 33210 5748 33212
rect 5804 33210 5828 33212
rect 5884 33210 5890 33212
rect 5644 33158 5646 33210
rect 5826 33158 5828 33210
rect 5582 33156 5588 33158
rect 5644 33156 5668 33158
rect 5724 33156 5748 33158
rect 5804 33156 5828 33158
rect 5884 33156 5890 33158
rect 5582 33136 5890 33156
rect 5582 32124 5890 32144
rect 5582 32122 5588 32124
rect 5644 32122 5668 32124
rect 5724 32122 5748 32124
rect 5804 32122 5828 32124
rect 5884 32122 5890 32124
rect 5644 32070 5646 32122
rect 5826 32070 5828 32122
rect 5582 32068 5588 32070
rect 5644 32068 5668 32070
rect 5724 32068 5748 32070
rect 5804 32068 5828 32070
rect 5884 32068 5890 32070
rect 5582 32048 5890 32068
rect 5582 31036 5890 31056
rect 5582 31034 5588 31036
rect 5644 31034 5668 31036
rect 5724 31034 5748 31036
rect 5804 31034 5828 31036
rect 5884 31034 5890 31036
rect 5644 30982 5646 31034
rect 5826 30982 5828 31034
rect 5582 30980 5588 30982
rect 5644 30980 5668 30982
rect 5724 30980 5748 30982
rect 5804 30980 5828 30982
rect 5884 30980 5890 30982
rect 5582 30960 5890 30980
rect 5582 29948 5890 29968
rect 5582 29946 5588 29948
rect 5644 29946 5668 29948
rect 5724 29946 5748 29948
rect 5804 29946 5828 29948
rect 5884 29946 5890 29948
rect 5644 29894 5646 29946
rect 5826 29894 5828 29946
rect 5582 29892 5588 29894
rect 5644 29892 5668 29894
rect 5724 29892 5748 29894
rect 5804 29892 5828 29894
rect 5884 29892 5890 29894
rect 5582 29872 5890 29892
rect 5582 28860 5890 28880
rect 5582 28858 5588 28860
rect 5644 28858 5668 28860
rect 5724 28858 5748 28860
rect 5804 28858 5828 28860
rect 5884 28858 5890 28860
rect 5644 28806 5646 28858
rect 5826 28806 5828 28858
rect 5582 28804 5588 28806
rect 5644 28804 5668 28806
rect 5724 28804 5748 28806
rect 5804 28804 5828 28806
rect 5884 28804 5890 28806
rect 5582 28784 5890 28804
rect 5582 27772 5890 27792
rect 5582 27770 5588 27772
rect 5644 27770 5668 27772
rect 5724 27770 5748 27772
rect 5804 27770 5828 27772
rect 5884 27770 5890 27772
rect 5644 27718 5646 27770
rect 5826 27718 5828 27770
rect 5582 27716 5588 27718
rect 5644 27716 5668 27718
rect 5724 27716 5748 27718
rect 5804 27716 5828 27718
rect 5884 27716 5890 27718
rect 5582 27696 5890 27716
rect 5582 26684 5890 26704
rect 5582 26682 5588 26684
rect 5644 26682 5668 26684
rect 5724 26682 5748 26684
rect 5804 26682 5828 26684
rect 5884 26682 5890 26684
rect 5644 26630 5646 26682
rect 5826 26630 5828 26682
rect 5582 26628 5588 26630
rect 5644 26628 5668 26630
rect 5724 26628 5748 26630
rect 5804 26628 5828 26630
rect 5884 26628 5890 26630
rect 5582 26608 5890 26628
rect 5582 25596 5890 25616
rect 5582 25594 5588 25596
rect 5644 25594 5668 25596
rect 5724 25594 5748 25596
rect 5804 25594 5828 25596
rect 5884 25594 5890 25596
rect 5644 25542 5646 25594
rect 5826 25542 5828 25594
rect 5582 25540 5588 25542
rect 5644 25540 5668 25542
rect 5724 25540 5748 25542
rect 5804 25540 5828 25542
rect 5884 25540 5890 25542
rect 5582 25520 5890 25540
rect 5540 25288 5592 25294
rect 5540 25230 5592 25236
rect 5552 24818 5580 25230
rect 5540 24812 5592 24818
rect 5540 24754 5592 24760
rect 5908 24812 5960 24818
rect 5908 24754 5960 24760
rect 5582 24508 5890 24528
rect 5582 24506 5588 24508
rect 5644 24506 5668 24508
rect 5724 24506 5748 24508
rect 5804 24506 5828 24508
rect 5884 24506 5890 24508
rect 5644 24454 5646 24506
rect 5826 24454 5828 24506
rect 5582 24452 5588 24454
rect 5644 24452 5668 24454
rect 5724 24452 5748 24454
rect 5804 24452 5828 24454
rect 5884 24452 5890 24454
rect 5582 24432 5890 24452
rect 5920 24206 5948 24754
rect 5908 24200 5960 24206
rect 5908 24142 5960 24148
rect 5448 24132 5500 24138
rect 5448 24074 5500 24080
rect 4712 22704 4764 22710
rect 4712 22646 4764 22652
rect 4724 21554 4752 22646
rect 4712 21548 4764 21554
rect 4712 21490 4764 21496
rect 4160 19848 4212 19854
rect 4160 19790 4212 19796
rect 4344 15904 4396 15910
rect 4344 15846 4396 15852
rect 4160 15360 4212 15366
rect 4160 15302 4212 15308
rect 4068 15156 4120 15162
rect 4068 15098 4120 15104
rect 4172 15094 4200 15302
rect 4160 15088 4212 15094
rect 4160 15030 4212 15036
rect 4356 15026 4384 15846
rect 4344 15020 4396 15026
rect 4344 14962 4396 14968
rect 3792 10056 3844 10062
rect 3792 9998 3844 10004
rect 3804 9586 3832 9998
rect 3792 9580 3844 9586
rect 3792 9522 3844 9528
rect 3976 7744 4028 7750
rect 3976 7686 4028 7692
rect 3988 7478 4016 7686
rect 3976 7472 4028 7478
rect 3976 7414 4028 7420
rect 3792 7336 3844 7342
rect 3792 7278 3844 7284
rect 4160 7336 4212 7342
rect 4160 7278 4212 7284
rect 3804 7002 3832 7278
rect 3792 6996 3844 7002
rect 3792 6938 3844 6944
rect 3698 3496 3754 3505
rect 4172 3482 4200 7278
rect 5264 4140 5316 4146
rect 5264 4082 5316 4088
rect 5276 4049 5304 4082
rect 5262 4040 5318 4049
rect 5262 3975 5318 3984
rect 5356 3936 5408 3942
rect 5356 3878 5408 3884
rect 5368 3602 5396 3878
rect 5460 3738 5488 24074
rect 5920 23730 5948 24142
rect 5908 23724 5960 23730
rect 5908 23666 5960 23672
rect 5582 23420 5890 23440
rect 5582 23418 5588 23420
rect 5644 23418 5668 23420
rect 5724 23418 5748 23420
rect 5804 23418 5828 23420
rect 5884 23418 5890 23420
rect 5644 23366 5646 23418
rect 5826 23366 5828 23418
rect 5582 23364 5588 23366
rect 5644 23364 5668 23366
rect 5724 23364 5748 23366
rect 5804 23364 5828 23366
rect 5884 23364 5890 23366
rect 5582 23344 5890 23364
rect 5582 22332 5890 22352
rect 5582 22330 5588 22332
rect 5644 22330 5668 22332
rect 5724 22330 5748 22332
rect 5804 22330 5828 22332
rect 5884 22330 5890 22332
rect 5644 22278 5646 22330
rect 5826 22278 5828 22330
rect 5582 22276 5588 22278
rect 5644 22276 5668 22278
rect 5724 22276 5748 22278
rect 5804 22276 5828 22278
rect 5884 22276 5890 22278
rect 5582 22256 5890 22276
rect 5582 21244 5890 21264
rect 5582 21242 5588 21244
rect 5644 21242 5668 21244
rect 5724 21242 5748 21244
rect 5804 21242 5828 21244
rect 5884 21242 5890 21244
rect 5644 21190 5646 21242
rect 5826 21190 5828 21242
rect 5582 21188 5588 21190
rect 5644 21188 5668 21190
rect 5724 21188 5748 21190
rect 5804 21188 5828 21190
rect 5884 21188 5890 21190
rect 5582 21168 5890 21188
rect 5582 20156 5890 20176
rect 5582 20154 5588 20156
rect 5644 20154 5668 20156
rect 5724 20154 5748 20156
rect 5804 20154 5828 20156
rect 5884 20154 5890 20156
rect 5644 20102 5646 20154
rect 5826 20102 5828 20154
rect 5582 20100 5588 20102
rect 5644 20100 5668 20102
rect 5724 20100 5748 20102
rect 5804 20100 5828 20102
rect 5884 20100 5890 20102
rect 5582 20080 5890 20100
rect 5582 19068 5890 19088
rect 5582 19066 5588 19068
rect 5644 19066 5668 19068
rect 5724 19066 5748 19068
rect 5804 19066 5828 19068
rect 5884 19066 5890 19068
rect 5644 19014 5646 19066
rect 5826 19014 5828 19066
rect 5582 19012 5588 19014
rect 5644 19012 5668 19014
rect 5724 19012 5748 19014
rect 5804 19012 5828 19014
rect 5884 19012 5890 19014
rect 5582 18992 5890 19012
rect 5582 17980 5890 18000
rect 5582 17978 5588 17980
rect 5644 17978 5668 17980
rect 5724 17978 5748 17980
rect 5804 17978 5828 17980
rect 5884 17978 5890 17980
rect 5644 17926 5646 17978
rect 5826 17926 5828 17978
rect 5582 17924 5588 17926
rect 5644 17924 5668 17926
rect 5724 17924 5748 17926
rect 5804 17924 5828 17926
rect 5884 17924 5890 17926
rect 5582 17904 5890 17924
rect 6564 17134 6592 46854
rect 6552 17128 6604 17134
rect 6552 17070 6604 17076
rect 5582 16892 5890 16912
rect 5582 16890 5588 16892
rect 5644 16890 5668 16892
rect 5724 16890 5748 16892
rect 5804 16890 5828 16892
rect 5884 16890 5890 16892
rect 5644 16838 5646 16890
rect 5826 16838 5828 16890
rect 5582 16836 5588 16838
rect 5644 16836 5668 16838
rect 5724 16836 5748 16838
rect 5804 16836 5828 16838
rect 5884 16836 5890 16838
rect 5582 16816 5890 16836
rect 7300 16250 7328 46854
rect 7852 46578 7880 46990
rect 7840 46572 7892 46578
rect 7840 46514 7892 46520
rect 8404 46510 8432 49200
rect 8024 46504 8076 46510
rect 8024 46446 8076 46452
rect 8392 46504 8444 46510
rect 8392 46446 8444 46452
rect 8036 46170 8064 46446
rect 9588 46368 9640 46374
rect 9588 46310 9640 46316
rect 8024 46164 8076 46170
rect 8024 46106 8076 46112
rect 9600 46034 9628 46310
rect 10152 46034 10180 49286
rect 10294 49200 10406 49286
rect 10938 49200 11050 50000
rect 11582 49200 11694 50000
rect 12226 49200 12338 50000
rect 12870 49200 12982 50000
rect 13514 49200 13626 50000
rect 14802 49200 14914 50000
rect 15446 49200 15558 50000
rect 16090 49200 16202 50000
rect 16734 49200 16846 50000
rect 17378 49200 17490 50000
rect 18022 49200 18134 50000
rect 18666 49200 18778 50000
rect 19954 49200 20066 50000
rect 20598 49200 20710 50000
rect 21242 49200 21354 50000
rect 21886 49200 21998 50000
rect 22530 49200 22642 50000
rect 23174 49200 23286 50000
rect 23818 49200 23930 50000
rect 25106 49200 25218 50000
rect 25750 49200 25862 50000
rect 26394 49200 26506 50000
rect 27038 49200 27150 50000
rect 27682 49314 27794 50000
rect 27682 49286 28028 49314
rect 27682 49200 27794 49286
rect 10214 46812 10522 46832
rect 10214 46810 10220 46812
rect 10276 46810 10300 46812
rect 10356 46810 10380 46812
rect 10436 46810 10460 46812
rect 10516 46810 10522 46812
rect 10276 46758 10278 46810
rect 10458 46758 10460 46810
rect 10214 46756 10220 46758
rect 10276 46756 10300 46758
rect 10356 46756 10380 46758
rect 10436 46756 10460 46758
rect 10516 46756 10522 46758
rect 10214 46736 10522 46756
rect 10980 46374 11008 49200
rect 11624 46918 11652 49200
rect 11612 46912 11664 46918
rect 11612 46854 11664 46860
rect 12532 46912 12584 46918
rect 12532 46854 12584 46860
rect 11704 46504 11756 46510
rect 11704 46446 11756 46452
rect 10968 46368 11020 46374
rect 10968 46310 11020 46316
rect 9588 46028 9640 46034
rect 9588 45970 9640 45976
rect 10140 46028 10192 46034
rect 10140 45970 10192 45976
rect 9864 45892 9916 45898
rect 9864 45834 9916 45840
rect 9876 45626 9904 45834
rect 10214 45724 10522 45744
rect 10214 45722 10220 45724
rect 10276 45722 10300 45724
rect 10356 45722 10380 45724
rect 10436 45722 10460 45724
rect 10516 45722 10522 45724
rect 10276 45670 10278 45722
rect 10458 45670 10460 45722
rect 10214 45668 10220 45670
rect 10276 45668 10300 45670
rect 10356 45668 10380 45670
rect 10436 45668 10460 45670
rect 10516 45668 10522 45670
rect 10214 45648 10522 45668
rect 9864 45620 9916 45626
rect 9864 45562 9916 45568
rect 11716 45558 11744 46446
rect 11704 45552 11756 45558
rect 11704 45494 11756 45500
rect 9956 45484 10008 45490
rect 9956 45426 10008 45432
rect 9968 41614 9996 45426
rect 12544 44946 12572 46854
rect 13452 46504 13504 46510
rect 13452 46446 13504 46452
rect 13464 46170 13492 46446
rect 13556 46442 13584 49200
rect 14844 47546 14872 49200
rect 14752 47518 14872 47546
rect 13820 47048 13872 47054
rect 13820 46990 13872 46996
rect 13832 46578 13860 46990
rect 13820 46572 13872 46578
rect 13820 46514 13872 46520
rect 13544 46436 13596 46442
rect 13544 46378 13596 46384
rect 13452 46164 13504 46170
rect 13452 46106 13504 46112
rect 14280 45960 14332 45966
rect 14280 45902 14332 45908
rect 14292 45422 14320 45902
rect 14752 45898 14780 47518
rect 14846 47356 15154 47376
rect 14846 47354 14852 47356
rect 14908 47354 14932 47356
rect 14988 47354 15012 47356
rect 15068 47354 15092 47356
rect 15148 47354 15154 47356
rect 14908 47302 14910 47354
rect 15090 47302 15092 47354
rect 14846 47300 14852 47302
rect 14908 47300 14932 47302
rect 14988 47300 15012 47302
rect 15068 47300 15092 47302
rect 15148 47300 15154 47302
rect 14846 47280 15154 47300
rect 16672 47048 16724 47054
rect 16672 46990 16724 46996
rect 16684 46578 16712 46990
rect 16672 46572 16724 46578
rect 16672 46514 16724 46520
rect 16776 46442 16804 49200
rect 18144 47048 18196 47054
rect 18144 46990 18196 46996
rect 16856 46504 16908 46510
rect 16856 46446 16908 46452
rect 16764 46436 16816 46442
rect 16764 46378 16816 46384
rect 14846 46268 15154 46288
rect 14846 46266 14852 46268
rect 14908 46266 14932 46268
rect 14988 46266 15012 46268
rect 15068 46266 15092 46268
rect 15148 46266 15154 46268
rect 14908 46214 14910 46266
rect 15090 46214 15092 46266
rect 14846 46212 14852 46214
rect 14908 46212 14932 46214
rect 14988 46212 15012 46214
rect 15068 46212 15092 46214
rect 15148 46212 15154 46214
rect 14846 46192 15154 46212
rect 16868 46170 16896 46446
rect 17592 46368 17644 46374
rect 17592 46310 17644 46316
rect 16856 46164 16908 46170
rect 16856 46106 16908 46112
rect 14464 45892 14516 45898
rect 14464 45834 14516 45840
rect 14740 45892 14792 45898
rect 14740 45834 14792 45840
rect 14476 45626 14504 45834
rect 14464 45620 14516 45626
rect 14464 45562 14516 45568
rect 14372 45484 14424 45490
rect 14372 45426 14424 45432
rect 14280 45416 14332 45422
rect 14280 45358 14332 45364
rect 14384 45014 14412 45426
rect 14846 45180 15154 45200
rect 14846 45178 14852 45180
rect 14908 45178 14932 45180
rect 14988 45178 15012 45180
rect 15068 45178 15092 45180
rect 15148 45178 15154 45180
rect 14908 45126 14910 45178
rect 15090 45126 15092 45178
rect 14846 45124 14852 45126
rect 14908 45124 14932 45126
rect 14988 45124 15012 45126
rect 15068 45124 15092 45126
rect 15148 45124 15154 45126
rect 14846 45104 15154 45124
rect 14372 45008 14424 45014
rect 14372 44950 14424 44956
rect 12532 44940 12584 44946
rect 12532 44882 12584 44888
rect 11612 44804 11664 44810
rect 11612 44746 11664 44752
rect 10214 44636 10522 44656
rect 10214 44634 10220 44636
rect 10276 44634 10300 44636
rect 10356 44634 10380 44636
rect 10436 44634 10460 44636
rect 10516 44634 10522 44636
rect 10276 44582 10278 44634
rect 10458 44582 10460 44634
rect 10214 44580 10220 44582
rect 10276 44580 10300 44582
rect 10356 44580 10380 44582
rect 10436 44580 10460 44582
rect 10516 44580 10522 44582
rect 10214 44560 10522 44580
rect 11624 44538 11652 44746
rect 11612 44532 11664 44538
rect 11612 44474 11664 44480
rect 11704 44396 11756 44402
rect 11704 44338 11756 44344
rect 10214 43548 10522 43568
rect 10214 43546 10220 43548
rect 10276 43546 10300 43548
rect 10356 43546 10380 43548
rect 10436 43546 10460 43548
rect 10516 43546 10522 43548
rect 10276 43494 10278 43546
rect 10458 43494 10460 43546
rect 10214 43492 10220 43494
rect 10276 43492 10300 43494
rect 10356 43492 10380 43494
rect 10436 43492 10460 43494
rect 10516 43492 10522 43494
rect 10214 43472 10522 43492
rect 10214 42460 10522 42480
rect 10214 42458 10220 42460
rect 10276 42458 10300 42460
rect 10356 42458 10380 42460
rect 10436 42458 10460 42460
rect 10516 42458 10522 42460
rect 10276 42406 10278 42458
rect 10458 42406 10460 42458
rect 10214 42404 10220 42406
rect 10276 42404 10300 42406
rect 10356 42404 10380 42406
rect 10436 42404 10460 42406
rect 10516 42404 10522 42406
rect 10214 42384 10522 42404
rect 9956 41608 10008 41614
rect 9956 41550 10008 41556
rect 10600 41608 10652 41614
rect 10600 41550 10652 41556
rect 10214 41372 10522 41392
rect 10214 41370 10220 41372
rect 10276 41370 10300 41372
rect 10356 41370 10380 41372
rect 10436 41370 10460 41372
rect 10516 41370 10522 41372
rect 10276 41318 10278 41370
rect 10458 41318 10460 41370
rect 10214 41316 10220 41318
rect 10276 41316 10300 41318
rect 10356 41316 10380 41318
rect 10436 41316 10460 41318
rect 10516 41316 10522 41318
rect 10214 41296 10522 41316
rect 10214 40284 10522 40304
rect 10214 40282 10220 40284
rect 10276 40282 10300 40284
rect 10356 40282 10380 40284
rect 10436 40282 10460 40284
rect 10516 40282 10522 40284
rect 10276 40230 10278 40282
rect 10458 40230 10460 40282
rect 10214 40228 10220 40230
rect 10276 40228 10300 40230
rect 10356 40228 10380 40230
rect 10436 40228 10460 40230
rect 10516 40228 10522 40230
rect 10214 40208 10522 40228
rect 10214 39196 10522 39216
rect 10214 39194 10220 39196
rect 10276 39194 10300 39196
rect 10356 39194 10380 39196
rect 10436 39194 10460 39196
rect 10516 39194 10522 39196
rect 10276 39142 10278 39194
rect 10458 39142 10460 39194
rect 10214 39140 10220 39142
rect 10276 39140 10300 39142
rect 10356 39140 10380 39142
rect 10436 39140 10460 39142
rect 10516 39140 10522 39142
rect 10214 39120 10522 39140
rect 10214 38108 10522 38128
rect 10214 38106 10220 38108
rect 10276 38106 10300 38108
rect 10356 38106 10380 38108
rect 10436 38106 10460 38108
rect 10516 38106 10522 38108
rect 10276 38054 10278 38106
rect 10458 38054 10460 38106
rect 10214 38052 10220 38054
rect 10276 38052 10300 38054
rect 10356 38052 10380 38054
rect 10436 38052 10460 38054
rect 10516 38052 10522 38054
rect 10214 38032 10522 38052
rect 10214 37020 10522 37040
rect 10214 37018 10220 37020
rect 10276 37018 10300 37020
rect 10356 37018 10380 37020
rect 10436 37018 10460 37020
rect 10516 37018 10522 37020
rect 10276 36966 10278 37018
rect 10458 36966 10460 37018
rect 10214 36964 10220 36966
rect 10276 36964 10300 36966
rect 10356 36964 10380 36966
rect 10436 36964 10460 36966
rect 10516 36964 10522 36966
rect 10214 36944 10522 36964
rect 10214 35932 10522 35952
rect 10214 35930 10220 35932
rect 10276 35930 10300 35932
rect 10356 35930 10380 35932
rect 10436 35930 10460 35932
rect 10516 35930 10522 35932
rect 10276 35878 10278 35930
rect 10458 35878 10460 35930
rect 10214 35876 10220 35878
rect 10276 35876 10300 35878
rect 10356 35876 10380 35878
rect 10436 35876 10460 35878
rect 10516 35876 10522 35878
rect 10214 35856 10522 35876
rect 10612 35193 10640 41550
rect 11716 35494 11744 44338
rect 14846 44092 15154 44112
rect 14846 44090 14852 44092
rect 14908 44090 14932 44092
rect 14988 44090 15012 44092
rect 15068 44090 15092 44092
rect 15148 44090 15154 44092
rect 14908 44038 14910 44090
rect 15090 44038 15092 44090
rect 14846 44036 14852 44038
rect 14908 44036 14932 44038
rect 14988 44036 15012 44038
rect 15068 44036 15092 44038
rect 15148 44036 15154 44038
rect 14846 44016 15154 44036
rect 14846 43004 15154 43024
rect 14846 43002 14852 43004
rect 14908 43002 14932 43004
rect 14988 43002 15012 43004
rect 15068 43002 15092 43004
rect 15148 43002 15154 43004
rect 14908 42950 14910 43002
rect 15090 42950 15092 43002
rect 14846 42948 14852 42950
rect 14908 42948 14932 42950
rect 14988 42948 15012 42950
rect 15068 42948 15092 42950
rect 15148 42948 15154 42950
rect 14846 42928 15154 42948
rect 14846 41916 15154 41936
rect 14846 41914 14852 41916
rect 14908 41914 14932 41916
rect 14988 41914 15012 41916
rect 15068 41914 15092 41916
rect 15148 41914 15154 41916
rect 14908 41862 14910 41914
rect 15090 41862 15092 41914
rect 14846 41860 14852 41862
rect 14908 41860 14932 41862
rect 14988 41860 15012 41862
rect 15068 41860 15092 41862
rect 15148 41860 15154 41862
rect 14846 41840 15154 41860
rect 14846 40828 15154 40848
rect 14846 40826 14852 40828
rect 14908 40826 14932 40828
rect 14988 40826 15012 40828
rect 15068 40826 15092 40828
rect 15148 40826 15154 40828
rect 14908 40774 14910 40826
rect 15090 40774 15092 40826
rect 14846 40772 14852 40774
rect 14908 40772 14932 40774
rect 14988 40772 15012 40774
rect 15068 40772 15092 40774
rect 15148 40772 15154 40774
rect 14846 40752 15154 40772
rect 14846 39740 15154 39760
rect 14846 39738 14852 39740
rect 14908 39738 14932 39740
rect 14988 39738 15012 39740
rect 15068 39738 15092 39740
rect 15148 39738 15154 39740
rect 14908 39686 14910 39738
rect 15090 39686 15092 39738
rect 14846 39684 14852 39686
rect 14908 39684 14932 39686
rect 14988 39684 15012 39686
rect 15068 39684 15092 39686
rect 15148 39684 15154 39686
rect 14846 39664 15154 39684
rect 14846 38652 15154 38672
rect 14846 38650 14852 38652
rect 14908 38650 14932 38652
rect 14988 38650 15012 38652
rect 15068 38650 15092 38652
rect 15148 38650 15154 38652
rect 14908 38598 14910 38650
rect 15090 38598 15092 38650
rect 14846 38596 14852 38598
rect 14908 38596 14932 38598
rect 14988 38596 15012 38598
rect 15068 38596 15092 38598
rect 15148 38596 15154 38598
rect 14846 38576 15154 38596
rect 14846 37564 15154 37584
rect 14846 37562 14852 37564
rect 14908 37562 14932 37564
rect 14988 37562 15012 37564
rect 15068 37562 15092 37564
rect 15148 37562 15154 37564
rect 14908 37510 14910 37562
rect 15090 37510 15092 37562
rect 14846 37508 14852 37510
rect 14908 37508 14932 37510
rect 14988 37508 15012 37510
rect 15068 37508 15092 37510
rect 15148 37508 15154 37510
rect 14846 37488 15154 37508
rect 16948 36576 17000 36582
rect 16948 36518 17000 36524
rect 14846 36476 15154 36496
rect 14846 36474 14852 36476
rect 14908 36474 14932 36476
rect 14988 36474 15012 36476
rect 15068 36474 15092 36476
rect 15148 36474 15154 36476
rect 14908 36422 14910 36474
rect 15090 36422 15092 36474
rect 14846 36420 14852 36422
rect 14908 36420 14932 36422
rect 14988 36420 15012 36422
rect 15068 36420 15092 36422
rect 15148 36420 15154 36422
rect 14846 36400 15154 36420
rect 16960 35766 16988 36518
rect 16948 35760 17000 35766
rect 16948 35702 17000 35708
rect 11704 35488 11756 35494
rect 11704 35430 11756 35436
rect 14846 35388 15154 35408
rect 14846 35386 14852 35388
rect 14908 35386 14932 35388
rect 14988 35386 15012 35388
rect 15068 35386 15092 35388
rect 15148 35386 15154 35388
rect 14908 35334 14910 35386
rect 15090 35334 15092 35386
rect 14846 35332 14852 35334
rect 14908 35332 14932 35334
rect 14988 35332 15012 35334
rect 15068 35332 15092 35334
rect 15148 35332 15154 35334
rect 14846 35312 15154 35332
rect 10598 35184 10654 35193
rect 10598 35119 10654 35128
rect 10214 34844 10522 34864
rect 10214 34842 10220 34844
rect 10276 34842 10300 34844
rect 10356 34842 10380 34844
rect 10436 34842 10460 34844
rect 10516 34842 10522 34844
rect 10276 34790 10278 34842
rect 10458 34790 10460 34842
rect 10214 34788 10220 34790
rect 10276 34788 10300 34790
rect 10356 34788 10380 34790
rect 10436 34788 10460 34790
rect 10516 34788 10522 34790
rect 10214 34768 10522 34788
rect 14846 34300 15154 34320
rect 14846 34298 14852 34300
rect 14908 34298 14932 34300
rect 14988 34298 15012 34300
rect 15068 34298 15092 34300
rect 15148 34298 15154 34300
rect 14908 34246 14910 34298
rect 15090 34246 15092 34298
rect 14846 34244 14852 34246
rect 14908 34244 14932 34246
rect 14988 34244 15012 34246
rect 15068 34244 15092 34246
rect 15148 34244 15154 34246
rect 14846 34224 15154 34244
rect 10214 33756 10522 33776
rect 10214 33754 10220 33756
rect 10276 33754 10300 33756
rect 10356 33754 10380 33756
rect 10436 33754 10460 33756
rect 10516 33754 10522 33756
rect 10276 33702 10278 33754
rect 10458 33702 10460 33754
rect 10214 33700 10220 33702
rect 10276 33700 10300 33702
rect 10356 33700 10380 33702
rect 10436 33700 10460 33702
rect 10516 33700 10522 33702
rect 10214 33680 10522 33700
rect 14846 33212 15154 33232
rect 14846 33210 14852 33212
rect 14908 33210 14932 33212
rect 14988 33210 15012 33212
rect 15068 33210 15092 33212
rect 15148 33210 15154 33212
rect 14908 33158 14910 33210
rect 15090 33158 15092 33210
rect 14846 33156 14852 33158
rect 14908 33156 14932 33158
rect 14988 33156 15012 33158
rect 15068 33156 15092 33158
rect 15148 33156 15154 33158
rect 14846 33136 15154 33156
rect 10214 32668 10522 32688
rect 10214 32666 10220 32668
rect 10276 32666 10300 32668
rect 10356 32666 10380 32668
rect 10436 32666 10460 32668
rect 10516 32666 10522 32668
rect 10276 32614 10278 32666
rect 10458 32614 10460 32666
rect 10214 32612 10220 32614
rect 10276 32612 10300 32614
rect 10356 32612 10380 32614
rect 10436 32612 10460 32614
rect 10516 32612 10522 32614
rect 10214 32592 10522 32612
rect 16764 32428 16816 32434
rect 16764 32370 16816 32376
rect 14846 32124 15154 32144
rect 14846 32122 14852 32124
rect 14908 32122 14932 32124
rect 14988 32122 15012 32124
rect 15068 32122 15092 32124
rect 15148 32122 15154 32124
rect 14908 32070 14910 32122
rect 15090 32070 15092 32122
rect 14846 32068 14852 32070
rect 14908 32068 14932 32070
rect 14988 32068 15012 32070
rect 15068 32068 15092 32070
rect 15148 32068 15154 32070
rect 14846 32048 15154 32068
rect 16776 31958 16804 32370
rect 16764 31952 16816 31958
rect 16764 31894 16816 31900
rect 17604 31890 17632 46310
rect 18052 45824 18104 45830
rect 18052 45766 18104 45772
rect 18064 45626 18092 45766
rect 18052 45620 18104 45626
rect 18052 45562 18104 45568
rect 18156 45490 18184 46990
rect 18236 45960 18288 45966
rect 18236 45902 18288 45908
rect 18144 45484 18196 45490
rect 18144 45426 18196 45432
rect 17960 36780 18012 36786
rect 17960 36722 18012 36728
rect 17972 36174 18000 36722
rect 17960 36168 18012 36174
rect 17960 36110 18012 36116
rect 17972 35698 18000 36110
rect 18248 35766 18276 45902
rect 18328 45824 18380 45830
rect 18328 45766 18380 45772
rect 18340 45558 18368 45766
rect 18328 45552 18380 45558
rect 18328 45494 18380 45500
rect 18708 45422 18736 49200
rect 19340 47048 19392 47054
rect 19340 46990 19392 46996
rect 19352 46578 19380 46990
rect 19478 46812 19786 46832
rect 19478 46810 19484 46812
rect 19540 46810 19564 46812
rect 19620 46810 19644 46812
rect 19700 46810 19724 46812
rect 19780 46810 19786 46812
rect 19540 46758 19542 46810
rect 19722 46758 19724 46810
rect 19478 46756 19484 46758
rect 19540 46756 19564 46758
rect 19620 46756 19644 46758
rect 19700 46756 19724 46758
rect 19780 46756 19786 46758
rect 19478 46736 19786 46756
rect 19340 46572 19392 46578
rect 19340 46514 19392 46520
rect 19996 46510 20024 49200
rect 19984 46504 20036 46510
rect 19984 46446 20036 46452
rect 19340 46436 19392 46442
rect 19340 46378 19392 46384
rect 18696 45416 18748 45422
rect 18696 45358 18748 45364
rect 19352 45082 19380 46378
rect 21284 46034 21312 49200
rect 21916 47048 21968 47054
rect 21916 46990 21968 46996
rect 20168 46028 20220 46034
rect 20168 45970 20220 45976
rect 21272 46028 21324 46034
rect 21272 45970 21324 45976
rect 19892 45892 19944 45898
rect 19892 45834 19944 45840
rect 19478 45724 19786 45744
rect 19478 45722 19484 45724
rect 19540 45722 19564 45724
rect 19620 45722 19644 45724
rect 19700 45722 19724 45724
rect 19780 45722 19786 45724
rect 19540 45670 19542 45722
rect 19722 45670 19724 45722
rect 19478 45668 19484 45670
rect 19540 45668 19564 45670
rect 19620 45668 19644 45670
rect 19700 45668 19724 45670
rect 19780 45668 19786 45670
rect 19478 45648 19786 45668
rect 19904 45626 19932 45834
rect 19892 45620 19944 45626
rect 19892 45562 19944 45568
rect 19524 45552 19576 45558
rect 19524 45494 19576 45500
rect 19340 45076 19392 45082
rect 19340 45018 19392 45024
rect 19536 44878 19564 45494
rect 20180 45082 20208 45970
rect 20444 45484 20496 45490
rect 20444 45426 20496 45432
rect 20168 45076 20220 45082
rect 20168 45018 20220 45024
rect 19340 44872 19392 44878
rect 19340 44814 19392 44820
rect 19524 44872 19576 44878
rect 19524 44814 19576 44820
rect 19352 40118 19380 44814
rect 19478 44636 19786 44656
rect 19478 44634 19484 44636
rect 19540 44634 19564 44636
rect 19620 44634 19644 44636
rect 19700 44634 19724 44636
rect 19780 44634 19786 44636
rect 19540 44582 19542 44634
rect 19722 44582 19724 44634
rect 19478 44580 19484 44582
rect 19540 44580 19564 44582
rect 19620 44580 19644 44582
rect 19700 44580 19724 44582
rect 19780 44580 19786 44582
rect 19478 44560 19786 44580
rect 19478 43548 19786 43568
rect 19478 43546 19484 43548
rect 19540 43546 19564 43548
rect 19620 43546 19644 43548
rect 19700 43546 19724 43548
rect 19780 43546 19786 43548
rect 19540 43494 19542 43546
rect 19722 43494 19724 43546
rect 19478 43492 19484 43494
rect 19540 43492 19564 43494
rect 19620 43492 19644 43494
rect 19700 43492 19724 43494
rect 19780 43492 19786 43494
rect 19478 43472 19786 43492
rect 19478 42460 19786 42480
rect 19478 42458 19484 42460
rect 19540 42458 19564 42460
rect 19620 42458 19644 42460
rect 19700 42458 19724 42460
rect 19780 42458 19786 42460
rect 19540 42406 19542 42458
rect 19722 42406 19724 42458
rect 19478 42404 19484 42406
rect 19540 42404 19564 42406
rect 19620 42404 19644 42406
rect 19700 42404 19724 42406
rect 19780 42404 19786 42406
rect 19478 42384 19786 42404
rect 19478 41372 19786 41392
rect 19478 41370 19484 41372
rect 19540 41370 19564 41372
rect 19620 41370 19644 41372
rect 19700 41370 19724 41372
rect 19780 41370 19786 41372
rect 19540 41318 19542 41370
rect 19722 41318 19724 41370
rect 19478 41316 19484 41318
rect 19540 41316 19564 41318
rect 19620 41316 19644 41318
rect 19700 41316 19724 41318
rect 19780 41316 19786 41318
rect 19478 41296 19786 41316
rect 19478 40284 19786 40304
rect 19478 40282 19484 40284
rect 19540 40282 19564 40284
rect 19620 40282 19644 40284
rect 19700 40282 19724 40284
rect 19780 40282 19786 40284
rect 19540 40230 19542 40282
rect 19722 40230 19724 40282
rect 19478 40228 19484 40230
rect 19540 40228 19564 40230
rect 19620 40228 19644 40230
rect 19700 40228 19724 40230
rect 19780 40228 19786 40230
rect 19478 40208 19786 40228
rect 19340 40112 19392 40118
rect 19340 40054 19392 40060
rect 19352 39114 19380 40054
rect 19478 39196 19786 39216
rect 19478 39194 19484 39196
rect 19540 39194 19564 39196
rect 19620 39194 19644 39196
rect 19700 39194 19724 39196
rect 19780 39194 19786 39196
rect 19540 39142 19542 39194
rect 19722 39142 19724 39194
rect 19478 39140 19484 39142
rect 19540 39140 19564 39142
rect 19620 39140 19644 39142
rect 19700 39140 19724 39142
rect 19780 39140 19786 39142
rect 19478 39120 19786 39140
rect 19260 39086 19380 39114
rect 18788 38344 18840 38350
rect 18788 38286 18840 38292
rect 18420 36712 18472 36718
rect 18420 36654 18472 36660
rect 18328 36100 18380 36106
rect 18328 36042 18380 36048
rect 18236 35760 18288 35766
rect 18236 35702 18288 35708
rect 17960 35692 18012 35698
rect 17960 35634 18012 35640
rect 17972 35086 18000 35634
rect 18340 35578 18368 36042
rect 18248 35550 18368 35578
rect 17960 35080 18012 35086
rect 17960 35022 18012 35028
rect 17972 34610 18000 35022
rect 17960 34604 18012 34610
rect 17960 34546 18012 34552
rect 17684 32224 17736 32230
rect 17684 32166 17736 32172
rect 17592 31884 17644 31890
rect 17592 31826 17644 31832
rect 16856 31816 16908 31822
rect 16856 31758 16908 31764
rect 10214 31580 10522 31600
rect 10214 31578 10220 31580
rect 10276 31578 10300 31580
rect 10356 31578 10380 31580
rect 10436 31578 10460 31580
rect 10516 31578 10522 31580
rect 10276 31526 10278 31578
rect 10458 31526 10460 31578
rect 10214 31524 10220 31526
rect 10276 31524 10300 31526
rect 10356 31524 10380 31526
rect 10436 31524 10460 31526
rect 10516 31524 10522 31526
rect 10214 31504 10522 31524
rect 16868 31482 16896 31758
rect 17696 31754 17724 32166
rect 17868 31884 17920 31890
rect 17868 31826 17920 31832
rect 17604 31726 17724 31754
rect 17604 31686 17632 31726
rect 17132 31680 17184 31686
rect 17132 31622 17184 31628
rect 17592 31680 17644 31686
rect 17592 31622 17644 31628
rect 16856 31476 16908 31482
rect 16856 31418 16908 31424
rect 17144 31414 17172 31622
rect 17132 31408 17184 31414
rect 17132 31350 17184 31356
rect 17224 31272 17276 31278
rect 17224 31214 17276 31220
rect 14846 31036 15154 31056
rect 14846 31034 14852 31036
rect 14908 31034 14932 31036
rect 14988 31034 15012 31036
rect 15068 31034 15092 31036
rect 15148 31034 15154 31036
rect 14908 30982 14910 31034
rect 15090 30982 15092 31034
rect 14846 30980 14852 30982
rect 14908 30980 14932 30982
rect 14988 30980 15012 30982
rect 15068 30980 15092 30982
rect 15148 30980 15154 30982
rect 14846 30960 15154 30980
rect 17236 30734 17264 31214
rect 14372 30728 14424 30734
rect 14372 30670 14424 30676
rect 17224 30728 17276 30734
rect 17224 30670 17276 30676
rect 10214 30492 10522 30512
rect 10214 30490 10220 30492
rect 10276 30490 10300 30492
rect 10356 30490 10380 30492
rect 10436 30490 10460 30492
rect 10516 30490 10522 30492
rect 10276 30438 10278 30490
rect 10458 30438 10460 30490
rect 10214 30436 10220 30438
rect 10276 30436 10300 30438
rect 10356 30436 10380 30438
rect 10436 30436 10460 30438
rect 10516 30436 10522 30438
rect 10214 30416 10522 30436
rect 14004 30184 14056 30190
rect 14004 30126 14056 30132
rect 14016 29578 14044 30126
rect 14004 29572 14056 29578
rect 14004 29514 14056 29520
rect 10214 29404 10522 29424
rect 10214 29402 10220 29404
rect 10276 29402 10300 29404
rect 10356 29402 10380 29404
rect 10436 29402 10460 29404
rect 10516 29402 10522 29404
rect 10276 29350 10278 29402
rect 10458 29350 10460 29402
rect 10214 29348 10220 29350
rect 10276 29348 10300 29350
rect 10356 29348 10380 29350
rect 10436 29348 10460 29350
rect 10516 29348 10522 29350
rect 10214 29328 10522 29348
rect 13360 29028 13412 29034
rect 13360 28970 13412 28976
rect 10214 28316 10522 28336
rect 10214 28314 10220 28316
rect 10276 28314 10300 28316
rect 10356 28314 10380 28316
rect 10436 28314 10460 28316
rect 10516 28314 10522 28316
rect 10276 28262 10278 28314
rect 10458 28262 10460 28314
rect 10214 28260 10220 28262
rect 10276 28260 10300 28262
rect 10356 28260 10380 28262
rect 10436 28260 10460 28262
rect 10516 28260 10522 28262
rect 10214 28240 10522 28260
rect 10214 27228 10522 27248
rect 10214 27226 10220 27228
rect 10276 27226 10300 27228
rect 10356 27226 10380 27228
rect 10436 27226 10460 27228
rect 10516 27226 10522 27228
rect 10276 27174 10278 27226
rect 10458 27174 10460 27226
rect 10214 27172 10220 27174
rect 10276 27172 10300 27174
rect 10356 27172 10380 27174
rect 10436 27172 10460 27174
rect 10516 27172 10522 27174
rect 10214 27152 10522 27172
rect 10214 26140 10522 26160
rect 10214 26138 10220 26140
rect 10276 26138 10300 26140
rect 10356 26138 10380 26140
rect 10436 26138 10460 26140
rect 10516 26138 10522 26140
rect 10276 26086 10278 26138
rect 10458 26086 10460 26138
rect 10214 26084 10220 26086
rect 10276 26084 10300 26086
rect 10356 26084 10380 26086
rect 10436 26084 10460 26086
rect 10516 26084 10522 26086
rect 10214 26064 10522 26084
rect 12532 25900 12584 25906
rect 12532 25842 12584 25848
rect 12716 25900 12768 25906
rect 12716 25842 12768 25848
rect 12164 25152 12216 25158
rect 12164 25094 12216 25100
rect 10214 25052 10522 25072
rect 10214 25050 10220 25052
rect 10276 25050 10300 25052
rect 10356 25050 10380 25052
rect 10436 25050 10460 25052
rect 10516 25050 10522 25052
rect 10276 24998 10278 25050
rect 10458 24998 10460 25050
rect 10214 24996 10220 24998
rect 10276 24996 10300 24998
rect 10356 24996 10380 24998
rect 10436 24996 10460 24998
rect 10516 24996 10522 24998
rect 10214 24976 10522 24996
rect 12176 24886 12204 25094
rect 12544 24954 12572 25842
rect 12532 24948 12584 24954
rect 12532 24890 12584 24896
rect 12164 24880 12216 24886
rect 12164 24822 12216 24828
rect 12440 24064 12492 24070
rect 12440 24006 12492 24012
rect 10214 23964 10522 23984
rect 10214 23962 10220 23964
rect 10276 23962 10300 23964
rect 10356 23962 10380 23964
rect 10436 23962 10460 23964
rect 10516 23962 10522 23964
rect 10276 23910 10278 23962
rect 10458 23910 10460 23962
rect 10214 23908 10220 23910
rect 10276 23908 10300 23910
rect 10356 23908 10380 23910
rect 10436 23908 10460 23910
rect 10516 23908 10522 23910
rect 10214 23888 10522 23908
rect 9496 23656 9548 23662
rect 9496 23598 9548 23604
rect 7288 16244 7340 16250
rect 7288 16186 7340 16192
rect 5582 15804 5890 15824
rect 5582 15802 5588 15804
rect 5644 15802 5668 15804
rect 5724 15802 5748 15804
rect 5804 15802 5828 15804
rect 5884 15802 5890 15804
rect 5644 15750 5646 15802
rect 5826 15750 5828 15802
rect 5582 15748 5588 15750
rect 5644 15748 5668 15750
rect 5724 15748 5748 15750
rect 5804 15748 5828 15750
rect 5884 15748 5890 15750
rect 5582 15728 5890 15748
rect 5582 14716 5890 14736
rect 5582 14714 5588 14716
rect 5644 14714 5668 14716
rect 5724 14714 5748 14716
rect 5804 14714 5828 14716
rect 5884 14714 5890 14716
rect 5644 14662 5646 14714
rect 5826 14662 5828 14714
rect 5582 14660 5588 14662
rect 5644 14660 5668 14662
rect 5724 14660 5748 14662
rect 5804 14660 5828 14662
rect 5884 14660 5890 14662
rect 5582 14640 5890 14660
rect 5582 13628 5890 13648
rect 5582 13626 5588 13628
rect 5644 13626 5668 13628
rect 5724 13626 5748 13628
rect 5804 13626 5828 13628
rect 5884 13626 5890 13628
rect 5644 13574 5646 13626
rect 5826 13574 5828 13626
rect 5582 13572 5588 13574
rect 5644 13572 5668 13574
rect 5724 13572 5748 13574
rect 5804 13572 5828 13574
rect 5884 13572 5890 13574
rect 5582 13552 5890 13572
rect 5582 12540 5890 12560
rect 5582 12538 5588 12540
rect 5644 12538 5668 12540
rect 5724 12538 5748 12540
rect 5804 12538 5828 12540
rect 5884 12538 5890 12540
rect 5644 12486 5646 12538
rect 5826 12486 5828 12538
rect 5582 12484 5588 12486
rect 5644 12484 5668 12486
rect 5724 12484 5748 12486
rect 5804 12484 5828 12486
rect 5884 12484 5890 12486
rect 5582 12464 5890 12484
rect 5582 11452 5890 11472
rect 5582 11450 5588 11452
rect 5644 11450 5668 11452
rect 5724 11450 5748 11452
rect 5804 11450 5828 11452
rect 5884 11450 5890 11452
rect 5644 11398 5646 11450
rect 5826 11398 5828 11450
rect 5582 11396 5588 11398
rect 5644 11396 5668 11398
rect 5724 11396 5748 11398
rect 5804 11396 5828 11398
rect 5884 11396 5890 11398
rect 5582 11376 5890 11396
rect 5582 10364 5890 10384
rect 5582 10362 5588 10364
rect 5644 10362 5668 10364
rect 5724 10362 5748 10364
rect 5804 10362 5828 10364
rect 5884 10362 5890 10364
rect 5644 10310 5646 10362
rect 5826 10310 5828 10362
rect 5582 10308 5588 10310
rect 5644 10308 5668 10310
rect 5724 10308 5748 10310
rect 5804 10308 5828 10310
rect 5884 10308 5890 10310
rect 5582 10288 5890 10308
rect 5582 9276 5890 9296
rect 5582 9274 5588 9276
rect 5644 9274 5668 9276
rect 5724 9274 5748 9276
rect 5804 9274 5828 9276
rect 5884 9274 5890 9276
rect 5644 9222 5646 9274
rect 5826 9222 5828 9274
rect 5582 9220 5588 9222
rect 5644 9220 5668 9222
rect 5724 9220 5748 9222
rect 5804 9220 5828 9222
rect 5884 9220 5890 9222
rect 5582 9200 5890 9220
rect 5582 8188 5890 8208
rect 5582 8186 5588 8188
rect 5644 8186 5668 8188
rect 5724 8186 5748 8188
rect 5804 8186 5828 8188
rect 5884 8186 5890 8188
rect 5644 8134 5646 8186
rect 5826 8134 5828 8186
rect 5582 8132 5588 8134
rect 5644 8132 5668 8134
rect 5724 8132 5748 8134
rect 5804 8132 5828 8134
rect 5884 8132 5890 8134
rect 5582 8112 5890 8132
rect 9220 7812 9272 7818
rect 9220 7754 9272 7760
rect 5582 7100 5890 7120
rect 5582 7098 5588 7100
rect 5644 7098 5668 7100
rect 5724 7098 5748 7100
rect 5804 7098 5828 7100
rect 5884 7098 5890 7100
rect 5644 7046 5646 7098
rect 5826 7046 5828 7098
rect 5582 7044 5588 7046
rect 5644 7044 5668 7046
rect 5724 7044 5748 7046
rect 5804 7044 5828 7046
rect 5884 7044 5890 7046
rect 5582 7024 5890 7044
rect 6184 6792 6236 6798
rect 6184 6734 6236 6740
rect 5582 6012 5890 6032
rect 5582 6010 5588 6012
rect 5644 6010 5668 6012
rect 5724 6010 5748 6012
rect 5804 6010 5828 6012
rect 5884 6010 5890 6012
rect 5644 5958 5646 6010
rect 5826 5958 5828 6010
rect 5582 5956 5588 5958
rect 5644 5956 5668 5958
rect 5724 5956 5748 5958
rect 5804 5956 5828 5958
rect 5884 5956 5890 5958
rect 5582 5936 5890 5956
rect 5582 4924 5890 4944
rect 5582 4922 5588 4924
rect 5644 4922 5668 4924
rect 5724 4922 5748 4924
rect 5804 4922 5828 4924
rect 5884 4922 5890 4924
rect 5644 4870 5646 4922
rect 5826 4870 5828 4922
rect 5582 4868 5588 4870
rect 5644 4868 5668 4870
rect 5724 4868 5748 4870
rect 5804 4868 5828 4870
rect 5884 4868 5890 4870
rect 5582 4848 5890 4868
rect 5582 3836 5890 3856
rect 5582 3834 5588 3836
rect 5644 3834 5668 3836
rect 5724 3834 5748 3836
rect 5804 3834 5828 3836
rect 5884 3834 5890 3836
rect 5644 3782 5646 3834
rect 5826 3782 5828 3834
rect 5582 3780 5588 3782
rect 5644 3780 5668 3782
rect 5724 3780 5748 3782
rect 5804 3780 5828 3782
rect 5884 3780 5890 3782
rect 5582 3760 5890 3780
rect 5448 3732 5500 3738
rect 5448 3674 5500 3680
rect 5356 3596 5408 3602
rect 5356 3538 5408 3544
rect 5908 3596 5960 3602
rect 5908 3538 5960 3544
rect 3698 3431 3754 3440
rect 3896 3454 4200 3482
rect 5172 3528 5224 3534
rect 5172 3470 5224 3476
rect 3424 2576 3476 2582
rect 3424 2518 3476 2524
rect 3436 2145 3464 2518
rect 3422 2136 3478 2145
rect 3422 2071 3478 2080
rect 3330 1456 3386 1465
rect 3330 1391 3386 1400
rect 3896 800 3924 3454
rect 4160 3392 4212 3398
rect 4160 3334 4212 3340
rect 4172 3126 4200 3334
rect 4160 3120 4212 3126
rect 4160 3062 4212 3068
rect 3976 2984 4028 2990
rect 3976 2926 4028 2932
rect 4528 2984 4580 2990
rect 4528 2926 4580 2932
rect 3988 2650 4016 2926
rect 3976 2644 4028 2650
rect 3976 2586 4028 2592
rect 4540 800 4568 2926
rect 5184 2650 5212 3470
rect 5582 2748 5890 2768
rect 5582 2746 5588 2748
rect 5644 2746 5668 2748
rect 5724 2746 5748 2748
rect 5804 2746 5828 2748
rect 5884 2746 5890 2748
rect 5644 2694 5646 2746
rect 5826 2694 5828 2746
rect 5582 2692 5588 2694
rect 5644 2692 5668 2694
rect 5724 2692 5748 2694
rect 5804 2692 5828 2694
rect 5884 2692 5890 2694
rect 5582 2672 5890 2692
rect 5172 2644 5224 2650
rect 5172 2586 5224 2592
rect 5920 1850 5948 3538
rect 6196 2446 6224 6734
rect 6276 5024 6328 5030
rect 6276 4966 6328 4972
rect 6288 4690 6316 4966
rect 6276 4684 6328 4690
rect 6276 4626 6328 4632
rect 9232 4146 9260 7754
rect 9220 4140 9272 4146
rect 9220 4082 9272 4088
rect 6368 3936 6420 3942
rect 6368 3878 6420 3884
rect 8668 3936 8720 3942
rect 8668 3878 8720 3884
rect 9312 3936 9364 3942
rect 9312 3878 9364 3884
rect 6380 3058 6408 3878
rect 8680 3058 8708 3878
rect 9324 3602 9352 3878
rect 9312 3596 9364 3602
rect 9312 3538 9364 3544
rect 8852 3392 8904 3398
rect 8852 3334 8904 3340
rect 8864 3126 8892 3334
rect 8852 3120 8904 3126
rect 8852 3062 8904 3068
rect 6368 3052 6420 3058
rect 6368 2994 6420 3000
rect 8668 3052 8720 3058
rect 8668 2994 8720 3000
rect 6552 2984 6604 2990
rect 6552 2926 6604 2932
rect 8392 2984 8444 2990
rect 8392 2926 8444 2932
rect 6460 2916 6512 2922
rect 6460 2858 6512 2864
rect 6184 2440 6236 2446
rect 6184 2382 6236 2388
rect 5828 1822 5948 1850
rect 5828 800 5856 1822
rect 6472 800 6500 2858
rect 6564 2650 6592 2926
rect 6552 2644 6604 2650
rect 6552 2586 6604 2592
rect 8404 800 8432 2926
rect 9508 2650 9536 23598
rect 12452 23118 12480 24006
rect 12532 23520 12584 23526
rect 12532 23462 12584 23468
rect 12164 23112 12216 23118
rect 12164 23054 12216 23060
rect 12440 23112 12492 23118
rect 12440 23054 12492 23060
rect 10214 22876 10522 22896
rect 10214 22874 10220 22876
rect 10276 22874 10300 22876
rect 10356 22874 10380 22876
rect 10436 22874 10460 22876
rect 10516 22874 10522 22876
rect 10276 22822 10278 22874
rect 10458 22822 10460 22874
rect 10214 22820 10220 22822
rect 10276 22820 10300 22822
rect 10356 22820 10380 22822
rect 10436 22820 10460 22822
rect 10516 22820 10522 22822
rect 10214 22800 10522 22820
rect 10214 21788 10522 21808
rect 10214 21786 10220 21788
rect 10276 21786 10300 21788
rect 10356 21786 10380 21788
rect 10436 21786 10460 21788
rect 10516 21786 10522 21788
rect 10276 21734 10278 21786
rect 10458 21734 10460 21786
rect 10214 21732 10220 21734
rect 10276 21732 10300 21734
rect 10356 21732 10380 21734
rect 10436 21732 10460 21734
rect 10516 21732 10522 21734
rect 10214 21712 10522 21732
rect 12072 20868 12124 20874
rect 12072 20810 12124 20816
rect 10214 20700 10522 20720
rect 10214 20698 10220 20700
rect 10276 20698 10300 20700
rect 10356 20698 10380 20700
rect 10436 20698 10460 20700
rect 10516 20698 10522 20700
rect 10276 20646 10278 20698
rect 10458 20646 10460 20698
rect 10214 20644 10220 20646
rect 10276 20644 10300 20646
rect 10356 20644 10380 20646
rect 10436 20644 10460 20646
rect 10516 20644 10522 20646
rect 10214 20624 10522 20644
rect 11888 20392 11940 20398
rect 11888 20334 11940 20340
rect 10214 19612 10522 19632
rect 10214 19610 10220 19612
rect 10276 19610 10300 19612
rect 10356 19610 10380 19612
rect 10436 19610 10460 19612
rect 10516 19610 10522 19612
rect 10276 19558 10278 19610
rect 10458 19558 10460 19610
rect 10214 19556 10220 19558
rect 10276 19556 10300 19558
rect 10356 19556 10380 19558
rect 10436 19556 10460 19558
rect 10516 19556 10522 19558
rect 10214 19536 10522 19556
rect 10214 18524 10522 18544
rect 10214 18522 10220 18524
rect 10276 18522 10300 18524
rect 10356 18522 10380 18524
rect 10436 18522 10460 18524
rect 10516 18522 10522 18524
rect 10276 18470 10278 18522
rect 10458 18470 10460 18522
rect 10214 18468 10220 18470
rect 10276 18468 10300 18470
rect 10356 18468 10380 18470
rect 10436 18468 10460 18470
rect 10516 18468 10522 18470
rect 10214 18448 10522 18468
rect 11244 18080 11296 18086
rect 11244 18022 11296 18028
rect 11256 17678 11284 18022
rect 11900 17678 11928 20334
rect 12084 20058 12112 20810
rect 12176 20534 12204 23054
rect 12544 22710 12572 23462
rect 12624 22976 12676 22982
rect 12624 22918 12676 22924
rect 12636 22778 12664 22918
rect 12624 22772 12676 22778
rect 12624 22714 12676 22720
rect 12728 22710 12756 25842
rect 13268 25696 13320 25702
rect 13268 25638 13320 25644
rect 13280 25294 13308 25638
rect 13268 25288 13320 25294
rect 13268 25230 13320 25236
rect 13372 24750 13400 28970
rect 13820 28416 13872 28422
rect 13820 28358 13872 28364
rect 13636 28076 13688 28082
rect 13636 28018 13688 28024
rect 13648 27674 13676 28018
rect 13636 27668 13688 27674
rect 13636 27610 13688 27616
rect 13832 27470 13860 28358
rect 14016 27878 14044 29514
rect 14384 28490 14412 30670
rect 14648 30660 14700 30666
rect 14648 30602 14700 30608
rect 14556 30048 14608 30054
rect 14556 29990 14608 29996
rect 14464 29776 14516 29782
rect 14464 29718 14516 29724
rect 14188 28484 14240 28490
rect 14188 28426 14240 28432
rect 14372 28484 14424 28490
rect 14372 28426 14424 28432
rect 14004 27872 14056 27878
rect 14004 27814 14056 27820
rect 13912 27600 13964 27606
rect 13912 27542 13964 27548
rect 13820 27464 13872 27470
rect 13820 27406 13872 27412
rect 13176 24744 13228 24750
rect 13176 24686 13228 24692
rect 13360 24744 13412 24750
rect 13360 24686 13412 24692
rect 12900 24200 12952 24206
rect 12900 24142 12952 24148
rect 12808 23656 12860 23662
rect 12808 23598 12860 23604
rect 12532 22704 12584 22710
rect 12532 22646 12584 22652
rect 12716 22704 12768 22710
rect 12716 22646 12768 22652
rect 12728 22098 12756 22646
rect 12716 22092 12768 22098
rect 12716 22034 12768 22040
rect 12728 20874 12756 22034
rect 12716 20868 12768 20874
rect 12716 20810 12768 20816
rect 12624 20800 12676 20806
rect 12624 20742 12676 20748
rect 12164 20528 12216 20534
rect 12164 20470 12216 20476
rect 12636 20466 12664 20742
rect 12624 20460 12676 20466
rect 12624 20402 12676 20408
rect 12072 20052 12124 20058
rect 12072 19994 12124 20000
rect 12820 19922 12848 23598
rect 12912 22778 12940 24142
rect 13188 23866 13216 24686
rect 13176 23860 13228 23866
rect 13176 23802 13228 23808
rect 13372 23662 13400 24686
rect 13544 23724 13596 23730
rect 13544 23666 13596 23672
rect 13360 23656 13412 23662
rect 13360 23598 13412 23604
rect 13556 23322 13584 23666
rect 13544 23316 13596 23322
rect 13544 23258 13596 23264
rect 12900 22772 12952 22778
rect 12900 22714 12952 22720
rect 13360 22432 13412 22438
rect 13360 22374 13412 22380
rect 13372 21554 13400 22374
rect 13924 22094 13952 27542
rect 14016 27470 14044 27814
rect 14200 27674 14228 28426
rect 14188 27668 14240 27674
rect 14188 27610 14240 27616
rect 14004 27464 14056 27470
rect 14004 27406 14056 27412
rect 14016 25838 14044 27406
rect 14384 27402 14412 28426
rect 14476 27606 14504 29718
rect 14568 29714 14596 29990
rect 14660 29850 14688 30602
rect 15476 30592 15528 30598
rect 15476 30534 15528 30540
rect 16672 30592 16724 30598
rect 16672 30534 16724 30540
rect 15488 30326 15516 30534
rect 15476 30320 15528 30326
rect 15476 30262 15528 30268
rect 16684 30258 16712 30534
rect 16672 30252 16724 30258
rect 16672 30194 16724 30200
rect 16120 30048 16172 30054
rect 16120 29990 16172 29996
rect 16948 30048 17000 30054
rect 16948 29990 17000 29996
rect 14846 29948 15154 29968
rect 14846 29946 14852 29948
rect 14908 29946 14932 29948
rect 14988 29946 15012 29948
rect 15068 29946 15092 29948
rect 15148 29946 15154 29948
rect 14908 29894 14910 29946
rect 15090 29894 15092 29946
rect 14846 29892 14852 29894
rect 14908 29892 14932 29894
rect 14988 29892 15012 29894
rect 15068 29892 15092 29894
rect 15148 29892 15154 29894
rect 14846 29872 15154 29892
rect 14648 29844 14700 29850
rect 14648 29786 14700 29792
rect 14556 29708 14608 29714
rect 14556 29650 14608 29656
rect 16132 29510 16160 29990
rect 16580 29844 16632 29850
rect 16580 29786 16632 29792
rect 16120 29504 16172 29510
rect 16120 29446 16172 29452
rect 14846 28860 15154 28880
rect 14846 28858 14852 28860
rect 14908 28858 14932 28860
rect 14988 28858 15012 28860
rect 15068 28858 15092 28860
rect 15148 28858 15154 28860
rect 14908 28806 14910 28858
rect 15090 28806 15092 28858
rect 14846 28804 14852 28806
rect 14908 28804 14932 28806
rect 14988 28804 15012 28806
rect 15068 28804 15092 28806
rect 15148 28804 15154 28806
rect 14846 28784 15154 28804
rect 14648 28144 14700 28150
rect 14648 28086 14700 28092
rect 15752 28144 15804 28150
rect 15752 28086 15804 28092
rect 14464 27600 14516 27606
rect 14464 27542 14516 27548
rect 14660 27538 14688 28086
rect 14740 27872 14792 27878
rect 14740 27814 14792 27820
rect 14648 27532 14700 27538
rect 14648 27474 14700 27480
rect 14372 27396 14424 27402
rect 14372 27338 14424 27344
rect 14752 27334 14780 27814
rect 14846 27772 15154 27792
rect 14846 27770 14852 27772
rect 14908 27770 14932 27772
rect 14988 27770 15012 27772
rect 15068 27770 15092 27772
rect 15148 27770 15154 27772
rect 14908 27718 14910 27770
rect 15090 27718 15092 27770
rect 14846 27716 14852 27718
rect 14908 27716 14932 27718
rect 14988 27716 15012 27718
rect 15068 27716 15092 27718
rect 15148 27716 15154 27718
rect 14846 27696 15154 27716
rect 15108 27464 15160 27470
rect 15108 27406 15160 27412
rect 14096 27328 14148 27334
rect 14096 27270 14148 27276
rect 14740 27328 14792 27334
rect 14740 27270 14792 27276
rect 14004 25832 14056 25838
rect 14004 25774 14056 25780
rect 14016 25362 14044 25774
rect 14004 25356 14056 25362
rect 14004 25298 14056 25304
rect 14108 22094 14136 27270
rect 15120 27062 15148 27406
rect 15108 27056 15160 27062
rect 15108 26998 15160 27004
rect 15660 26920 15712 26926
rect 15660 26862 15712 26868
rect 14846 26684 15154 26704
rect 14846 26682 14852 26684
rect 14908 26682 14932 26684
rect 14988 26682 15012 26684
rect 15068 26682 15092 26684
rect 15148 26682 15154 26684
rect 14908 26630 14910 26682
rect 15090 26630 15092 26682
rect 14846 26628 14852 26630
rect 14908 26628 14932 26630
rect 14988 26628 15012 26630
rect 15068 26628 15092 26630
rect 15148 26628 15154 26630
rect 14846 26608 15154 26628
rect 15672 26382 15700 26862
rect 14740 26376 14792 26382
rect 14740 26318 14792 26324
rect 15568 26376 15620 26382
rect 15568 26318 15620 26324
rect 15660 26376 15712 26382
rect 15660 26318 15712 26324
rect 14556 26240 14608 26246
rect 14556 26182 14608 26188
rect 14568 25974 14596 26182
rect 14556 25968 14608 25974
rect 14556 25910 14608 25916
rect 14752 25498 14780 26318
rect 15384 26240 15436 26246
rect 15384 26182 15436 26188
rect 14846 25596 15154 25616
rect 14846 25594 14852 25596
rect 14908 25594 14932 25596
rect 14988 25594 15012 25596
rect 15068 25594 15092 25596
rect 15148 25594 15154 25596
rect 14908 25542 14910 25594
rect 15090 25542 15092 25594
rect 14846 25540 14852 25542
rect 14908 25540 14932 25542
rect 14988 25540 15012 25542
rect 15068 25540 15092 25542
rect 15148 25540 15154 25542
rect 14846 25520 15154 25540
rect 15396 25498 15424 26182
rect 15580 26042 15608 26318
rect 15568 26036 15620 26042
rect 15568 25978 15620 25984
rect 14740 25492 14792 25498
rect 14740 25434 14792 25440
rect 15384 25492 15436 25498
rect 15384 25434 15436 25440
rect 15200 25152 15252 25158
rect 15200 25094 15252 25100
rect 15476 25152 15528 25158
rect 15476 25094 15528 25100
rect 15212 24954 15240 25094
rect 15200 24948 15252 24954
rect 15200 24890 15252 24896
rect 15488 24818 15516 25094
rect 15476 24812 15528 24818
rect 15528 24772 15608 24800
rect 15476 24754 15528 24760
rect 14846 24508 15154 24528
rect 14846 24506 14852 24508
rect 14908 24506 14932 24508
rect 14988 24506 15012 24508
rect 15068 24506 15092 24508
rect 15148 24506 15154 24508
rect 14908 24454 14910 24506
rect 15090 24454 15092 24506
rect 14846 24452 14852 24454
rect 14908 24452 14932 24454
rect 14988 24452 15012 24454
rect 15068 24452 15092 24454
rect 15148 24452 15154 24454
rect 14846 24432 15154 24452
rect 15292 24200 15344 24206
rect 15292 24142 15344 24148
rect 15108 24064 15160 24070
rect 15108 24006 15160 24012
rect 15120 23798 15148 24006
rect 15108 23792 15160 23798
rect 15108 23734 15160 23740
rect 14740 23656 14792 23662
rect 14740 23598 14792 23604
rect 14752 23050 14780 23598
rect 14846 23420 15154 23440
rect 14846 23418 14852 23420
rect 14908 23418 14932 23420
rect 14988 23418 15012 23420
rect 15068 23418 15092 23420
rect 15148 23418 15154 23420
rect 14908 23366 14910 23418
rect 15090 23366 15092 23418
rect 14846 23364 14852 23366
rect 14908 23364 14932 23366
rect 14988 23364 15012 23366
rect 15068 23364 15092 23366
rect 15148 23364 15154 23366
rect 14846 23344 15154 23364
rect 15304 23322 15332 24142
rect 15292 23316 15344 23322
rect 15292 23258 15344 23264
rect 14740 23044 14792 23050
rect 14740 22986 14792 22992
rect 14752 22642 14780 22986
rect 14464 22636 14516 22642
rect 14464 22578 14516 22584
rect 14740 22636 14792 22642
rect 14740 22578 14792 22584
rect 14476 22234 14504 22578
rect 14846 22332 15154 22352
rect 14846 22330 14852 22332
rect 14908 22330 14932 22332
rect 14988 22330 15012 22332
rect 15068 22330 15092 22332
rect 15148 22330 15154 22332
rect 14908 22278 14910 22330
rect 15090 22278 15092 22330
rect 14846 22276 14852 22278
rect 14908 22276 14932 22278
rect 14988 22276 15012 22278
rect 15068 22276 15092 22278
rect 15148 22276 15154 22278
rect 14846 22256 15154 22276
rect 14464 22228 14516 22234
rect 14464 22170 14516 22176
rect 13832 22066 13952 22094
rect 14016 22066 14136 22094
rect 13360 21548 13412 21554
rect 13360 21490 13412 21496
rect 12808 19916 12860 19922
rect 12808 19858 12860 19864
rect 12716 19712 12768 19718
rect 12716 19654 12768 19660
rect 12728 18630 12756 19654
rect 12716 18624 12768 18630
rect 12716 18566 12768 18572
rect 13372 18290 13400 21490
rect 12348 18284 12400 18290
rect 12348 18226 12400 18232
rect 12440 18284 12492 18290
rect 12440 18226 12492 18232
rect 13360 18284 13412 18290
rect 13360 18226 13412 18232
rect 11244 17672 11296 17678
rect 11244 17614 11296 17620
rect 11888 17672 11940 17678
rect 11888 17614 11940 17620
rect 10214 17436 10522 17456
rect 10214 17434 10220 17436
rect 10276 17434 10300 17436
rect 10356 17434 10380 17436
rect 10436 17434 10460 17436
rect 10516 17434 10522 17436
rect 10276 17382 10278 17434
rect 10458 17382 10460 17434
rect 10214 17380 10220 17382
rect 10276 17380 10300 17382
rect 10356 17380 10380 17382
rect 10436 17380 10460 17382
rect 10516 17380 10522 17382
rect 10214 17360 10522 17380
rect 10214 16348 10522 16368
rect 10214 16346 10220 16348
rect 10276 16346 10300 16348
rect 10356 16346 10380 16348
rect 10436 16346 10460 16348
rect 10516 16346 10522 16348
rect 10276 16294 10278 16346
rect 10458 16294 10460 16346
rect 10214 16292 10220 16294
rect 10276 16292 10300 16294
rect 10356 16292 10380 16294
rect 10436 16292 10460 16294
rect 10516 16292 10522 16294
rect 10214 16272 10522 16292
rect 10214 15260 10522 15280
rect 10214 15258 10220 15260
rect 10276 15258 10300 15260
rect 10356 15258 10380 15260
rect 10436 15258 10460 15260
rect 10516 15258 10522 15260
rect 10276 15206 10278 15258
rect 10458 15206 10460 15258
rect 10214 15204 10220 15206
rect 10276 15204 10300 15206
rect 10356 15204 10380 15206
rect 10436 15204 10460 15206
rect 10516 15204 10522 15206
rect 10214 15184 10522 15204
rect 11900 15026 11928 17614
rect 12360 17338 12388 18226
rect 12348 17332 12400 17338
rect 12348 17274 12400 17280
rect 12164 15904 12216 15910
rect 12164 15846 12216 15852
rect 12176 15502 12204 15846
rect 12452 15570 12480 18226
rect 13268 18080 13320 18086
rect 13268 18022 13320 18028
rect 13280 17542 13308 18022
rect 13268 17536 13320 17542
rect 13268 17478 13320 17484
rect 13280 17338 13308 17478
rect 13268 17332 13320 17338
rect 13268 17274 13320 17280
rect 12900 17128 12952 17134
rect 12900 17070 12952 17076
rect 12912 16046 12940 17070
rect 13280 17066 13308 17274
rect 13372 17270 13400 18226
rect 13360 17264 13412 17270
rect 13360 17206 13412 17212
rect 13268 17060 13320 17066
rect 13268 17002 13320 17008
rect 13360 16108 13412 16114
rect 13360 16050 13412 16056
rect 12900 16040 12952 16046
rect 12900 15982 12952 15988
rect 13372 15638 13400 16050
rect 13360 15632 13412 15638
rect 13360 15574 13412 15580
rect 12440 15564 12492 15570
rect 12440 15506 12492 15512
rect 12164 15496 12216 15502
rect 12164 15438 12216 15444
rect 12808 15360 12860 15366
rect 12808 15302 12860 15308
rect 12820 15094 12848 15302
rect 13372 15162 13400 15574
rect 13360 15156 13412 15162
rect 13360 15098 13412 15104
rect 12808 15088 12860 15094
rect 12808 15030 12860 15036
rect 11888 15020 11940 15026
rect 11888 14962 11940 14968
rect 10214 14172 10522 14192
rect 10214 14170 10220 14172
rect 10276 14170 10300 14172
rect 10356 14170 10380 14172
rect 10436 14170 10460 14172
rect 10516 14170 10522 14172
rect 10276 14118 10278 14170
rect 10458 14118 10460 14170
rect 10214 14116 10220 14118
rect 10276 14116 10300 14118
rect 10356 14116 10380 14118
rect 10436 14116 10460 14118
rect 10516 14116 10522 14118
rect 10214 14096 10522 14116
rect 11900 13938 11928 14962
rect 11888 13932 11940 13938
rect 11888 13874 11940 13880
rect 10214 13084 10522 13104
rect 10214 13082 10220 13084
rect 10276 13082 10300 13084
rect 10356 13082 10380 13084
rect 10436 13082 10460 13084
rect 10516 13082 10522 13084
rect 10276 13030 10278 13082
rect 10458 13030 10460 13082
rect 10214 13028 10220 13030
rect 10276 13028 10300 13030
rect 10356 13028 10380 13030
rect 10436 13028 10460 13030
rect 10516 13028 10522 13030
rect 10214 13008 10522 13028
rect 10214 11996 10522 12016
rect 10214 11994 10220 11996
rect 10276 11994 10300 11996
rect 10356 11994 10380 11996
rect 10436 11994 10460 11996
rect 10516 11994 10522 11996
rect 10276 11942 10278 11994
rect 10458 11942 10460 11994
rect 10214 11940 10220 11942
rect 10276 11940 10300 11942
rect 10356 11940 10380 11942
rect 10436 11940 10460 11942
rect 10516 11940 10522 11942
rect 10214 11920 10522 11940
rect 13832 11218 13860 22066
rect 13912 17604 13964 17610
rect 13912 17546 13964 17552
rect 13924 17338 13952 17546
rect 13912 17332 13964 17338
rect 13912 17274 13964 17280
rect 14016 17066 14044 22066
rect 14096 22024 14148 22030
rect 14096 21966 14148 21972
rect 14108 21078 14136 21966
rect 15580 21554 15608 24772
rect 15672 24070 15700 26318
rect 15764 25226 15792 28086
rect 15936 27872 15988 27878
rect 15936 27814 15988 27820
rect 15948 27130 15976 27814
rect 15936 27124 15988 27130
rect 15936 27066 15988 27072
rect 15936 26988 15988 26994
rect 15936 26930 15988 26936
rect 15948 26858 15976 26930
rect 15936 26852 15988 26858
rect 15936 26794 15988 26800
rect 15948 26314 15976 26794
rect 15936 26308 15988 26314
rect 15936 26250 15988 26256
rect 15948 25294 15976 26250
rect 15936 25288 15988 25294
rect 15936 25230 15988 25236
rect 15752 25220 15804 25226
rect 15752 25162 15804 25168
rect 16028 25220 16080 25226
rect 16028 25162 16080 25168
rect 15660 24064 15712 24070
rect 15660 24006 15712 24012
rect 15672 23254 15700 24006
rect 15660 23248 15712 23254
rect 15660 23190 15712 23196
rect 15384 21548 15436 21554
rect 15384 21490 15436 21496
rect 15568 21548 15620 21554
rect 15568 21490 15620 21496
rect 14740 21344 14792 21350
rect 14740 21286 14792 21292
rect 14752 21146 14780 21286
rect 14846 21244 15154 21264
rect 14846 21242 14852 21244
rect 14908 21242 14932 21244
rect 14988 21242 15012 21244
rect 15068 21242 15092 21244
rect 15148 21242 15154 21244
rect 14908 21190 14910 21242
rect 15090 21190 15092 21242
rect 14846 21188 14852 21190
rect 14908 21188 14932 21190
rect 14988 21188 15012 21190
rect 15068 21188 15092 21190
rect 15148 21188 15154 21190
rect 14846 21168 15154 21188
rect 14740 21140 14792 21146
rect 14740 21082 14792 21088
rect 14096 21072 14148 21078
rect 14096 21014 14148 21020
rect 14280 20936 14332 20942
rect 14280 20878 14332 20884
rect 14096 20800 14148 20806
rect 14096 20742 14148 20748
rect 14108 20534 14136 20742
rect 14096 20528 14148 20534
rect 14096 20470 14148 20476
rect 14096 20256 14148 20262
rect 14096 20198 14148 20204
rect 14108 19786 14136 20198
rect 14292 20058 14320 20878
rect 14740 20800 14792 20806
rect 14740 20742 14792 20748
rect 15292 20800 15344 20806
rect 15292 20742 15344 20748
rect 14280 20052 14332 20058
rect 14280 19994 14332 20000
rect 14752 19854 14780 20742
rect 15200 20256 15252 20262
rect 15200 20198 15252 20204
rect 14846 20156 15154 20176
rect 14846 20154 14852 20156
rect 14908 20154 14932 20156
rect 14988 20154 15012 20156
rect 15068 20154 15092 20156
rect 15148 20154 15154 20156
rect 14908 20102 14910 20154
rect 15090 20102 15092 20154
rect 14846 20100 14852 20102
rect 14908 20100 14932 20102
rect 14988 20100 15012 20102
rect 15068 20100 15092 20102
rect 15148 20100 15154 20102
rect 14846 20080 15154 20100
rect 14188 19848 14240 19854
rect 14188 19790 14240 19796
rect 14740 19848 14792 19854
rect 14740 19790 14792 19796
rect 14096 19780 14148 19786
rect 14096 19722 14148 19728
rect 14108 19258 14136 19722
rect 14200 19360 14228 19790
rect 15212 19378 15240 20198
rect 15304 20058 15332 20742
rect 15396 20262 15424 21490
rect 15476 20868 15528 20874
rect 15476 20810 15528 20816
rect 15384 20256 15436 20262
rect 15384 20198 15436 20204
rect 15292 20052 15344 20058
rect 15292 19994 15344 20000
rect 14280 19372 14332 19378
rect 14200 19332 14280 19360
rect 14280 19314 14332 19320
rect 15200 19372 15252 19378
rect 15200 19314 15252 19320
rect 14108 19230 14228 19258
rect 14096 18080 14148 18086
rect 14096 18022 14148 18028
rect 14108 17270 14136 18022
rect 14200 17678 14228 19230
rect 14188 17672 14240 17678
rect 14188 17614 14240 17620
rect 14096 17264 14148 17270
rect 14096 17206 14148 17212
rect 14004 17060 14056 17066
rect 14004 17002 14056 17008
rect 14200 16794 14228 17614
rect 14292 17542 14320 19314
rect 14846 19068 15154 19088
rect 14846 19066 14852 19068
rect 14908 19066 14932 19068
rect 14988 19066 15012 19068
rect 15068 19066 15092 19068
rect 15148 19066 15154 19068
rect 14908 19014 14910 19066
rect 15090 19014 15092 19066
rect 14846 19012 14852 19014
rect 14908 19012 14932 19014
rect 14988 19012 15012 19014
rect 15068 19012 15092 19014
rect 15148 19012 15154 19014
rect 14846 18992 15154 19012
rect 14660 18290 14872 18306
rect 14372 18284 14424 18290
rect 14556 18284 14608 18290
rect 14372 18226 14424 18232
rect 14476 18244 14556 18272
rect 14384 17678 14412 18226
rect 14372 17672 14424 17678
rect 14372 17614 14424 17620
rect 14280 17536 14332 17542
rect 14280 17478 14332 17484
rect 14188 16788 14240 16794
rect 14188 16730 14240 16736
rect 14292 16658 14320 17478
rect 14188 16652 14240 16658
rect 14188 16594 14240 16600
rect 14280 16652 14332 16658
rect 14280 16594 14332 16600
rect 14096 16584 14148 16590
rect 14096 16526 14148 16532
rect 14108 15706 14136 16526
rect 14096 15700 14148 15706
rect 14096 15642 14148 15648
rect 14200 15638 14228 16594
rect 14188 15632 14240 15638
rect 14188 15574 14240 15580
rect 14384 15570 14412 17614
rect 14476 17134 14504 18244
rect 14556 18226 14608 18232
rect 14660 18284 14884 18290
rect 14660 18278 14832 18284
rect 14556 18148 14608 18154
rect 14556 18090 14608 18096
rect 14568 17338 14596 18090
rect 14660 17542 14688 18278
rect 14832 18226 14884 18232
rect 14740 18216 14792 18222
rect 14740 18158 14792 18164
rect 14752 17746 14780 18158
rect 14846 17980 15154 18000
rect 14846 17978 14852 17980
rect 14908 17978 14932 17980
rect 14988 17978 15012 17980
rect 15068 17978 15092 17980
rect 15148 17978 15154 17980
rect 14908 17926 14910 17978
rect 15090 17926 15092 17978
rect 14846 17924 14852 17926
rect 14908 17924 14932 17926
rect 14988 17924 15012 17926
rect 15068 17924 15092 17926
rect 15148 17924 15154 17926
rect 14846 17904 15154 17924
rect 14740 17740 14792 17746
rect 14740 17682 14792 17688
rect 14648 17536 14700 17542
rect 14648 17478 14700 17484
rect 14556 17332 14608 17338
rect 14556 17274 14608 17280
rect 14464 17128 14516 17134
rect 14464 17070 14516 17076
rect 14568 16794 14596 17274
rect 14660 17202 14688 17478
rect 14752 17338 14780 17682
rect 14740 17332 14792 17338
rect 14740 17274 14792 17280
rect 14648 17196 14700 17202
rect 14648 17138 14700 17144
rect 14846 16892 15154 16912
rect 14846 16890 14852 16892
rect 14908 16890 14932 16892
rect 14988 16890 15012 16892
rect 15068 16890 15092 16892
rect 15148 16890 15154 16892
rect 14908 16838 14910 16890
rect 15090 16838 15092 16890
rect 14846 16836 14852 16838
rect 14908 16836 14932 16838
rect 14988 16836 15012 16838
rect 15068 16836 15092 16838
rect 15148 16836 15154 16838
rect 14846 16816 15154 16836
rect 14556 16788 14608 16794
rect 14556 16730 14608 16736
rect 14556 16040 14608 16046
rect 14556 15982 14608 15988
rect 14372 15564 14424 15570
rect 14372 15506 14424 15512
rect 14568 15434 14596 15982
rect 14846 15804 15154 15824
rect 14846 15802 14852 15804
rect 14908 15802 14932 15804
rect 14988 15802 15012 15804
rect 15068 15802 15092 15804
rect 15148 15802 15154 15804
rect 14908 15750 14910 15802
rect 15090 15750 15092 15802
rect 14846 15748 14852 15750
rect 14908 15748 14932 15750
rect 14988 15748 15012 15750
rect 15068 15748 15092 15750
rect 15148 15748 15154 15750
rect 14846 15728 15154 15748
rect 15016 15632 15068 15638
rect 15016 15574 15068 15580
rect 14556 15428 14608 15434
rect 14556 15370 14608 15376
rect 14280 14272 14332 14278
rect 14280 14214 14332 14220
rect 14096 13932 14148 13938
rect 14096 13874 14148 13880
rect 14108 13530 14136 13874
rect 14096 13524 14148 13530
rect 14096 13466 14148 13472
rect 14292 13326 14320 14214
rect 14568 13870 14596 15370
rect 15028 15026 15056 15574
rect 15304 15026 15332 19994
rect 15488 19922 15516 20810
rect 15580 20466 15608 21490
rect 15764 20874 15792 25162
rect 16040 24070 16068 25162
rect 16028 24064 16080 24070
rect 16028 24006 16080 24012
rect 16132 22094 16160 29446
rect 16592 29034 16620 29786
rect 16960 29646 16988 29990
rect 16948 29640 17000 29646
rect 16948 29582 17000 29588
rect 16580 29028 16632 29034
rect 16580 28970 16632 28976
rect 16764 28008 16816 28014
rect 16764 27950 16816 27956
rect 16672 27872 16724 27878
rect 16672 27814 16724 27820
rect 16684 27470 16712 27814
rect 16672 27464 16724 27470
rect 16672 27406 16724 27412
rect 16776 27130 16804 27950
rect 16764 27124 16816 27130
rect 16764 27066 16816 27072
rect 16488 26444 16540 26450
rect 16488 26386 16540 26392
rect 16500 25430 16528 26386
rect 16580 26376 16632 26382
rect 16580 26318 16632 26324
rect 16488 25424 16540 25430
rect 16488 25366 16540 25372
rect 16212 25152 16264 25158
rect 16212 25094 16264 25100
rect 16224 24342 16252 25094
rect 16592 24750 16620 26318
rect 16672 24812 16724 24818
rect 16672 24754 16724 24760
rect 16580 24744 16632 24750
rect 16580 24686 16632 24692
rect 16580 24608 16632 24614
rect 16580 24550 16632 24556
rect 16212 24336 16264 24342
rect 16212 24278 16264 24284
rect 16592 24206 16620 24550
rect 16684 24410 16712 24754
rect 16948 24744 17000 24750
rect 16948 24686 17000 24692
rect 16672 24404 16724 24410
rect 16672 24346 16724 24352
rect 16580 24200 16632 24206
rect 16580 24142 16632 24148
rect 16592 23526 16620 24142
rect 16856 24132 16908 24138
rect 16856 24074 16908 24080
rect 16764 24064 16816 24070
rect 16764 24006 16816 24012
rect 16776 23730 16804 24006
rect 16764 23724 16816 23730
rect 16764 23666 16816 23672
rect 16580 23520 16632 23526
rect 16580 23462 16632 23468
rect 16592 23118 16620 23462
rect 16672 23316 16724 23322
rect 16672 23258 16724 23264
rect 16580 23112 16632 23118
rect 16580 23054 16632 23060
rect 16132 22066 16252 22094
rect 16028 20936 16080 20942
rect 16028 20878 16080 20884
rect 15752 20868 15804 20874
rect 15752 20810 15804 20816
rect 15568 20460 15620 20466
rect 15568 20402 15620 20408
rect 15936 20460 15988 20466
rect 15936 20402 15988 20408
rect 15752 20256 15804 20262
rect 15752 20198 15804 20204
rect 15476 19916 15528 19922
rect 15476 19858 15528 19864
rect 15764 19854 15792 20198
rect 15844 19916 15896 19922
rect 15844 19858 15896 19864
rect 15752 19848 15804 19854
rect 15752 19790 15804 19796
rect 15384 19780 15436 19786
rect 15384 19722 15436 19728
rect 15396 16590 15424 19722
rect 15568 17196 15620 17202
rect 15568 17138 15620 17144
rect 15476 17128 15528 17134
rect 15476 17070 15528 17076
rect 15488 16658 15516 17070
rect 15580 17066 15608 17138
rect 15568 17060 15620 17066
rect 15568 17002 15620 17008
rect 15476 16652 15528 16658
rect 15476 16594 15528 16600
rect 15384 16584 15436 16590
rect 15384 16526 15436 16532
rect 15396 15502 15424 16526
rect 15384 15496 15436 15502
rect 15384 15438 15436 15444
rect 15488 15450 15516 16594
rect 15660 16516 15712 16522
rect 15660 16458 15712 16464
rect 15672 16250 15700 16458
rect 15660 16244 15712 16250
rect 15660 16186 15712 16192
rect 15672 15484 15700 16186
rect 15752 15496 15804 15502
rect 15672 15456 15752 15484
rect 15488 15422 15608 15450
rect 15752 15438 15804 15444
rect 15476 15360 15528 15366
rect 15476 15302 15528 15308
rect 15016 15020 15068 15026
rect 15016 14962 15068 14968
rect 15292 15020 15344 15026
rect 15292 14962 15344 14968
rect 15200 14816 15252 14822
rect 15200 14758 15252 14764
rect 14846 14716 15154 14736
rect 14846 14714 14852 14716
rect 14908 14714 14932 14716
rect 14988 14714 15012 14716
rect 15068 14714 15092 14716
rect 15148 14714 15154 14716
rect 14908 14662 14910 14714
rect 15090 14662 15092 14714
rect 14846 14660 14852 14662
rect 14908 14660 14932 14662
rect 14988 14660 15012 14662
rect 15068 14660 15092 14662
rect 15148 14660 15154 14662
rect 14846 14640 15154 14660
rect 15212 14346 15240 14758
rect 15488 14618 15516 15302
rect 15476 14612 15528 14618
rect 15476 14554 15528 14560
rect 15200 14340 15252 14346
rect 15200 14282 15252 14288
rect 15384 14340 15436 14346
rect 15384 14282 15436 14288
rect 14740 14000 14792 14006
rect 14740 13942 14792 13948
rect 14556 13864 14608 13870
rect 14556 13806 14608 13812
rect 14280 13320 14332 13326
rect 14280 13262 14332 13268
rect 14752 12850 14780 13942
rect 14846 13628 15154 13648
rect 14846 13626 14852 13628
rect 14908 13626 14932 13628
rect 14988 13626 15012 13628
rect 15068 13626 15092 13628
rect 15148 13626 15154 13628
rect 14908 13574 14910 13626
rect 15090 13574 15092 13626
rect 14846 13572 14852 13574
rect 14908 13572 14932 13574
rect 14988 13572 15012 13574
rect 15068 13572 15092 13574
rect 15148 13572 15154 13574
rect 14846 13552 15154 13572
rect 15396 13258 15424 14282
rect 15488 13938 15516 14554
rect 15580 14414 15608 15422
rect 15856 15314 15884 19858
rect 15948 19854 15976 20402
rect 16040 20262 16068 20878
rect 16028 20256 16080 20262
rect 16028 20198 16080 20204
rect 15936 19848 15988 19854
rect 15936 19790 15988 19796
rect 16040 16114 16068 20198
rect 16120 17536 16172 17542
rect 16120 17478 16172 17484
rect 16132 16794 16160 17478
rect 16224 16810 16252 22066
rect 16684 19990 16712 23258
rect 16764 23044 16816 23050
rect 16764 22986 16816 22992
rect 16776 21622 16804 22986
rect 16764 21616 16816 21622
rect 16764 21558 16816 21564
rect 16776 21146 16804 21558
rect 16764 21140 16816 21146
rect 16764 21082 16816 21088
rect 16868 20942 16896 24074
rect 16960 23050 16988 24686
rect 17132 23724 17184 23730
rect 17132 23666 17184 23672
rect 17144 23118 17172 23666
rect 17132 23112 17184 23118
rect 17132 23054 17184 23060
rect 16948 23044 17000 23050
rect 16948 22986 17000 22992
rect 17236 22098 17264 30670
rect 17316 30660 17368 30666
rect 17316 30602 17368 30608
rect 17328 30394 17356 30602
rect 17316 30388 17368 30394
rect 17316 30330 17368 30336
rect 17604 28490 17632 31622
rect 17776 30320 17828 30326
rect 17776 30262 17828 30268
rect 17788 29510 17816 30262
rect 17880 30190 17908 31826
rect 17868 30184 17920 30190
rect 17868 30126 17920 30132
rect 17880 29850 17908 30126
rect 17868 29844 17920 29850
rect 17868 29786 17920 29792
rect 17776 29504 17828 29510
rect 17776 29446 17828 29452
rect 17592 28484 17644 28490
rect 17592 28426 17644 28432
rect 17316 27600 17368 27606
rect 17316 27542 17368 27548
rect 17328 26994 17356 27542
rect 17316 26988 17368 26994
rect 17316 26930 17368 26936
rect 17604 26858 17632 28426
rect 17788 28014 17816 29446
rect 17868 28688 17920 28694
rect 17868 28630 17920 28636
rect 17776 28008 17828 28014
rect 17776 27950 17828 27956
rect 17684 27940 17736 27946
rect 17684 27882 17736 27888
rect 17592 26852 17644 26858
rect 17592 26794 17644 26800
rect 17696 26450 17724 27882
rect 17788 26518 17816 27950
rect 17880 27538 17908 28630
rect 18052 28076 18104 28082
rect 18052 28018 18104 28024
rect 18064 27878 18092 28018
rect 18052 27872 18104 27878
rect 18052 27814 18104 27820
rect 17868 27532 17920 27538
rect 17868 27474 17920 27480
rect 17880 26994 17908 27474
rect 17868 26988 17920 26994
rect 17868 26930 17920 26936
rect 17776 26512 17828 26518
rect 17776 26454 17828 26460
rect 17684 26444 17736 26450
rect 17684 26386 17736 26392
rect 17868 25900 17920 25906
rect 17868 25842 17920 25848
rect 17776 25696 17828 25702
rect 17776 25638 17828 25644
rect 17408 24812 17460 24818
rect 17408 24754 17460 24760
rect 17684 24812 17736 24818
rect 17684 24754 17736 24760
rect 17316 24744 17368 24750
rect 17316 24686 17368 24692
rect 17328 24614 17356 24686
rect 17316 24608 17368 24614
rect 17316 24550 17368 24556
rect 17328 23050 17356 24550
rect 17420 24070 17448 24754
rect 17408 24064 17460 24070
rect 17408 24006 17460 24012
rect 17420 23050 17448 24006
rect 17696 23866 17724 24754
rect 17684 23860 17736 23866
rect 17684 23802 17736 23808
rect 17696 23322 17724 23802
rect 17684 23316 17736 23322
rect 17684 23258 17736 23264
rect 17316 23044 17368 23050
rect 17316 22986 17368 22992
rect 17408 23044 17460 23050
rect 17408 22986 17460 22992
rect 17684 22976 17736 22982
rect 17684 22918 17736 22924
rect 17224 22092 17276 22098
rect 17224 22034 17276 22040
rect 17236 21690 17264 22034
rect 17224 21684 17276 21690
rect 17224 21626 17276 21632
rect 17696 21622 17724 22918
rect 17684 21616 17736 21622
rect 17684 21558 17736 21564
rect 17316 21548 17368 21554
rect 17316 21490 17368 21496
rect 16856 20936 16908 20942
rect 16856 20878 16908 20884
rect 16868 20534 16896 20878
rect 17328 20806 17356 21490
rect 17788 20942 17816 25638
rect 17880 24954 17908 25842
rect 18064 25838 18092 27814
rect 18144 26784 18196 26790
rect 18144 26726 18196 26732
rect 18156 25906 18184 26726
rect 18144 25900 18196 25906
rect 18144 25842 18196 25848
rect 18052 25832 18104 25838
rect 18052 25774 18104 25780
rect 17868 24948 17920 24954
rect 17868 24890 17920 24896
rect 17868 24812 17920 24818
rect 17868 24754 17920 24760
rect 17880 23866 17908 24754
rect 17868 23860 17920 23866
rect 17868 23802 17920 23808
rect 18144 23520 18196 23526
rect 18144 23462 18196 23468
rect 18156 23118 18184 23462
rect 18144 23112 18196 23118
rect 18144 23054 18196 23060
rect 18144 21684 18196 21690
rect 18144 21626 18196 21632
rect 18052 21548 18104 21554
rect 18052 21490 18104 21496
rect 18064 20942 18092 21490
rect 18156 20942 18184 21626
rect 17776 20936 17828 20942
rect 17776 20878 17828 20884
rect 18052 20936 18104 20942
rect 18052 20878 18104 20884
rect 18144 20936 18196 20942
rect 18144 20878 18196 20884
rect 17316 20800 17368 20806
rect 17316 20742 17368 20748
rect 16856 20528 16908 20534
rect 16856 20470 16908 20476
rect 16672 19984 16724 19990
rect 16672 19926 16724 19932
rect 16488 19168 16540 19174
rect 16488 19110 16540 19116
rect 16500 18766 16528 19110
rect 16488 18760 16540 18766
rect 16488 18702 16540 18708
rect 16304 18692 16356 18698
rect 16304 18634 16356 18640
rect 16316 18426 16344 18634
rect 16304 18420 16356 18426
rect 16304 18362 16356 18368
rect 16316 17814 16344 18362
rect 16684 17882 16712 19926
rect 16868 19446 16896 20470
rect 17328 19786 17356 20742
rect 17684 20256 17736 20262
rect 17684 20198 17736 20204
rect 17408 19848 17460 19854
rect 17408 19790 17460 19796
rect 17316 19780 17368 19786
rect 17316 19722 17368 19728
rect 17420 19530 17448 19790
rect 17696 19786 17724 20198
rect 17684 19780 17736 19786
rect 17684 19722 17736 19728
rect 17420 19502 17540 19530
rect 16856 19440 16908 19446
rect 16856 19382 16908 19388
rect 17408 19440 17460 19446
rect 17408 19382 17460 19388
rect 16868 18272 16896 19382
rect 17316 19168 17368 19174
rect 17316 19110 17368 19116
rect 17328 18834 17356 19110
rect 17316 18828 17368 18834
rect 17316 18770 17368 18776
rect 16948 18284 17000 18290
rect 16868 18244 16948 18272
rect 16948 18226 17000 18232
rect 17420 18222 17448 19382
rect 17512 18970 17540 19502
rect 18064 19334 18092 20878
rect 17972 19306 18092 19334
rect 17868 19168 17920 19174
rect 17868 19110 17920 19116
rect 17500 18964 17552 18970
rect 17500 18906 17552 18912
rect 17776 18828 17828 18834
rect 17776 18770 17828 18776
rect 17408 18216 17460 18222
rect 17408 18158 17460 18164
rect 16672 17876 16724 17882
rect 16672 17818 16724 17824
rect 16304 17808 16356 17814
rect 16304 17750 16356 17756
rect 16120 16788 16172 16794
rect 16224 16782 16344 16810
rect 16120 16730 16172 16736
rect 16212 16448 16264 16454
rect 16212 16390 16264 16396
rect 16224 16114 16252 16390
rect 16028 16108 16080 16114
rect 16028 16050 16080 16056
rect 16212 16108 16264 16114
rect 16212 16050 16264 16056
rect 16224 15570 16252 16050
rect 16212 15564 16264 15570
rect 16212 15506 16264 15512
rect 16316 15434 16344 16782
rect 16488 15972 16540 15978
rect 16488 15914 16540 15920
rect 16304 15428 16356 15434
rect 16304 15370 16356 15376
rect 15672 15286 15884 15314
rect 15568 14408 15620 14414
rect 15568 14350 15620 14356
rect 15476 13932 15528 13938
rect 15476 13874 15528 13880
rect 15488 13326 15516 13874
rect 15568 13728 15620 13734
rect 15568 13670 15620 13676
rect 15476 13320 15528 13326
rect 15476 13262 15528 13268
rect 15384 13252 15436 13258
rect 15384 13194 15436 13200
rect 15580 13190 15608 13670
rect 15568 13184 15620 13190
rect 15568 13126 15620 13132
rect 15672 13002 15700 15286
rect 16500 14958 16528 15914
rect 16488 14952 16540 14958
rect 16488 14894 16540 14900
rect 16120 14408 16172 14414
rect 16120 14350 16172 14356
rect 15752 13184 15804 13190
rect 15752 13126 15804 13132
rect 15488 12974 15700 13002
rect 14740 12844 14792 12850
rect 14740 12786 14792 12792
rect 14846 12540 15154 12560
rect 14846 12538 14852 12540
rect 14908 12538 14932 12540
rect 14988 12538 15012 12540
rect 15068 12538 15092 12540
rect 15148 12538 15154 12540
rect 14908 12486 14910 12538
rect 15090 12486 15092 12538
rect 14846 12484 14852 12486
rect 14908 12484 14932 12486
rect 14988 12484 15012 12486
rect 15068 12484 15092 12486
rect 15148 12484 15154 12486
rect 14846 12464 15154 12484
rect 15488 11762 15516 12974
rect 15568 12844 15620 12850
rect 15568 12786 15620 12792
rect 15580 12442 15608 12786
rect 15568 12436 15620 12442
rect 15568 12378 15620 12384
rect 15764 12238 15792 13126
rect 16132 12986 16160 14350
rect 16684 14346 16712 17818
rect 17316 17536 17368 17542
rect 17316 17478 17368 17484
rect 16856 17196 16908 17202
rect 16856 17138 16908 17144
rect 16868 14618 16896 17138
rect 17328 16590 17356 17478
rect 17420 16794 17448 18158
rect 17408 16788 17460 16794
rect 17408 16730 17460 16736
rect 17592 16652 17644 16658
rect 17592 16594 17644 16600
rect 17316 16584 17368 16590
rect 17316 16526 17368 16532
rect 16856 14612 16908 14618
rect 16856 14554 16908 14560
rect 16672 14340 16724 14346
rect 16672 14282 16724 14288
rect 16684 14074 16712 14282
rect 16672 14068 16724 14074
rect 16672 14010 16724 14016
rect 16868 14006 16896 14554
rect 16856 14000 16908 14006
rect 16856 13942 16908 13948
rect 16868 13326 16896 13942
rect 17132 13728 17184 13734
rect 17132 13670 17184 13676
rect 17408 13728 17460 13734
rect 17408 13670 17460 13676
rect 16856 13320 16908 13326
rect 16856 13262 16908 13268
rect 16120 12980 16172 12986
rect 16120 12922 16172 12928
rect 17144 12782 17172 13670
rect 17224 13252 17276 13258
rect 17224 13194 17276 13200
rect 17316 13252 17368 13258
rect 17316 13194 17368 13200
rect 17132 12776 17184 12782
rect 17132 12718 17184 12724
rect 17236 12442 17264 13194
rect 17328 12918 17356 13194
rect 17316 12912 17368 12918
rect 17316 12854 17368 12860
rect 17224 12436 17276 12442
rect 17224 12378 17276 12384
rect 15752 12232 15804 12238
rect 15752 12174 15804 12180
rect 15476 11756 15528 11762
rect 15476 11698 15528 11704
rect 14846 11452 15154 11472
rect 14846 11450 14852 11452
rect 14908 11450 14932 11452
rect 14988 11450 15012 11452
rect 15068 11450 15092 11452
rect 15148 11450 15154 11452
rect 14908 11398 14910 11450
rect 15090 11398 15092 11450
rect 14846 11396 14852 11398
rect 14908 11396 14932 11398
rect 14988 11396 15012 11398
rect 15068 11396 15092 11398
rect 15148 11396 15154 11398
rect 14846 11376 15154 11396
rect 17328 11218 17356 12854
rect 17420 12238 17448 13670
rect 17604 13326 17632 16594
rect 17684 15904 17736 15910
rect 17684 15846 17736 15852
rect 17696 15638 17724 15846
rect 17684 15632 17736 15638
rect 17684 15574 17736 15580
rect 17592 13320 17644 13326
rect 17592 13262 17644 13268
rect 17408 12232 17460 12238
rect 17408 12174 17460 12180
rect 17592 11552 17644 11558
rect 17592 11494 17644 11500
rect 13820 11212 13872 11218
rect 13820 11154 13872 11160
rect 16948 11212 17000 11218
rect 16948 11154 17000 11160
rect 17316 11212 17368 11218
rect 17316 11154 17368 11160
rect 16580 11144 16632 11150
rect 16580 11086 16632 11092
rect 15568 11008 15620 11014
rect 15568 10950 15620 10956
rect 15936 11008 15988 11014
rect 15936 10950 15988 10956
rect 10214 10908 10522 10928
rect 10214 10906 10220 10908
rect 10276 10906 10300 10908
rect 10356 10906 10380 10908
rect 10436 10906 10460 10908
rect 10516 10906 10522 10908
rect 10276 10854 10278 10906
rect 10458 10854 10460 10906
rect 10214 10852 10220 10854
rect 10276 10852 10300 10854
rect 10356 10852 10380 10854
rect 10436 10852 10460 10854
rect 10516 10852 10522 10854
rect 10214 10832 10522 10852
rect 14846 10364 15154 10384
rect 14846 10362 14852 10364
rect 14908 10362 14932 10364
rect 14988 10362 15012 10364
rect 15068 10362 15092 10364
rect 15148 10362 15154 10364
rect 14908 10310 14910 10362
rect 15090 10310 15092 10362
rect 14846 10308 14852 10310
rect 14908 10308 14932 10310
rect 14988 10308 15012 10310
rect 15068 10308 15092 10310
rect 15148 10308 15154 10310
rect 14846 10288 15154 10308
rect 15580 10130 15608 10950
rect 15948 10674 15976 10950
rect 15936 10668 15988 10674
rect 15936 10610 15988 10616
rect 16592 10266 16620 11086
rect 16580 10260 16632 10266
rect 16580 10202 16632 10208
rect 15568 10124 15620 10130
rect 15568 10066 15620 10072
rect 10214 9820 10522 9840
rect 10214 9818 10220 9820
rect 10276 9818 10300 9820
rect 10356 9818 10380 9820
rect 10436 9818 10460 9820
rect 10516 9818 10522 9820
rect 10276 9766 10278 9818
rect 10458 9766 10460 9818
rect 10214 9764 10220 9766
rect 10276 9764 10300 9766
rect 10356 9764 10380 9766
rect 10436 9764 10460 9766
rect 10516 9764 10522 9766
rect 10214 9744 10522 9764
rect 14846 9276 15154 9296
rect 14846 9274 14852 9276
rect 14908 9274 14932 9276
rect 14988 9274 15012 9276
rect 15068 9274 15092 9276
rect 15148 9274 15154 9276
rect 14908 9222 14910 9274
rect 15090 9222 15092 9274
rect 14846 9220 14852 9222
rect 14908 9220 14932 9222
rect 14988 9220 15012 9222
rect 15068 9220 15092 9222
rect 15148 9220 15154 9222
rect 14846 9200 15154 9220
rect 10214 8732 10522 8752
rect 10214 8730 10220 8732
rect 10276 8730 10300 8732
rect 10356 8730 10380 8732
rect 10436 8730 10460 8732
rect 10516 8730 10522 8732
rect 10276 8678 10278 8730
rect 10458 8678 10460 8730
rect 10214 8676 10220 8678
rect 10276 8676 10300 8678
rect 10356 8676 10380 8678
rect 10436 8676 10460 8678
rect 10516 8676 10522 8678
rect 10214 8656 10522 8676
rect 14846 8188 15154 8208
rect 14846 8186 14852 8188
rect 14908 8186 14932 8188
rect 14988 8186 15012 8188
rect 15068 8186 15092 8188
rect 15148 8186 15154 8188
rect 14908 8134 14910 8186
rect 15090 8134 15092 8186
rect 14846 8132 14852 8134
rect 14908 8132 14932 8134
rect 14988 8132 15012 8134
rect 15068 8132 15092 8134
rect 15148 8132 15154 8134
rect 14846 8112 15154 8132
rect 10214 7644 10522 7664
rect 10214 7642 10220 7644
rect 10276 7642 10300 7644
rect 10356 7642 10380 7644
rect 10436 7642 10460 7644
rect 10516 7642 10522 7644
rect 10276 7590 10278 7642
rect 10458 7590 10460 7642
rect 10214 7588 10220 7590
rect 10276 7588 10300 7590
rect 10356 7588 10380 7590
rect 10436 7588 10460 7590
rect 10516 7588 10522 7590
rect 10214 7568 10522 7588
rect 14846 7100 15154 7120
rect 14846 7098 14852 7100
rect 14908 7098 14932 7100
rect 14988 7098 15012 7100
rect 15068 7098 15092 7100
rect 15148 7098 15154 7100
rect 14908 7046 14910 7098
rect 15090 7046 15092 7098
rect 14846 7044 14852 7046
rect 14908 7044 14932 7046
rect 14988 7044 15012 7046
rect 15068 7044 15092 7046
rect 15148 7044 15154 7046
rect 14846 7024 15154 7044
rect 10214 6556 10522 6576
rect 10214 6554 10220 6556
rect 10276 6554 10300 6556
rect 10356 6554 10380 6556
rect 10436 6554 10460 6556
rect 10516 6554 10522 6556
rect 10276 6502 10278 6554
rect 10458 6502 10460 6554
rect 10214 6500 10220 6502
rect 10276 6500 10300 6502
rect 10356 6500 10380 6502
rect 10436 6500 10460 6502
rect 10516 6500 10522 6502
rect 10214 6480 10522 6500
rect 14846 6012 15154 6032
rect 14846 6010 14852 6012
rect 14908 6010 14932 6012
rect 14988 6010 15012 6012
rect 15068 6010 15092 6012
rect 15148 6010 15154 6012
rect 14908 5958 14910 6010
rect 15090 5958 15092 6010
rect 14846 5956 14852 5958
rect 14908 5956 14932 5958
rect 14988 5956 15012 5958
rect 15068 5956 15092 5958
rect 15148 5956 15154 5958
rect 14846 5936 15154 5956
rect 10214 5468 10522 5488
rect 10214 5466 10220 5468
rect 10276 5466 10300 5468
rect 10356 5466 10380 5468
rect 10436 5466 10460 5468
rect 10516 5466 10522 5468
rect 10276 5414 10278 5466
rect 10458 5414 10460 5466
rect 10214 5412 10220 5414
rect 10276 5412 10300 5414
rect 10356 5412 10380 5414
rect 10436 5412 10460 5414
rect 10516 5412 10522 5414
rect 10214 5392 10522 5412
rect 14846 4924 15154 4944
rect 14846 4922 14852 4924
rect 14908 4922 14932 4924
rect 14988 4922 15012 4924
rect 15068 4922 15092 4924
rect 15148 4922 15154 4924
rect 14908 4870 14910 4922
rect 15090 4870 15092 4922
rect 14846 4868 14852 4870
rect 14908 4868 14932 4870
rect 14988 4868 15012 4870
rect 15068 4868 15092 4870
rect 15148 4868 15154 4870
rect 14846 4848 15154 4868
rect 10214 4380 10522 4400
rect 10214 4378 10220 4380
rect 10276 4378 10300 4380
rect 10356 4378 10380 4380
rect 10436 4378 10460 4380
rect 10516 4378 10522 4380
rect 10276 4326 10278 4378
rect 10458 4326 10460 4378
rect 10214 4324 10220 4326
rect 10276 4324 10300 4326
rect 10356 4324 10380 4326
rect 10436 4324 10460 4326
rect 10516 4324 10522 4326
rect 10214 4304 10522 4324
rect 12900 4140 12952 4146
rect 12900 4082 12952 4088
rect 12624 4072 12676 4078
rect 12624 4014 12676 4020
rect 11704 3936 11756 3942
rect 11704 3878 11756 3884
rect 9680 3596 9732 3602
rect 9680 3538 9732 3544
rect 9496 2644 9548 2650
rect 9496 2586 9548 2592
rect 9036 2372 9088 2378
rect 9036 2314 9088 2320
rect 9048 800 9076 2314
rect 9692 800 9720 3538
rect 11520 3528 11572 3534
rect 11520 3470 11572 3476
rect 10214 3292 10522 3312
rect 10214 3290 10220 3292
rect 10276 3290 10300 3292
rect 10356 3290 10380 3292
rect 10436 3290 10460 3292
rect 10516 3290 10522 3292
rect 10276 3238 10278 3290
rect 10458 3238 10460 3290
rect 10214 3236 10220 3238
rect 10276 3236 10300 3238
rect 10356 3236 10380 3238
rect 10436 3236 10460 3238
rect 10516 3236 10522 3238
rect 10214 3216 10522 3236
rect 11532 3058 11560 3470
rect 11716 3126 11744 3878
rect 12636 3738 12664 4014
rect 12912 3942 12940 4082
rect 13176 4072 13228 4078
rect 13176 4014 13228 4020
rect 13544 4072 13596 4078
rect 13544 4014 13596 4020
rect 12900 3936 12952 3942
rect 12900 3878 12952 3884
rect 13188 3738 13216 4014
rect 12624 3732 12676 3738
rect 12624 3674 12676 3680
rect 13176 3732 13228 3738
rect 13176 3674 13228 3680
rect 13084 3528 13136 3534
rect 13084 3470 13136 3476
rect 13096 3194 13124 3470
rect 13084 3188 13136 3194
rect 13084 3130 13136 3136
rect 11704 3120 11756 3126
rect 11704 3062 11756 3068
rect 11520 3052 11572 3058
rect 11520 2994 11572 3000
rect 10968 2916 11020 2922
rect 10968 2858 11020 2864
rect 10214 2204 10522 2224
rect 10214 2202 10220 2204
rect 10276 2202 10300 2204
rect 10356 2202 10380 2204
rect 10436 2202 10460 2204
rect 10516 2202 10522 2204
rect 10276 2150 10278 2202
rect 10458 2150 10460 2202
rect 10214 2148 10220 2150
rect 10276 2148 10300 2150
rect 10356 2148 10380 2150
rect 10436 2148 10460 2150
rect 10516 2148 10522 2150
rect 10214 2128 10522 2148
rect 10980 800 11008 2858
rect 13556 800 13584 4014
rect 14846 3836 15154 3856
rect 14846 3834 14852 3836
rect 14908 3834 14932 3836
rect 14988 3834 15012 3836
rect 15068 3834 15092 3836
rect 15148 3834 15154 3836
rect 14908 3782 14910 3834
rect 15090 3782 15092 3834
rect 14846 3780 14852 3782
rect 14908 3780 14932 3782
rect 14988 3780 15012 3782
rect 15068 3780 15092 3782
rect 15148 3780 15154 3782
rect 14846 3760 15154 3780
rect 14646 3632 14702 3641
rect 14646 3567 14702 3576
rect 14660 3534 14688 3567
rect 14648 3528 14700 3534
rect 14648 3470 14700 3476
rect 16304 3528 16356 3534
rect 16304 3470 16356 3476
rect 16672 3528 16724 3534
rect 16672 3470 16724 3476
rect 14280 3460 14332 3466
rect 14280 3402 14332 3408
rect 14292 3058 14320 3402
rect 14464 3392 14516 3398
rect 14464 3334 14516 3340
rect 14476 3126 14504 3334
rect 14464 3120 14516 3126
rect 14464 3062 14516 3068
rect 14280 3052 14332 3058
rect 14280 2994 14332 3000
rect 14740 2984 14792 2990
rect 14740 2926 14792 2932
rect 14752 1578 14780 2926
rect 16316 2854 16344 3470
rect 16684 3058 16712 3470
rect 16856 3392 16908 3398
rect 16856 3334 16908 3340
rect 16868 3126 16896 3334
rect 16856 3120 16908 3126
rect 16856 3062 16908 3068
rect 16672 3052 16724 3058
rect 16672 2994 16724 3000
rect 16764 2916 16816 2922
rect 16764 2858 16816 2864
rect 16028 2848 16080 2854
rect 16028 2790 16080 2796
rect 16304 2848 16356 2854
rect 16304 2790 16356 2796
rect 14846 2748 15154 2768
rect 14846 2746 14852 2748
rect 14908 2746 14932 2748
rect 14988 2746 15012 2748
rect 15068 2746 15092 2748
rect 15148 2746 15154 2748
rect 14908 2694 14910 2746
rect 15090 2694 15092 2746
rect 14846 2692 14852 2694
rect 14908 2692 14932 2694
rect 14988 2692 15012 2694
rect 15068 2692 15092 2694
rect 15148 2692 15154 2694
rect 14846 2672 15154 2692
rect 16040 2446 16068 2790
rect 16028 2440 16080 2446
rect 16028 2382 16080 2388
rect 16120 2440 16172 2446
rect 16120 2382 16172 2388
rect 14752 1550 14872 1578
rect 14844 800 14872 1550
rect 16132 800 16160 2382
rect 16776 800 16804 2858
rect 16960 2774 16988 11154
rect 17328 10742 17356 11154
rect 17604 11150 17632 11494
rect 17592 11144 17644 11150
rect 17592 11086 17644 11092
rect 17696 10810 17724 15574
rect 17788 13938 17816 18770
rect 17880 18290 17908 19110
rect 17868 18284 17920 18290
rect 17868 18226 17920 18232
rect 17880 16658 17908 18226
rect 17972 16998 18000 19306
rect 18156 18986 18184 20878
rect 18064 18958 18184 18986
rect 18064 17542 18092 18958
rect 18052 17536 18104 17542
rect 18052 17478 18104 17484
rect 17960 16992 18012 16998
rect 17960 16934 18012 16940
rect 17868 16652 17920 16658
rect 17868 16594 17920 16600
rect 18064 16250 18092 17478
rect 18144 17128 18196 17134
rect 18144 17070 18196 17076
rect 18156 16794 18184 17070
rect 18144 16788 18196 16794
rect 18144 16730 18196 16736
rect 18052 16244 18104 16250
rect 18052 16186 18104 16192
rect 17868 14068 17920 14074
rect 17868 14010 17920 14016
rect 17776 13932 17828 13938
rect 17776 13874 17828 13880
rect 17788 12850 17816 13874
rect 17776 12844 17828 12850
rect 17776 12786 17828 12792
rect 17880 11762 17908 14010
rect 17868 11756 17920 11762
rect 17868 11698 17920 11704
rect 17684 10804 17736 10810
rect 17684 10746 17736 10752
rect 17316 10736 17368 10742
rect 17316 10678 17368 10684
rect 17696 10062 17724 10746
rect 17684 10056 17736 10062
rect 17684 9998 17736 10004
rect 17500 9920 17552 9926
rect 17500 9862 17552 9868
rect 16868 2746 16988 2774
rect 16868 2650 16896 2746
rect 17512 2650 17540 9862
rect 17684 5024 17736 5030
rect 17684 4966 17736 4972
rect 17696 4554 17724 4966
rect 17684 4548 17736 4554
rect 17684 4490 17736 4496
rect 18248 4078 18276 35550
rect 18326 35184 18382 35193
rect 18326 35119 18328 35128
rect 18380 35119 18382 35128
rect 18328 35090 18380 35096
rect 18328 33584 18380 33590
rect 18328 33526 18380 33532
rect 18340 32502 18368 33526
rect 18328 32496 18380 32502
rect 18328 32438 18380 32444
rect 18340 31346 18368 32438
rect 18328 31340 18380 31346
rect 18328 31282 18380 31288
rect 18328 27872 18380 27878
rect 18328 27814 18380 27820
rect 18340 26994 18368 27814
rect 18328 26988 18380 26994
rect 18328 26930 18380 26936
rect 18340 26586 18368 26930
rect 18432 26874 18460 36654
rect 18696 35760 18748 35766
rect 18696 35702 18748 35708
rect 18512 31680 18564 31686
rect 18512 31622 18564 31628
rect 18524 31414 18552 31622
rect 18512 31408 18564 31414
rect 18512 31350 18564 31356
rect 18512 28416 18564 28422
rect 18512 28358 18564 28364
rect 18524 28082 18552 28358
rect 18512 28076 18564 28082
rect 18512 28018 18564 28024
rect 18604 28076 18656 28082
rect 18604 28018 18656 28024
rect 18616 26994 18644 28018
rect 18708 27130 18736 35702
rect 18800 35698 18828 38286
rect 19260 37890 19288 39086
rect 19340 38956 19392 38962
rect 19340 38898 19392 38904
rect 19892 38956 19944 38962
rect 19892 38898 19944 38904
rect 19352 38010 19380 38898
rect 19524 38752 19576 38758
rect 19524 38694 19576 38700
rect 19536 38350 19564 38694
rect 19524 38344 19576 38350
rect 19524 38286 19576 38292
rect 19478 38108 19786 38128
rect 19478 38106 19484 38108
rect 19540 38106 19564 38108
rect 19620 38106 19644 38108
rect 19700 38106 19724 38108
rect 19780 38106 19786 38108
rect 19540 38054 19542 38106
rect 19722 38054 19724 38106
rect 19478 38052 19484 38054
rect 19540 38052 19564 38054
rect 19620 38052 19644 38054
rect 19700 38052 19724 38054
rect 19780 38052 19786 38054
rect 19478 38032 19786 38052
rect 19340 38004 19392 38010
rect 19340 37946 19392 37952
rect 19260 37862 19380 37890
rect 19352 36106 19380 37862
rect 19904 37466 19932 38898
rect 20168 37868 20220 37874
rect 20220 37828 20300 37856
rect 20168 37810 20220 37816
rect 20076 37800 20128 37806
rect 20076 37742 20128 37748
rect 19892 37460 19944 37466
rect 19892 37402 19944 37408
rect 19478 37020 19786 37040
rect 19478 37018 19484 37020
rect 19540 37018 19564 37020
rect 19620 37018 19644 37020
rect 19700 37018 19724 37020
rect 19780 37018 19786 37020
rect 19540 36966 19542 37018
rect 19722 36966 19724 37018
rect 19478 36964 19484 36966
rect 19540 36964 19564 36966
rect 19620 36964 19644 36966
rect 19700 36964 19724 36966
rect 19780 36964 19786 36966
rect 19478 36944 19786 36964
rect 20088 36378 20116 37742
rect 20168 37256 20220 37262
rect 20168 37198 20220 37204
rect 20076 36372 20128 36378
rect 20076 36314 20128 36320
rect 19340 36100 19392 36106
rect 19340 36042 19392 36048
rect 19892 36100 19944 36106
rect 19892 36042 19944 36048
rect 19478 35932 19786 35952
rect 19478 35930 19484 35932
rect 19540 35930 19564 35932
rect 19620 35930 19644 35932
rect 19700 35930 19724 35932
rect 19780 35930 19786 35932
rect 19540 35878 19542 35930
rect 19722 35878 19724 35930
rect 19478 35876 19484 35878
rect 19540 35876 19564 35878
rect 19620 35876 19644 35878
rect 19700 35876 19724 35878
rect 19780 35876 19786 35878
rect 19478 35856 19786 35876
rect 18788 35692 18840 35698
rect 18788 35634 18840 35640
rect 19340 35692 19392 35698
rect 19340 35634 19392 35640
rect 18800 33590 18828 35634
rect 18788 33584 18840 33590
rect 18788 33526 18840 33532
rect 19352 33114 19380 35634
rect 19904 34950 19932 36042
rect 19892 34944 19944 34950
rect 19892 34886 19944 34892
rect 19478 34844 19786 34864
rect 19478 34842 19484 34844
rect 19540 34842 19564 34844
rect 19620 34842 19644 34844
rect 19700 34842 19724 34844
rect 19780 34842 19786 34844
rect 19540 34790 19542 34842
rect 19722 34790 19724 34842
rect 19478 34788 19484 34790
rect 19540 34788 19564 34790
rect 19620 34788 19644 34790
rect 19700 34788 19724 34790
rect 19780 34788 19786 34790
rect 19478 34768 19786 34788
rect 19904 34610 19932 34886
rect 19892 34604 19944 34610
rect 19892 34546 19944 34552
rect 20180 34202 20208 37198
rect 20272 37126 20300 37828
rect 20352 37800 20404 37806
rect 20352 37742 20404 37748
rect 20260 37120 20312 37126
rect 20260 37062 20312 37068
rect 20168 34196 20220 34202
rect 20168 34138 20220 34144
rect 19892 33924 19944 33930
rect 19892 33866 19944 33872
rect 19478 33756 19786 33776
rect 19478 33754 19484 33756
rect 19540 33754 19564 33756
rect 19620 33754 19644 33756
rect 19700 33754 19724 33756
rect 19780 33754 19786 33756
rect 19540 33702 19542 33754
rect 19722 33702 19724 33754
rect 19478 33700 19484 33702
rect 19540 33700 19564 33702
rect 19620 33700 19644 33702
rect 19700 33700 19724 33702
rect 19780 33700 19786 33702
rect 19478 33680 19786 33700
rect 19904 33522 19932 33866
rect 20168 33856 20220 33862
rect 20168 33798 20220 33804
rect 20180 33522 20208 33798
rect 19892 33516 19944 33522
rect 19892 33458 19944 33464
rect 20168 33516 20220 33522
rect 20168 33458 20220 33464
rect 19340 33108 19392 33114
rect 19340 33050 19392 33056
rect 19478 32668 19786 32688
rect 19478 32666 19484 32668
rect 19540 32666 19564 32668
rect 19620 32666 19644 32668
rect 19700 32666 19724 32668
rect 19780 32666 19786 32668
rect 19540 32614 19542 32666
rect 19722 32614 19724 32666
rect 19478 32612 19484 32614
rect 19540 32612 19564 32614
rect 19620 32612 19644 32614
rect 19700 32612 19724 32614
rect 19780 32612 19786 32614
rect 19478 32592 19786 32612
rect 19616 32224 19668 32230
rect 19616 32166 19668 32172
rect 19628 31822 19656 32166
rect 19616 31816 19668 31822
rect 19616 31758 19668 31764
rect 19478 31580 19786 31600
rect 19478 31578 19484 31580
rect 19540 31578 19564 31580
rect 19620 31578 19644 31580
rect 19700 31578 19724 31580
rect 19780 31578 19786 31580
rect 19540 31526 19542 31578
rect 19722 31526 19724 31578
rect 19478 31524 19484 31526
rect 19540 31524 19564 31526
rect 19620 31524 19644 31526
rect 19700 31524 19724 31526
rect 19780 31524 19786 31526
rect 19478 31504 19786 31524
rect 19248 31136 19300 31142
rect 19248 31078 19300 31084
rect 19260 30666 19288 31078
rect 19340 30864 19392 30870
rect 19340 30806 19392 30812
rect 19248 30660 19300 30666
rect 19248 30602 19300 30608
rect 18972 30184 19024 30190
rect 18972 30126 19024 30132
rect 18788 27872 18840 27878
rect 18788 27814 18840 27820
rect 18696 27124 18748 27130
rect 18696 27066 18748 27072
rect 18604 26988 18656 26994
rect 18604 26930 18656 26936
rect 18432 26846 18644 26874
rect 18328 26580 18380 26586
rect 18328 26522 18380 26528
rect 18512 26308 18564 26314
rect 18512 26250 18564 26256
rect 18420 23248 18472 23254
rect 18420 23190 18472 23196
rect 18432 21690 18460 23190
rect 18420 21684 18472 21690
rect 18420 21626 18472 21632
rect 18524 21434 18552 26250
rect 18432 21406 18552 21434
rect 18432 20602 18460 21406
rect 18512 21344 18564 21350
rect 18512 21286 18564 21292
rect 18524 21010 18552 21286
rect 18512 21004 18564 21010
rect 18512 20946 18564 20952
rect 18420 20596 18472 20602
rect 18420 20538 18472 20544
rect 18432 19938 18460 20538
rect 18524 20466 18552 20946
rect 18512 20460 18564 20466
rect 18512 20402 18564 20408
rect 18340 19910 18460 19938
rect 18340 19854 18368 19910
rect 18328 19848 18380 19854
rect 18328 19790 18380 19796
rect 18328 18624 18380 18630
rect 18328 18566 18380 18572
rect 18340 18358 18368 18566
rect 18328 18352 18380 18358
rect 18328 18294 18380 18300
rect 18328 18080 18380 18086
rect 18328 18022 18380 18028
rect 18340 17678 18368 18022
rect 18328 17672 18380 17678
rect 18328 17614 18380 17620
rect 18328 15496 18380 15502
rect 18328 15438 18380 15444
rect 18420 15496 18472 15502
rect 18420 15438 18472 15444
rect 18340 15162 18368 15438
rect 18328 15156 18380 15162
rect 18328 15098 18380 15104
rect 18328 13932 18380 13938
rect 18328 13874 18380 13880
rect 18340 13190 18368 13874
rect 18328 13184 18380 13190
rect 18328 13126 18380 13132
rect 18340 12918 18368 13126
rect 18328 12912 18380 12918
rect 18328 12854 18380 12860
rect 18432 11898 18460 15438
rect 18420 11892 18472 11898
rect 18420 11834 18472 11840
rect 18616 5710 18644 26846
rect 18800 25974 18828 27814
rect 18984 25974 19012 30126
rect 19064 30116 19116 30122
rect 19064 30058 19116 30064
rect 19076 29306 19104 30058
rect 19260 29646 19288 30602
rect 19352 30258 19380 30806
rect 19478 30492 19786 30512
rect 19478 30490 19484 30492
rect 19540 30490 19564 30492
rect 19620 30490 19644 30492
rect 19700 30490 19724 30492
rect 19780 30490 19786 30492
rect 19540 30438 19542 30490
rect 19722 30438 19724 30490
rect 19478 30436 19484 30438
rect 19540 30436 19564 30438
rect 19620 30436 19644 30438
rect 19700 30436 19724 30438
rect 19780 30436 19786 30438
rect 19478 30416 19786 30436
rect 19340 30252 19392 30258
rect 19340 30194 19392 30200
rect 19800 30252 19852 30258
rect 19800 30194 19852 30200
rect 19340 30048 19392 30054
rect 19340 29990 19392 29996
rect 19352 29646 19380 29990
rect 19812 29646 19840 30194
rect 19248 29640 19300 29646
rect 19248 29582 19300 29588
rect 19340 29640 19392 29646
rect 19340 29582 19392 29588
rect 19800 29640 19852 29646
rect 19800 29582 19852 29588
rect 19478 29404 19786 29424
rect 19478 29402 19484 29404
rect 19540 29402 19564 29404
rect 19620 29402 19644 29404
rect 19700 29402 19724 29404
rect 19780 29402 19786 29404
rect 19540 29350 19542 29402
rect 19722 29350 19724 29402
rect 19478 29348 19484 29350
rect 19540 29348 19564 29350
rect 19620 29348 19644 29350
rect 19700 29348 19724 29350
rect 19780 29348 19786 29350
rect 19478 29328 19786 29348
rect 19064 29300 19116 29306
rect 19064 29242 19116 29248
rect 19478 28316 19786 28336
rect 19478 28314 19484 28316
rect 19540 28314 19564 28316
rect 19620 28314 19644 28316
rect 19700 28314 19724 28316
rect 19780 28314 19786 28316
rect 19540 28262 19542 28314
rect 19722 28262 19724 28314
rect 19478 28260 19484 28262
rect 19540 28260 19564 28262
rect 19620 28260 19644 28262
rect 19700 28260 19724 28262
rect 19780 28260 19786 28262
rect 19478 28240 19786 28260
rect 19248 27872 19300 27878
rect 19248 27814 19300 27820
rect 19156 26988 19208 26994
rect 19156 26930 19208 26936
rect 19064 26512 19116 26518
rect 19064 26454 19116 26460
rect 18788 25968 18840 25974
rect 18788 25910 18840 25916
rect 18972 25968 19024 25974
rect 18972 25910 19024 25916
rect 18800 23050 18828 25910
rect 19076 25906 19104 26454
rect 19168 26042 19196 26930
rect 19260 26382 19288 27814
rect 19478 27228 19786 27248
rect 19478 27226 19484 27228
rect 19540 27226 19564 27228
rect 19620 27226 19644 27228
rect 19700 27226 19724 27228
rect 19780 27226 19786 27228
rect 19540 27174 19542 27226
rect 19722 27174 19724 27226
rect 19478 27172 19484 27174
rect 19540 27172 19564 27174
rect 19620 27172 19644 27174
rect 19700 27172 19724 27174
rect 19780 27172 19786 27174
rect 19478 27152 19786 27172
rect 19904 26382 19932 33458
rect 19984 33312 20036 33318
rect 19984 33254 20036 33260
rect 19996 33046 20024 33254
rect 19984 33040 20036 33046
rect 19984 32982 20036 32988
rect 19996 32450 20024 32982
rect 20168 32904 20220 32910
rect 20168 32846 20220 32852
rect 20180 32570 20208 32846
rect 20168 32564 20220 32570
rect 20168 32506 20220 32512
rect 20272 32502 20300 37062
rect 20260 32496 20312 32502
rect 19996 32434 20116 32450
rect 20260 32438 20312 32444
rect 19996 32428 20128 32434
rect 19996 32422 20076 32428
rect 20076 32370 20128 32376
rect 20088 32042 20116 32370
rect 20088 32014 20208 32042
rect 20076 31816 20128 31822
rect 20076 31758 20128 31764
rect 20088 31142 20116 31758
rect 20180 31346 20208 32014
rect 20168 31340 20220 31346
rect 20168 31282 20220 31288
rect 20076 31136 20128 31142
rect 20076 31078 20128 31084
rect 19984 30660 20036 30666
rect 19984 30602 20036 30608
rect 19996 30394 20024 30602
rect 19984 30388 20036 30394
rect 19984 30330 20036 30336
rect 19248 26376 19300 26382
rect 19248 26318 19300 26324
rect 19892 26376 19944 26382
rect 19892 26318 19944 26324
rect 19478 26140 19786 26160
rect 19478 26138 19484 26140
rect 19540 26138 19564 26140
rect 19620 26138 19644 26140
rect 19700 26138 19724 26140
rect 19780 26138 19786 26140
rect 19540 26086 19542 26138
rect 19722 26086 19724 26138
rect 19478 26084 19484 26086
rect 19540 26084 19564 26086
rect 19620 26084 19644 26086
rect 19700 26084 19724 26086
rect 19780 26084 19786 26086
rect 19478 26064 19786 26084
rect 19156 26036 19208 26042
rect 19156 25978 19208 25984
rect 19064 25900 19116 25906
rect 19064 25842 19116 25848
rect 19340 25900 19392 25906
rect 19340 25842 19392 25848
rect 18880 24608 18932 24614
rect 18880 24550 18932 24556
rect 18892 23050 18920 24550
rect 19064 24200 19116 24206
rect 19064 24142 19116 24148
rect 18972 23112 19024 23118
rect 18972 23054 19024 23060
rect 18788 23044 18840 23050
rect 18788 22986 18840 22992
rect 18880 23044 18932 23050
rect 18880 22986 18932 22992
rect 18892 22642 18920 22986
rect 18984 22778 19012 23054
rect 18972 22772 19024 22778
rect 18972 22714 19024 22720
rect 18880 22636 18932 22642
rect 18880 22578 18932 22584
rect 18972 22636 19024 22642
rect 18972 22578 19024 22584
rect 18984 21350 19012 22578
rect 19076 21622 19104 24142
rect 19352 21690 19380 25842
rect 19478 25052 19786 25072
rect 19478 25050 19484 25052
rect 19540 25050 19564 25052
rect 19620 25050 19644 25052
rect 19700 25050 19724 25052
rect 19780 25050 19786 25052
rect 19540 24998 19542 25050
rect 19722 24998 19724 25050
rect 19478 24996 19484 24998
rect 19540 24996 19564 24998
rect 19620 24996 19644 24998
rect 19700 24996 19724 24998
rect 19780 24996 19786 24998
rect 19478 24976 19786 24996
rect 19904 24410 19932 26318
rect 19996 24614 20024 30330
rect 20088 27606 20116 31078
rect 20180 30258 20208 31282
rect 20260 30660 20312 30666
rect 20260 30602 20312 30608
rect 20272 30258 20300 30602
rect 20168 30252 20220 30258
rect 20168 30194 20220 30200
rect 20260 30252 20312 30258
rect 20260 30194 20312 30200
rect 20180 29850 20208 30194
rect 20168 29844 20220 29850
rect 20168 29786 20220 29792
rect 20168 29504 20220 29510
rect 20272 29492 20300 30194
rect 20220 29464 20300 29492
rect 20168 29446 20220 29452
rect 20180 28082 20208 29446
rect 20168 28076 20220 28082
rect 20168 28018 20220 28024
rect 20076 27600 20128 27606
rect 20076 27542 20128 27548
rect 20168 27464 20220 27470
rect 20168 27406 20220 27412
rect 20180 27130 20208 27406
rect 20364 27334 20392 37742
rect 20456 34678 20484 45426
rect 21928 45082 21956 46990
rect 22008 46368 22060 46374
rect 22008 46310 22060 46316
rect 22020 46034 22048 46310
rect 22572 46034 22600 49200
rect 23216 47122 23244 49200
rect 23204 47116 23256 47122
rect 23204 47058 23256 47064
rect 22744 46980 22796 46986
rect 22744 46922 22796 46928
rect 22008 46028 22060 46034
rect 22008 45970 22060 45976
rect 22560 46028 22612 46034
rect 22560 45970 22612 45976
rect 22192 45892 22244 45898
rect 22192 45834 22244 45840
rect 22204 45626 22232 45834
rect 22192 45620 22244 45626
rect 22192 45562 22244 45568
rect 22756 45558 22784 46922
rect 23860 46714 23888 49200
rect 26146 49056 26202 49065
rect 26146 48991 26202 49000
rect 25594 47696 25650 47705
rect 25594 47631 25650 47640
rect 24110 47356 24418 47376
rect 24110 47354 24116 47356
rect 24172 47354 24196 47356
rect 24252 47354 24276 47356
rect 24332 47354 24356 47356
rect 24412 47354 24418 47356
rect 24172 47302 24174 47354
rect 24354 47302 24356 47354
rect 24110 47300 24116 47302
rect 24172 47300 24196 47302
rect 24252 47300 24276 47302
rect 24332 47300 24356 47302
rect 24412 47300 24418 47302
rect 24110 47280 24418 47300
rect 23848 46708 23900 46714
rect 23848 46650 23900 46656
rect 25608 46646 25636 47631
rect 25596 46640 25648 46646
rect 25596 46582 25648 46588
rect 23756 46504 23808 46510
rect 23756 46446 23808 46452
rect 23940 46504 23992 46510
rect 23940 46446 23992 46452
rect 23768 46170 23796 46446
rect 23756 46164 23808 46170
rect 23756 46106 23808 46112
rect 23952 45558 23980 46446
rect 25962 46336 26018 46345
rect 24110 46268 24418 46288
rect 25962 46271 26018 46280
rect 24110 46266 24116 46268
rect 24172 46266 24196 46268
rect 24252 46266 24276 46268
rect 24332 46266 24356 46268
rect 24412 46266 24418 46268
rect 24172 46214 24174 46266
rect 24354 46214 24356 46266
rect 24110 46212 24116 46214
rect 24172 46212 24196 46214
rect 24252 46212 24276 46214
rect 24332 46212 24356 46214
rect 24412 46212 24418 46214
rect 24110 46192 24418 46212
rect 25780 45960 25832 45966
rect 25780 45902 25832 45908
rect 22744 45552 22796 45558
rect 22744 45494 22796 45500
rect 23940 45552 23992 45558
rect 23940 45494 23992 45500
rect 22008 45484 22060 45490
rect 22008 45426 22060 45432
rect 23296 45484 23348 45490
rect 23296 45426 23348 45432
rect 21916 45076 21968 45082
rect 21916 45018 21968 45024
rect 22020 44305 22048 45426
rect 22006 44296 22062 44305
rect 22006 44231 22062 44240
rect 21824 39568 21876 39574
rect 21824 39510 21876 39516
rect 20812 39432 20864 39438
rect 20812 39374 20864 39380
rect 21180 39432 21232 39438
rect 21180 39374 21232 39380
rect 21272 39432 21324 39438
rect 21272 39374 21324 39380
rect 20536 39296 20588 39302
rect 20536 39238 20588 39244
rect 20548 38350 20576 39238
rect 20824 39030 20852 39374
rect 20904 39296 20956 39302
rect 20904 39238 20956 39244
rect 20812 39024 20864 39030
rect 20812 38966 20864 38972
rect 20824 38842 20852 38966
rect 20732 38814 20852 38842
rect 20536 38344 20588 38350
rect 20536 38286 20588 38292
rect 20548 37942 20576 38286
rect 20536 37936 20588 37942
rect 20536 37878 20588 37884
rect 20548 37738 20576 37878
rect 20536 37732 20588 37738
rect 20536 37674 20588 37680
rect 20548 37194 20576 37674
rect 20536 37188 20588 37194
rect 20536 37130 20588 37136
rect 20732 36174 20760 38814
rect 20812 38752 20864 38758
rect 20812 38694 20864 38700
rect 20824 38418 20852 38694
rect 20812 38412 20864 38418
rect 20812 38354 20864 38360
rect 20812 37664 20864 37670
rect 20812 37606 20864 37612
rect 20720 36168 20772 36174
rect 20720 36110 20772 36116
rect 20732 35766 20760 36110
rect 20720 35760 20772 35766
rect 20720 35702 20772 35708
rect 20720 35284 20772 35290
rect 20720 35226 20772 35232
rect 20444 34672 20496 34678
rect 20444 34614 20496 34620
rect 20628 34536 20680 34542
rect 20628 34478 20680 34484
rect 20444 34128 20496 34134
rect 20444 34070 20496 34076
rect 20456 31822 20484 34070
rect 20536 33924 20588 33930
rect 20536 33866 20588 33872
rect 20548 33386 20576 33866
rect 20536 33380 20588 33386
rect 20536 33322 20588 33328
rect 20548 31958 20576 33322
rect 20640 33046 20668 34478
rect 20732 33998 20760 35226
rect 20720 33992 20772 33998
rect 20720 33934 20772 33940
rect 20628 33040 20680 33046
rect 20628 32982 20680 32988
rect 20720 32836 20772 32842
rect 20720 32778 20772 32784
rect 20732 32366 20760 32778
rect 20720 32360 20772 32366
rect 20720 32302 20772 32308
rect 20536 31952 20588 31958
rect 20536 31894 20588 31900
rect 20732 31890 20760 32302
rect 20720 31884 20772 31890
rect 20720 31826 20772 31832
rect 20444 31816 20496 31822
rect 20444 31758 20496 31764
rect 20456 29646 20484 31758
rect 20444 29640 20496 29646
rect 20444 29582 20496 29588
rect 20732 28218 20760 31826
rect 20824 30734 20852 37606
rect 20916 37262 20944 39238
rect 20996 38820 21048 38826
rect 20996 38762 21048 38768
rect 20904 37256 20956 37262
rect 20904 37198 20956 37204
rect 21008 37126 21036 38762
rect 21192 38010 21220 39374
rect 21284 38894 21312 39374
rect 21836 38962 21864 39510
rect 21824 38956 21876 38962
rect 21824 38898 21876 38904
rect 22376 38956 22428 38962
rect 22376 38898 22428 38904
rect 21272 38888 21324 38894
rect 21272 38830 21324 38836
rect 22100 38888 22152 38894
rect 22100 38830 22152 38836
rect 21180 38004 21232 38010
rect 21180 37946 21232 37952
rect 20996 37120 21048 37126
rect 20996 37062 21048 37068
rect 20904 36168 20956 36174
rect 20904 36110 20956 36116
rect 20916 35034 20944 36110
rect 20996 36100 21048 36106
rect 20996 36042 21048 36048
rect 21008 35834 21036 36042
rect 20996 35828 21048 35834
rect 20996 35770 21048 35776
rect 21008 35680 21036 35770
rect 21088 35692 21140 35698
rect 21008 35652 21088 35680
rect 21008 35154 21036 35652
rect 21088 35634 21140 35640
rect 21192 35290 21220 37946
rect 21284 37942 21312 38830
rect 21364 38752 21416 38758
rect 21364 38694 21416 38700
rect 21272 37936 21324 37942
rect 21272 37878 21324 37884
rect 21272 36032 21324 36038
rect 21272 35974 21324 35980
rect 21180 35284 21232 35290
rect 21180 35226 21232 35232
rect 20996 35148 21048 35154
rect 20996 35090 21048 35096
rect 20916 35006 21036 35034
rect 21284 35018 21312 35974
rect 21008 34678 21036 35006
rect 21272 35012 21324 35018
rect 21272 34954 21324 34960
rect 21088 34944 21140 34950
rect 21088 34886 21140 34892
rect 21100 34678 21128 34886
rect 21284 34678 21312 34954
rect 20996 34672 21048 34678
rect 20996 34614 21048 34620
rect 21088 34672 21140 34678
rect 21088 34614 21140 34620
rect 21272 34672 21324 34678
rect 21272 34614 21324 34620
rect 20904 34604 20956 34610
rect 20904 34546 20956 34552
rect 20916 34202 20944 34546
rect 20904 34196 20956 34202
rect 20904 34138 20956 34144
rect 20916 33862 20944 34138
rect 20904 33856 20956 33862
rect 20904 33798 20956 33804
rect 20904 30864 20956 30870
rect 20904 30806 20956 30812
rect 20812 30728 20864 30734
rect 20812 30670 20864 30676
rect 20812 30252 20864 30258
rect 20916 30240 20944 30806
rect 20864 30212 20944 30240
rect 20812 30194 20864 30200
rect 20812 30116 20864 30122
rect 20812 30058 20864 30064
rect 20824 29782 20852 30058
rect 20812 29776 20864 29782
rect 20812 29718 20864 29724
rect 20720 28212 20772 28218
rect 20720 28154 20772 28160
rect 20536 28076 20588 28082
rect 20536 28018 20588 28024
rect 20548 27538 20576 28018
rect 20732 27538 20760 28154
rect 20824 28082 20852 29718
rect 21008 29714 21036 34614
rect 21284 34066 21312 34614
rect 21088 34060 21140 34066
rect 21088 34002 21140 34008
rect 21272 34060 21324 34066
rect 21272 34002 21324 34008
rect 21100 32434 21128 34002
rect 21088 32428 21140 32434
rect 21088 32370 21140 32376
rect 21180 32428 21232 32434
rect 21180 32370 21232 32376
rect 20996 29708 21048 29714
rect 20996 29650 21048 29656
rect 20812 28076 20864 28082
rect 20812 28018 20864 28024
rect 20536 27532 20588 27538
rect 20536 27474 20588 27480
rect 20720 27532 20772 27538
rect 20720 27474 20772 27480
rect 20444 27464 20496 27470
rect 20444 27406 20496 27412
rect 20352 27328 20404 27334
rect 20352 27270 20404 27276
rect 20168 27124 20220 27130
rect 20168 27066 20220 27072
rect 20364 26382 20392 27270
rect 20352 26376 20404 26382
rect 20352 26318 20404 26324
rect 20456 26314 20484 27406
rect 20444 26308 20496 26314
rect 20444 26250 20496 26256
rect 19984 24608 20036 24614
rect 19984 24550 20036 24556
rect 19892 24404 19944 24410
rect 19892 24346 19944 24352
rect 19478 23964 19786 23984
rect 19478 23962 19484 23964
rect 19540 23962 19564 23964
rect 19620 23962 19644 23964
rect 19700 23962 19724 23964
rect 19780 23962 19786 23964
rect 19540 23910 19542 23962
rect 19722 23910 19724 23962
rect 19478 23908 19484 23910
rect 19540 23908 19564 23910
rect 19620 23908 19644 23910
rect 19700 23908 19724 23910
rect 19780 23908 19786 23910
rect 19478 23888 19786 23908
rect 19800 23724 19852 23730
rect 19800 23666 19852 23672
rect 19812 23322 19840 23666
rect 19800 23316 19852 23322
rect 19800 23258 19852 23264
rect 19478 22876 19786 22896
rect 19478 22874 19484 22876
rect 19540 22874 19564 22876
rect 19620 22874 19644 22876
rect 19700 22874 19724 22876
rect 19780 22874 19786 22876
rect 19540 22822 19542 22874
rect 19722 22822 19724 22874
rect 19478 22820 19484 22822
rect 19540 22820 19564 22822
rect 19620 22820 19644 22822
rect 19700 22820 19724 22822
rect 19780 22820 19786 22822
rect 19478 22800 19786 22820
rect 19478 21788 19786 21808
rect 19478 21786 19484 21788
rect 19540 21786 19564 21788
rect 19620 21786 19644 21788
rect 19700 21786 19724 21788
rect 19780 21786 19786 21788
rect 19540 21734 19542 21786
rect 19722 21734 19724 21786
rect 19478 21732 19484 21734
rect 19540 21732 19564 21734
rect 19620 21732 19644 21734
rect 19700 21732 19724 21734
rect 19780 21732 19786 21734
rect 19478 21712 19786 21732
rect 19340 21684 19392 21690
rect 19340 21626 19392 21632
rect 19064 21616 19116 21622
rect 19064 21558 19116 21564
rect 18972 21344 19024 21350
rect 18972 21286 19024 21292
rect 18788 20936 18840 20942
rect 18788 20878 18840 20884
rect 18696 20868 18748 20874
rect 18696 20810 18748 20816
rect 18708 20602 18736 20810
rect 18696 20596 18748 20602
rect 18696 20538 18748 20544
rect 18800 20466 18828 20878
rect 18788 20460 18840 20466
rect 18788 20402 18840 20408
rect 18800 17882 18828 20402
rect 18984 19990 19012 21286
rect 19076 21146 19104 21558
rect 19064 21140 19116 21146
rect 19064 21082 19116 21088
rect 19478 20700 19786 20720
rect 19478 20698 19484 20700
rect 19540 20698 19564 20700
rect 19620 20698 19644 20700
rect 19700 20698 19724 20700
rect 19780 20698 19786 20700
rect 19540 20646 19542 20698
rect 19722 20646 19724 20698
rect 19478 20644 19484 20646
rect 19540 20644 19564 20646
rect 19620 20644 19644 20646
rect 19700 20644 19724 20646
rect 19780 20644 19786 20646
rect 19478 20624 19786 20644
rect 18972 19984 19024 19990
rect 18972 19926 19024 19932
rect 19478 19612 19786 19632
rect 19478 19610 19484 19612
rect 19540 19610 19564 19612
rect 19620 19610 19644 19612
rect 19700 19610 19724 19612
rect 19780 19610 19786 19612
rect 19540 19558 19542 19610
rect 19722 19558 19724 19610
rect 19478 19556 19484 19558
rect 19540 19556 19564 19558
rect 19620 19556 19644 19558
rect 19700 19556 19724 19558
rect 19780 19556 19786 19558
rect 19478 19536 19786 19556
rect 19996 19446 20024 24550
rect 20260 24132 20312 24138
rect 20260 24074 20312 24080
rect 20076 23520 20128 23526
rect 20076 23462 20128 23468
rect 20088 22642 20116 23462
rect 20272 22778 20300 24074
rect 20456 23118 20484 26250
rect 20812 23724 20864 23730
rect 20812 23666 20864 23672
rect 20720 23656 20772 23662
rect 20720 23598 20772 23604
rect 20536 23588 20588 23594
rect 20536 23530 20588 23536
rect 20548 23186 20576 23530
rect 20536 23180 20588 23186
rect 20536 23122 20588 23128
rect 20444 23112 20496 23118
rect 20444 23054 20496 23060
rect 20260 22772 20312 22778
rect 20260 22714 20312 22720
rect 20076 22636 20128 22642
rect 20076 22578 20128 22584
rect 20168 22024 20220 22030
rect 20168 21966 20220 21972
rect 20180 21554 20208 21966
rect 20456 21554 20484 23054
rect 20732 22574 20760 23598
rect 20824 23186 20852 23666
rect 21100 23322 21128 32370
rect 21192 31822 21220 32370
rect 21272 32360 21324 32366
rect 21272 32302 21324 32308
rect 21180 31816 21232 31822
rect 21180 31758 21232 31764
rect 21284 23322 21312 32302
rect 21376 30938 21404 38694
rect 22112 37466 22140 38830
rect 22284 38752 22336 38758
rect 22284 38694 22336 38700
rect 22296 37874 22324 38694
rect 22284 37868 22336 37874
rect 22284 37810 22336 37816
rect 22388 37738 22416 38898
rect 22836 38276 22888 38282
rect 22836 38218 22888 38224
rect 22560 38208 22612 38214
rect 22560 38150 22612 38156
rect 22572 37874 22600 38150
rect 22848 38010 22876 38218
rect 22836 38004 22888 38010
rect 22836 37946 22888 37952
rect 22560 37868 22612 37874
rect 22560 37810 22612 37816
rect 22376 37732 22428 37738
rect 22376 37674 22428 37680
rect 22100 37460 22152 37466
rect 22100 37402 22152 37408
rect 22388 37194 22416 37674
rect 22744 37664 22796 37670
rect 22744 37606 22796 37612
rect 22560 37256 22612 37262
rect 22560 37198 22612 37204
rect 22376 37188 22428 37194
rect 22376 37130 22428 37136
rect 21456 37120 21508 37126
rect 21456 37062 21508 37068
rect 21364 30932 21416 30938
rect 21364 30874 21416 30880
rect 21376 30190 21404 30874
rect 21364 30184 21416 30190
rect 21364 30126 21416 30132
rect 21468 29782 21496 37062
rect 22388 36242 22416 37130
rect 22468 36576 22520 36582
rect 22468 36518 22520 36524
rect 22480 36310 22508 36518
rect 22468 36304 22520 36310
rect 22468 36246 22520 36252
rect 22376 36236 22428 36242
rect 22376 36178 22428 36184
rect 22192 36168 22244 36174
rect 22192 36110 22244 36116
rect 21548 35760 21600 35766
rect 21548 35702 21600 35708
rect 21560 35494 21588 35702
rect 21548 35488 21600 35494
rect 21548 35430 21600 35436
rect 22204 35290 22232 36110
rect 22388 36038 22416 36178
rect 22376 36032 22428 36038
rect 22376 35974 22428 35980
rect 22284 35624 22336 35630
rect 22284 35566 22336 35572
rect 22192 35284 22244 35290
rect 22192 35226 22244 35232
rect 22296 35170 22324 35566
rect 22204 35142 22324 35170
rect 22100 34944 22152 34950
rect 22100 34886 22152 34892
rect 21824 33992 21876 33998
rect 21822 33960 21824 33969
rect 21876 33960 21878 33969
rect 21822 33895 21878 33904
rect 21732 32904 21784 32910
rect 21732 32846 21784 32852
rect 21548 32428 21600 32434
rect 21548 32370 21600 32376
rect 21560 31226 21588 32370
rect 21744 32230 21772 32846
rect 21732 32224 21784 32230
rect 21732 32166 21784 32172
rect 21744 31754 21772 32166
rect 22112 31822 22140 34886
rect 22204 34610 22232 35142
rect 22192 34604 22244 34610
rect 22192 34546 22244 34552
rect 22204 34066 22232 34546
rect 22192 34060 22244 34066
rect 22192 34002 22244 34008
rect 22388 33046 22416 35974
rect 22480 35698 22508 36246
rect 22468 35692 22520 35698
rect 22468 35634 22520 35640
rect 22480 33998 22508 35634
rect 22572 35154 22600 37198
rect 22652 36780 22704 36786
rect 22652 36722 22704 36728
rect 22664 35562 22692 36722
rect 22756 36174 22784 37606
rect 23308 36718 23336 45426
rect 25792 45422 25820 45902
rect 25976 45422 26004 46271
rect 26160 46034 26188 48991
rect 26240 46980 26292 46986
rect 26240 46922 26292 46928
rect 26252 46714 26280 46922
rect 27080 46918 27108 49200
rect 27068 46912 27120 46918
rect 27068 46854 27120 46860
rect 26240 46708 26292 46714
rect 26240 46650 26292 46656
rect 26976 46572 27028 46578
rect 26976 46514 27028 46520
rect 26424 46368 26476 46374
rect 26424 46310 26476 46316
rect 26148 46028 26200 46034
rect 26148 45970 26200 45976
rect 26240 45824 26292 45830
rect 26240 45766 26292 45772
rect 26252 45558 26280 45766
rect 26240 45552 26292 45558
rect 26240 45494 26292 45500
rect 26436 45490 26464 46310
rect 26988 46102 27016 46514
rect 27896 46368 27948 46374
rect 27896 46310 27948 46316
rect 26976 46096 27028 46102
rect 26976 46038 27028 46044
rect 26884 45824 26936 45830
rect 26884 45766 26936 45772
rect 26424 45484 26476 45490
rect 26424 45426 26476 45432
rect 25780 45416 25832 45422
rect 25780 45358 25832 45364
rect 25964 45416 26016 45422
rect 25964 45358 26016 45364
rect 24110 45180 24418 45200
rect 24110 45178 24116 45180
rect 24172 45178 24196 45180
rect 24252 45178 24276 45180
rect 24332 45178 24356 45180
rect 24412 45178 24418 45180
rect 24172 45126 24174 45178
rect 24354 45126 24356 45178
rect 24110 45124 24116 45126
rect 24172 45124 24196 45126
rect 24252 45124 24276 45126
rect 24332 45124 24356 45126
rect 24412 45124 24418 45126
rect 24110 45104 24418 45124
rect 26332 44192 26384 44198
rect 26332 44134 26384 44140
rect 24110 44092 24418 44112
rect 24110 44090 24116 44092
rect 24172 44090 24196 44092
rect 24252 44090 24276 44092
rect 24332 44090 24356 44092
rect 24412 44090 24418 44092
rect 24172 44038 24174 44090
rect 24354 44038 24356 44090
rect 24110 44036 24116 44038
rect 24172 44036 24196 44038
rect 24252 44036 24276 44038
rect 24332 44036 24356 44038
rect 24412 44036 24418 44038
rect 24110 44016 24418 44036
rect 24110 43004 24418 43024
rect 24110 43002 24116 43004
rect 24172 43002 24196 43004
rect 24252 43002 24276 43004
rect 24332 43002 24356 43004
rect 24412 43002 24418 43004
rect 24172 42950 24174 43002
rect 24354 42950 24356 43002
rect 24110 42948 24116 42950
rect 24172 42948 24196 42950
rect 24252 42948 24276 42950
rect 24332 42948 24356 42950
rect 24412 42948 24418 42950
rect 24110 42928 24418 42948
rect 26344 42770 26372 44134
rect 26516 43104 26568 43110
rect 26516 43046 26568 43052
rect 26528 42770 26556 43046
rect 26332 42764 26384 42770
rect 26332 42706 26384 42712
rect 26516 42764 26568 42770
rect 26516 42706 26568 42712
rect 26054 42256 26110 42265
rect 26054 42191 26110 42200
rect 24110 41916 24418 41936
rect 24110 41914 24116 41916
rect 24172 41914 24196 41916
rect 24252 41914 24276 41916
rect 24332 41914 24356 41916
rect 24412 41914 24418 41916
rect 24172 41862 24174 41914
rect 24354 41862 24356 41914
rect 24110 41860 24116 41862
rect 24172 41860 24196 41862
rect 24252 41860 24276 41862
rect 24332 41860 24356 41862
rect 24412 41860 24418 41862
rect 24110 41840 24418 41860
rect 25962 41576 26018 41585
rect 25962 41511 26018 41520
rect 25976 41070 26004 41511
rect 25964 41064 26016 41070
rect 25964 41006 26016 41012
rect 24110 40828 24418 40848
rect 24110 40826 24116 40828
rect 24172 40826 24196 40828
rect 24252 40826 24276 40828
rect 24332 40826 24356 40828
rect 24412 40826 24418 40828
rect 24172 40774 24174 40826
rect 24354 40774 24356 40826
rect 24110 40772 24116 40774
rect 24172 40772 24196 40774
rect 24252 40772 24276 40774
rect 24332 40772 24356 40774
rect 24412 40772 24418 40774
rect 24110 40752 24418 40772
rect 24110 39740 24418 39760
rect 24110 39738 24116 39740
rect 24172 39738 24196 39740
rect 24252 39738 24276 39740
rect 24332 39738 24356 39740
rect 24412 39738 24418 39740
rect 24172 39686 24174 39738
rect 24354 39686 24356 39738
rect 24110 39684 24116 39686
rect 24172 39684 24196 39686
rect 24252 39684 24276 39686
rect 24332 39684 24356 39686
rect 24412 39684 24418 39686
rect 24110 39664 24418 39684
rect 24110 38652 24418 38672
rect 24110 38650 24116 38652
rect 24172 38650 24196 38652
rect 24252 38650 24276 38652
rect 24332 38650 24356 38652
rect 24412 38650 24418 38652
rect 24172 38598 24174 38650
rect 24354 38598 24356 38650
rect 24110 38596 24116 38598
rect 24172 38596 24196 38598
rect 24252 38596 24276 38598
rect 24332 38596 24356 38598
rect 24412 38596 24418 38598
rect 24110 38576 24418 38596
rect 23756 38344 23808 38350
rect 23756 38286 23808 38292
rect 23296 36712 23348 36718
rect 23296 36654 23348 36660
rect 22744 36168 22796 36174
rect 22744 36110 22796 36116
rect 22652 35556 22704 35562
rect 22652 35498 22704 35504
rect 22756 35306 22784 36110
rect 23768 35494 23796 38286
rect 24110 37564 24418 37584
rect 24110 37562 24116 37564
rect 24172 37562 24196 37564
rect 24252 37562 24276 37564
rect 24332 37562 24356 37564
rect 24412 37562 24418 37564
rect 24172 37510 24174 37562
rect 24354 37510 24356 37562
rect 24110 37508 24116 37510
rect 24172 37508 24196 37510
rect 24252 37508 24276 37510
rect 24332 37508 24356 37510
rect 24412 37508 24418 37510
rect 24110 37488 24418 37508
rect 24110 36476 24418 36496
rect 24110 36474 24116 36476
rect 24172 36474 24196 36476
rect 24252 36474 24276 36476
rect 24332 36474 24356 36476
rect 24412 36474 24418 36476
rect 24172 36422 24174 36474
rect 24354 36422 24356 36474
rect 24110 36420 24116 36422
rect 24172 36420 24196 36422
rect 24252 36420 24276 36422
rect 24332 36420 24356 36422
rect 24412 36420 24418 36422
rect 24110 36400 24418 36420
rect 25228 36168 25280 36174
rect 25228 36110 25280 36116
rect 24400 36032 24452 36038
rect 24400 35974 24452 35980
rect 24412 35766 24440 35974
rect 25240 35834 25268 36110
rect 25596 36100 25648 36106
rect 25596 36042 25648 36048
rect 25228 35828 25280 35834
rect 25228 35770 25280 35776
rect 24400 35760 24452 35766
rect 24400 35702 24452 35708
rect 25608 35698 25636 36042
rect 25596 35692 25648 35698
rect 25596 35634 25648 35640
rect 23112 35488 23164 35494
rect 23112 35430 23164 35436
rect 23296 35488 23348 35494
rect 23296 35430 23348 35436
rect 23480 35488 23532 35494
rect 23480 35430 23532 35436
rect 23756 35488 23808 35494
rect 23756 35430 23808 35436
rect 24676 35488 24728 35494
rect 24676 35430 24728 35436
rect 22756 35278 22876 35306
rect 22560 35148 22612 35154
rect 22560 35090 22612 35096
rect 22468 33992 22520 33998
rect 22468 33934 22520 33940
rect 22376 33040 22428 33046
rect 22376 32982 22428 32988
rect 22572 32994 22600 35090
rect 22652 34060 22704 34066
rect 22652 34002 22704 34008
rect 22664 33590 22692 34002
rect 22652 33584 22704 33590
rect 22652 33526 22704 33532
rect 22744 33312 22796 33318
rect 22744 33254 22796 33260
rect 22572 32966 22692 32994
rect 22376 32904 22428 32910
rect 22376 32846 22428 32852
rect 22560 32904 22612 32910
rect 22560 32846 22612 32852
rect 22388 32337 22416 32846
rect 22468 32360 22520 32366
rect 22374 32328 22430 32337
rect 22468 32302 22520 32308
rect 22374 32263 22430 32272
rect 22284 32224 22336 32230
rect 22284 32166 22336 32172
rect 22100 31816 22152 31822
rect 22100 31758 22152 31764
rect 21744 31726 21864 31754
rect 21560 31198 21772 31226
rect 21640 30660 21692 30666
rect 21640 30602 21692 30608
rect 21456 29776 21508 29782
rect 21456 29718 21508 29724
rect 21456 29640 21508 29646
rect 21456 29582 21508 29588
rect 21468 28558 21496 29582
rect 21456 28552 21508 28558
rect 21456 28494 21508 28500
rect 21364 27600 21416 27606
rect 21364 27542 21416 27548
rect 21376 27402 21404 27542
rect 21364 27396 21416 27402
rect 21364 27338 21416 27344
rect 21468 27062 21496 28494
rect 21652 27606 21680 30602
rect 21744 30122 21772 31198
rect 21836 30258 21864 31726
rect 22112 31346 22140 31758
rect 22296 31754 22324 32166
rect 22480 31822 22508 32302
rect 22572 32026 22600 32846
rect 22560 32020 22612 32026
rect 22560 31962 22612 31968
rect 22664 31890 22692 32966
rect 22756 32910 22784 33254
rect 22744 32904 22796 32910
rect 22744 32846 22796 32852
rect 22756 32366 22784 32846
rect 22744 32360 22796 32366
rect 22744 32302 22796 32308
rect 22652 31884 22704 31890
rect 22652 31826 22704 31832
rect 22468 31816 22520 31822
rect 22468 31758 22520 31764
rect 22192 31748 22324 31754
rect 22244 31726 22324 31748
rect 22848 31754 22876 35278
rect 23124 35086 23152 35430
rect 23112 35080 23164 35086
rect 23112 35022 23164 35028
rect 23308 34406 23336 35430
rect 23296 34400 23348 34406
rect 23296 34342 23348 34348
rect 23308 34134 23336 34342
rect 23296 34128 23348 34134
rect 23296 34070 23348 34076
rect 23388 33992 23440 33998
rect 23388 33934 23440 33940
rect 23400 32842 23428 33934
rect 23492 33318 23520 35430
rect 24110 35388 24418 35408
rect 24110 35386 24116 35388
rect 24172 35386 24196 35388
rect 24252 35386 24276 35388
rect 24332 35386 24356 35388
rect 24412 35386 24418 35388
rect 24172 35334 24174 35386
rect 24354 35334 24356 35386
rect 24110 35332 24116 35334
rect 24172 35332 24196 35334
rect 24252 35332 24276 35334
rect 24332 35332 24356 35334
rect 24412 35332 24418 35334
rect 24110 35312 24418 35332
rect 23572 35216 23624 35222
rect 23572 35158 23624 35164
rect 23584 34202 23612 35158
rect 24688 35154 24716 35430
rect 23664 35148 23716 35154
rect 23664 35090 23716 35096
rect 24676 35148 24728 35154
rect 24676 35090 24728 35096
rect 23572 34196 23624 34202
rect 23572 34138 23624 34144
rect 23572 33584 23624 33590
rect 23572 33526 23624 33532
rect 23480 33312 23532 33318
rect 23480 33254 23532 33260
rect 23388 32836 23440 32842
rect 23388 32778 23440 32784
rect 23112 31884 23164 31890
rect 23112 31826 23164 31832
rect 22848 31726 23060 31754
rect 22192 31690 22244 31696
rect 22100 31340 22152 31346
rect 22100 31282 22152 31288
rect 22468 31340 22520 31346
rect 22468 31282 22520 31288
rect 21916 31136 21968 31142
rect 21916 31078 21968 31084
rect 21928 30802 21956 31078
rect 22112 30870 22140 31282
rect 22100 30864 22152 30870
rect 22100 30806 22152 30812
rect 21916 30796 21968 30802
rect 21916 30738 21968 30744
rect 21824 30252 21876 30258
rect 21824 30194 21876 30200
rect 21732 30116 21784 30122
rect 21732 30058 21784 30064
rect 21744 29646 21772 30058
rect 21836 29866 21864 30194
rect 21928 30190 21956 30738
rect 22480 30394 22508 31282
rect 22468 30388 22520 30394
rect 22468 30330 22520 30336
rect 22008 30252 22060 30258
rect 22008 30194 22060 30200
rect 21916 30184 21968 30190
rect 21916 30126 21968 30132
rect 21836 29838 21956 29866
rect 22020 29850 22048 30194
rect 21824 29708 21876 29714
rect 21824 29650 21876 29656
rect 21732 29640 21784 29646
rect 21732 29582 21784 29588
rect 21640 27600 21692 27606
rect 21640 27542 21692 27548
rect 21640 27396 21692 27402
rect 21640 27338 21692 27344
rect 21548 27328 21600 27334
rect 21548 27270 21600 27276
rect 21456 27056 21508 27062
rect 21456 26998 21508 27004
rect 21560 26586 21588 27270
rect 21548 26580 21600 26586
rect 21548 26522 21600 26528
rect 21560 26450 21588 26522
rect 21548 26444 21600 26450
rect 21548 26386 21600 26392
rect 21364 26376 21416 26382
rect 21416 26324 21588 26330
rect 21364 26318 21588 26324
rect 21376 26302 21588 26318
rect 21456 24064 21508 24070
rect 21456 24006 21508 24012
rect 21364 23860 21416 23866
rect 21364 23802 21416 23808
rect 21088 23316 21140 23322
rect 21088 23258 21140 23264
rect 21272 23316 21324 23322
rect 21272 23258 21324 23264
rect 20812 23180 20864 23186
rect 20812 23122 20864 23128
rect 20720 22568 20772 22574
rect 20720 22510 20772 22516
rect 20168 21548 20220 21554
rect 20168 21490 20220 21496
rect 20444 21548 20496 21554
rect 20444 21490 20496 21496
rect 20180 20806 20208 21490
rect 20456 20942 20484 21490
rect 20444 20936 20496 20942
rect 20444 20878 20496 20884
rect 20168 20800 20220 20806
rect 20168 20742 20220 20748
rect 19984 19440 20036 19446
rect 19984 19382 20036 19388
rect 19340 19236 19392 19242
rect 19340 19178 19392 19184
rect 19352 18086 19380 19178
rect 19478 18524 19786 18544
rect 19478 18522 19484 18524
rect 19540 18522 19564 18524
rect 19620 18522 19644 18524
rect 19700 18522 19724 18524
rect 19780 18522 19786 18524
rect 19540 18470 19542 18522
rect 19722 18470 19724 18522
rect 19478 18468 19484 18470
rect 19540 18468 19564 18470
rect 19620 18468 19644 18470
rect 19700 18468 19724 18470
rect 19780 18468 19786 18470
rect 19478 18448 19786 18468
rect 19340 18080 19392 18086
rect 19340 18022 19392 18028
rect 18788 17876 18840 17882
rect 18788 17818 18840 17824
rect 19352 16658 19380 18022
rect 19892 17604 19944 17610
rect 19892 17546 19944 17552
rect 19478 17436 19786 17456
rect 19478 17434 19484 17436
rect 19540 17434 19564 17436
rect 19620 17434 19644 17436
rect 19700 17434 19724 17436
rect 19780 17434 19786 17436
rect 19540 17382 19542 17434
rect 19722 17382 19724 17434
rect 19478 17380 19484 17382
rect 19540 17380 19564 17382
rect 19620 17380 19644 17382
rect 19700 17380 19724 17382
rect 19780 17380 19786 17382
rect 19478 17360 19786 17380
rect 19340 16652 19392 16658
rect 19340 16594 19392 16600
rect 19340 16448 19392 16454
rect 19340 16390 19392 16396
rect 19248 16176 19300 16182
rect 19248 16118 19300 16124
rect 18696 16040 18748 16046
rect 18696 15982 18748 15988
rect 18708 15706 18736 15982
rect 19260 15706 19288 16118
rect 18696 15700 18748 15706
rect 18696 15642 18748 15648
rect 19248 15700 19300 15706
rect 19248 15642 19300 15648
rect 19156 15632 19208 15638
rect 19156 15574 19208 15580
rect 19352 15586 19380 16390
rect 19478 16348 19786 16368
rect 19478 16346 19484 16348
rect 19540 16346 19564 16348
rect 19620 16346 19644 16348
rect 19700 16346 19724 16348
rect 19780 16346 19786 16348
rect 19540 16294 19542 16346
rect 19722 16294 19724 16346
rect 19478 16292 19484 16294
rect 19540 16292 19564 16294
rect 19620 16292 19644 16294
rect 19700 16292 19724 16294
rect 19780 16292 19786 16294
rect 19478 16272 19786 16292
rect 19904 16250 19932 17546
rect 20180 17202 20208 20742
rect 20732 20262 20760 22510
rect 20824 21894 20852 23122
rect 21088 22976 21140 22982
rect 21376 22930 21404 23802
rect 21468 23730 21496 24006
rect 21456 23724 21508 23730
rect 21456 23666 21508 23672
rect 21560 23526 21588 26302
rect 21652 23526 21680 27338
rect 21744 23798 21772 29582
rect 21836 28762 21864 29650
rect 21824 28756 21876 28762
rect 21824 28698 21876 28704
rect 21836 28150 21864 28698
rect 21824 28144 21876 28150
rect 21824 28086 21876 28092
rect 21836 28014 21864 28086
rect 21824 28008 21876 28014
rect 21824 27950 21876 27956
rect 21928 26874 21956 29838
rect 22008 29844 22060 29850
rect 22008 29786 22060 29792
rect 23032 29714 23060 31726
rect 23020 29708 23072 29714
rect 23020 29650 23072 29656
rect 22560 29640 22612 29646
rect 22612 29600 22692 29628
rect 22560 29582 22612 29588
rect 22100 28552 22152 28558
rect 22100 28494 22152 28500
rect 22112 28218 22140 28494
rect 22664 28422 22692 29600
rect 22744 28552 22796 28558
rect 22744 28494 22796 28500
rect 22560 28416 22612 28422
rect 22560 28358 22612 28364
rect 22652 28416 22704 28422
rect 22652 28358 22704 28364
rect 22100 28212 22152 28218
rect 22100 28154 22152 28160
rect 22572 28150 22600 28358
rect 22560 28144 22612 28150
rect 22560 28086 22612 28092
rect 22376 28076 22428 28082
rect 22376 28018 22428 28024
rect 22388 27470 22416 28018
rect 22664 27996 22692 28358
rect 22572 27968 22692 27996
rect 22572 27878 22600 27968
rect 22560 27872 22612 27878
rect 22560 27814 22612 27820
rect 22376 27464 22428 27470
rect 22376 27406 22428 27412
rect 22192 26988 22244 26994
rect 22192 26930 22244 26936
rect 21836 26846 21956 26874
rect 21836 24834 21864 26846
rect 21916 26784 21968 26790
rect 21916 26726 21968 26732
rect 21928 26450 21956 26726
rect 21916 26444 21968 26450
rect 21916 26386 21968 26392
rect 22008 26240 22060 26246
rect 22060 26188 22140 26194
rect 22008 26182 22140 26188
rect 22020 26166 22140 26182
rect 21836 24806 22048 24834
rect 21824 24744 21876 24750
rect 21824 24686 21876 24692
rect 21836 24206 21864 24686
rect 21824 24200 21876 24206
rect 21824 24142 21876 24148
rect 21732 23792 21784 23798
rect 21732 23734 21784 23740
rect 21916 23792 21968 23798
rect 21916 23734 21968 23740
rect 21824 23588 21876 23594
rect 21824 23530 21876 23536
rect 21548 23520 21600 23526
rect 21548 23462 21600 23468
rect 21640 23520 21692 23526
rect 21640 23462 21692 23468
rect 21456 23180 21508 23186
rect 21456 23122 21508 23128
rect 21468 23050 21496 23122
rect 21456 23044 21508 23050
rect 21456 22986 21508 22992
rect 21088 22918 21140 22924
rect 20904 22024 20956 22030
rect 20904 21966 20956 21972
rect 20812 21888 20864 21894
rect 20812 21830 20864 21836
rect 20824 21622 20852 21830
rect 20812 21616 20864 21622
rect 20812 21558 20864 21564
rect 20812 21344 20864 21350
rect 20812 21286 20864 21292
rect 20824 20534 20852 21286
rect 20812 20528 20864 20534
rect 20812 20470 20864 20476
rect 20720 20256 20772 20262
rect 20720 20198 20772 20204
rect 20916 19854 20944 21966
rect 21100 21026 21128 22918
rect 21284 22902 21404 22930
rect 21100 20998 21220 21026
rect 21088 20936 21140 20942
rect 21088 20878 21140 20884
rect 21100 20602 21128 20878
rect 21088 20596 21140 20602
rect 21088 20538 21140 20544
rect 20996 20528 21048 20534
rect 20996 20470 21048 20476
rect 21008 20262 21036 20470
rect 20996 20256 21048 20262
rect 20996 20198 21048 20204
rect 20904 19848 20956 19854
rect 20904 19790 20956 19796
rect 21008 19174 21036 20198
rect 21100 19854 21128 20538
rect 21088 19848 21140 19854
rect 21088 19790 21140 19796
rect 20996 19168 21048 19174
rect 20996 19110 21048 19116
rect 20812 18420 20864 18426
rect 20812 18362 20864 18368
rect 20628 18080 20680 18086
rect 20628 18022 20680 18028
rect 20640 17610 20668 18022
rect 20628 17604 20680 17610
rect 20628 17546 20680 17552
rect 20168 17196 20220 17202
rect 20168 17138 20220 17144
rect 20628 17196 20680 17202
rect 20628 17138 20680 17144
rect 20260 16992 20312 16998
rect 20260 16934 20312 16940
rect 19984 16652 20036 16658
rect 19984 16594 20036 16600
rect 19892 16244 19944 16250
rect 19892 16186 19944 16192
rect 19892 16040 19944 16046
rect 19892 15982 19944 15988
rect 19168 15366 19196 15574
rect 19352 15558 19564 15586
rect 19536 15502 19564 15558
rect 19432 15496 19484 15502
rect 19352 15444 19432 15450
rect 19352 15438 19484 15444
rect 19524 15496 19576 15502
rect 19524 15438 19576 15444
rect 19352 15422 19472 15438
rect 18696 15360 18748 15366
rect 18696 15302 18748 15308
rect 19156 15360 19208 15366
rect 19156 15302 19208 15308
rect 18708 14074 18736 15302
rect 19352 14822 19380 15422
rect 19478 15260 19786 15280
rect 19478 15258 19484 15260
rect 19540 15258 19564 15260
rect 19620 15258 19644 15260
rect 19700 15258 19724 15260
rect 19780 15258 19786 15260
rect 19540 15206 19542 15258
rect 19722 15206 19724 15258
rect 19478 15204 19484 15206
rect 19540 15204 19564 15206
rect 19620 15204 19644 15206
rect 19700 15204 19724 15206
rect 19780 15204 19786 15206
rect 19478 15184 19786 15204
rect 19340 14816 19392 14822
rect 19340 14758 19392 14764
rect 19340 14476 19392 14482
rect 19340 14418 19392 14424
rect 18696 14068 18748 14074
rect 18696 14010 18748 14016
rect 18696 12232 18748 12238
rect 19352 12186 19380 14418
rect 19478 14172 19786 14192
rect 19478 14170 19484 14172
rect 19540 14170 19564 14172
rect 19620 14170 19644 14172
rect 19700 14170 19724 14172
rect 19780 14170 19786 14172
rect 19540 14118 19542 14170
rect 19722 14118 19724 14170
rect 19478 14116 19484 14118
rect 19540 14116 19564 14118
rect 19620 14116 19644 14118
rect 19700 14116 19724 14118
rect 19780 14116 19786 14118
rect 19478 14096 19786 14116
rect 19800 13932 19852 13938
rect 19800 13874 19852 13880
rect 19812 13530 19840 13874
rect 19800 13524 19852 13530
rect 19800 13466 19852 13472
rect 19478 13084 19786 13104
rect 19478 13082 19484 13084
rect 19540 13082 19564 13084
rect 19620 13082 19644 13084
rect 19700 13082 19724 13084
rect 19780 13082 19786 13084
rect 19540 13030 19542 13082
rect 19722 13030 19724 13082
rect 19478 13028 19484 13030
rect 19540 13028 19564 13030
rect 19620 13028 19644 13030
rect 19700 13028 19724 13030
rect 19780 13028 19786 13030
rect 19478 13008 19786 13028
rect 18696 12174 18748 12180
rect 18708 11762 18736 12174
rect 19260 12158 19380 12186
rect 18696 11756 18748 11762
rect 18696 11698 18748 11704
rect 18708 11354 18736 11698
rect 18696 11348 18748 11354
rect 18696 11290 18748 11296
rect 19260 11082 19288 12158
rect 19340 12096 19392 12102
rect 19340 12038 19392 12044
rect 19352 11830 19380 12038
rect 19478 11996 19786 12016
rect 19478 11994 19484 11996
rect 19540 11994 19564 11996
rect 19620 11994 19644 11996
rect 19700 11994 19724 11996
rect 19780 11994 19786 11996
rect 19540 11942 19542 11994
rect 19722 11942 19724 11994
rect 19478 11940 19484 11942
rect 19540 11940 19564 11942
rect 19620 11940 19644 11942
rect 19700 11940 19724 11942
rect 19780 11940 19786 11942
rect 19478 11920 19786 11940
rect 19904 11898 19932 15982
rect 19996 15094 20024 16594
rect 20272 16590 20300 16934
rect 20260 16584 20312 16590
rect 20260 16526 20312 16532
rect 20640 15638 20668 17138
rect 20824 16658 20852 18362
rect 21008 17678 21036 19110
rect 21192 18290 21220 20998
rect 21284 18766 21312 22902
rect 21468 22710 21496 22986
rect 21456 22704 21508 22710
rect 21456 22646 21508 22652
rect 21560 22094 21588 23462
rect 21376 22066 21588 22094
rect 21376 21962 21404 22066
rect 21652 22030 21680 23462
rect 21836 23186 21864 23530
rect 21824 23180 21876 23186
rect 21824 23122 21876 23128
rect 21928 23050 21956 23734
rect 22020 23662 22048 24806
rect 22112 24750 22140 26166
rect 22204 25498 22232 26930
rect 22572 25906 22600 27814
rect 22652 27464 22704 27470
rect 22652 27406 22704 27412
rect 22560 25900 22612 25906
rect 22560 25842 22612 25848
rect 22192 25492 22244 25498
rect 22192 25434 22244 25440
rect 22100 24744 22152 24750
rect 22100 24686 22152 24692
rect 22376 24132 22428 24138
rect 22376 24074 22428 24080
rect 22388 23866 22416 24074
rect 22376 23860 22428 23866
rect 22376 23802 22428 23808
rect 22008 23656 22060 23662
rect 22008 23598 22060 23604
rect 22100 23520 22152 23526
rect 22006 23488 22062 23497
rect 22100 23462 22152 23468
rect 22006 23423 22062 23432
rect 21916 23044 21968 23050
rect 21916 22986 21968 22992
rect 21824 22976 21876 22982
rect 21824 22918 21876 22924
rect 21640 22024 21692 22030
rect 21640 21966 21692 21972
rect 21364 21956 21416 21962
rect 21364 21898 21416 21904
rect 21364 21684 21416 21690
rect 21364 21626 21416 21632
rect 21376 20058 21404 21626
rect 21732 21344 21784 21350
rect 21732 21286 21784 21292
rect 21744 20942 21772 21286
rect 21456 20936 21508 20942
rect 21456 20878 21508 20884
rect 21732 20936 21784 20942
rect 21732 20878 21784 20884
rect 21468 20534 21496 20878
rect 21456 20528 21508 20534
rect 21456 20470 21508 20476
rect 21364 20052 21416 20058
rect 21364 19994 21416 20000
rect 21836 18970 21864 22918
rect 21928 22710 21956 22986
rect 21916 22704 21968 22710
rect 21916 22646 21968 22652
rect 22020 22438 22048 23423
rect 22008 22432 22060 22438
rect 22008 22374 22060 22380
rect 22006 21584 22062 21593
rect 22006 21519 22008 21528
rect 22060 21519 22062 21528
rect 22008 21490 22060 21496
rect 21824 18964 21876 18970
rect 21824 18906 21876 18912
rect 22020 18766 22048 21490
rect 21272 18760 21324 18766
rect 21272 18702 21324 18708
rect 21916 18760 21968 18766
rect 21916 18702 21968 18708
rect 22008 18760 22060 18766
rect 22008 18702 22060 18708
rect 21180 18284 21232 18290
rect 21180 18226 21232 18232
rect 21088 18216 21140 18222
rect 21284 18170 21312 18702
rect 21928 18426 21956 18702
rect 21916 18420 21968 18426
rect 21916 18362 21968 18368
rect 22020 18290 22048 18702
rect 22112 18358 22140 23462
rect 22572 23050 22600 25842
rect 22664 25838 22692 27406
rect 22756 26858 22784 28494
rect 23032 28082 23060 29650
rect 23124 29646 23152 31826
rect 23492 31142 23520 33254
rect 23584 33114 23612 33526
rect 23572 33108 23624 33114
rect 23572 33050 23624 33056
rect 23676 33046 23704 35090
rect 24688 34678 24716 35090
rect 25608 35018 25636 35634
rect 25872 35624 25924 35630
rect 25872 35566 25924 35572
rect 25596 35012 25648 35018
rect 25596 34954 25648 34960
rect 24860 34944 24912 34950
rect 24860 34886 24912 34892
rect 24676 34672 24728 34678
rect 24676 34614 24728 34620
rect 24110 34300 24418 34320
rect 24110 34298 24116 34300
rect 24172 34298 24196 34300
rect 24252 34298 24276 34300
rect 24332 34298 24356 34300
rect 24412 34298 24418 34300
rect 24172 34246 24174 34298
rect 24354 34246 24356 34298
rect 24110 34244 24116 34246
rect 24172 34244 24196 34246
rect 24252 34244 24276 34246
rect 24332 34244 24356 34246
rect 24412 34244 24418 34246
rect 24110 34224 24418 34244
rect 23848 33924 23900 33930
rect 23848 33866 23900 33872
rect 24584 33924 24636 33930
rect 24584 33866 24636 33872
rect 23664 33040 23716 33046
rect 23664 32982 23716 32988
rect 23664 32768 23716 32774
rect 23664 32710 23716 32716
rect 23676 32434 23704 32710
rect 23664 32428 23716 32434
rect 23664 32370 23716 32376
rect 23676 32026 23704 32370
rect 23664 32020 23716 32026
rect 23664 31962 23716 31968
rect 23860 31822 23888 33866
rect 24596 33658 24624 33866
rect 24584 33652 24636 33658
rect 24584 33594 24636 33600
rect 24110 33212 24418 33232
rect 24110 33210 24116 33212
rect 24172 33210 24196 33212
rect 24252 33210 24276 33212
rect 24332 33210 24356 33212
rect 24412 33210 24418 33212
rect 24172 33158 24174 33210
rect 24354 33158 24356 33210
rect 24110 33156 24116 33158
rect 24172 33156 24196 33158
rect 24252 33156 24276 33158
rect 24332 33156 24356 33158
rect 24412 33156 24418 33158
rect 24110 33136 24418 33156
rect 24110 32124 24418 32144
rect 24110 32122 24116 32124
rect 24172 32122 24196 32124
rect 24252 32122 24276 32124
rect 24332 32122 24356 32124
rect 24412 32122 24418 32124
rect 24172 32070 24174 32122
rect 24354 32070 24356 32122
rect 24110 32068 24116 32070
rect 24172 32068 24196 32070
rect 24252 32068 24276 32070
rect 24332 32068 24356 32070
rect 24412 32068 24418 32070
rect 24110 32048 24418 32068
rect 23848 31816 23900 31822
rect 23848 31758 23900 31764
rect 23860 31482 23888 31758
rect 24872 31754 24900 34886
rect 25044 34400 25096 34406
rect 25044 34342 25096 34348
rect 25056 33998 25084 34342
rect 25044 33992 25096 33998
rect 25044 33934 25096 33940
rect 25136 33856 25188 33862
rect 25136 33798 25188 33804
rect 25148 33522 25176 33798
rect 25136 33516 25188 33522
rect 25136 33458 25188 33464
rect 24872 31726 24992 31754
rect 23848 31476 23900 31482
rect 23848 31418 23900 31424
rect 23480 31136 23532 31142
rect 23480 31078 23532 31084
rect 23492 30122 23520 31078
rect 24110 31036 24418 31056
rect 24110 31034 24116 31036
rect 24172 31034 24196 31036
rect 24252 31034 24276 31036
rect 24332 31034 24356 31036
rect 24412 31034 24418 31036
rect 24172 30982 24174 31034
rect 24354 30982 24356 31034
rect 24110 30980 24116 30982
rect 24172 30980 24196 30982
rect 24252 30980 24276 30982
rect 24332 30980 24356 30982
rect 24412 30980 24418 30982
rect 24110 30960 24418 30980
rect 24860 30728 24912 30734
rect 24860 30670 24912 30676
rect 23480 30116 23532 30122
rect 23480 30058 23532 30064
rect 24032 30116 24084 30122
rect 24032 30058 24084 30064
rect 23664 29708 23716 29714
rect 23664 29650 23716 29656
rect 23112 29640 23164 29646
rect 23112 29582 23164 29588
rect 23572 29640 23624 29646
rect 23572 29582 23624 29588
rect 23020 28076 23072 28082
rect 23020 28018 23072 28024
rect 22836 27056 22888 27062
rect 22836 26998 22888 27004
rect 22744 26852 22796 26858
rect 22744 26794 22796 26800
rect 22756 26382 22784 26794
rect 22744 26376 22796 26382
rect 22744 26318 22796 26324
rect 22756 26042 22784 26318
rect 22848 26314 22876 26998
rect 22928 26988 22980 26994
rect 22928 26930 22980 26936
rect 22836 26308 22888 26314
rect 22836 26250 22888 26256
rect 22744 26036 22796 26042
rect 22744 25978 22796 25984
rect 22652 25832 22704 25838
rect 22652 25774 22704 25780
rect 22756 25362 22784 25978
rect 22848 25378 22876 26250
rect 22940 25498 22968 26930
rect 23032 25906 23060 28018
rect 23124 27606 23152 29582
rect 23296 28552 23348 28558
rect 23348 28500 23428 28506
rect 23296 28494 23428 28500
rect 23308 28478 23428 28494
rect 23296 28416 23348 28422
rect 23296 28358 23348 28364
rect 23204 28076 23256 28082
rect 23204 28018 23256 28024
rect 23216 27674 23244 28018
rect 23204 27668 23256 27674
rect 23204 27610 23256 27616
rect 23112 27600 23164 27606
rect 23112 27542 23164 27548
rect 23020 25900 23072 25906
rect 23020 25842 23072 25848
rect 22928 25492 22980 25498
rect 22928 25434 22980 25440
rect 22848 25362 22968 25378
rect 22744 25356 22796 25362
rect 22848 25356 22980 25362
rect 22848 25350 22928 25356
rect 22744 25298 22796 25304
rect 22928 25298 22980 25304
rect 23032 24410 23060 25842
rect 23124 25362 23152 27542
rect 23308 27334 23336 28358
rect 23400 27470 23428 28478
rect 23584 28082 23612 29582
rect 23676 28762 23704 29650
rect 24044 29646 24072 30058
rect 24110 29948 24418 29968
rect 24110 29946 24116 29948
rect 24172 29946 24196 29948
rect 24252 29946 24276 29948
rect 24332 29946 24356 29948
rect 24412 29946 24418 29948
rect 24172 29894 24174 29946
rect 24354 29894 24356 29946
rect 24110 29892 24116 29894
rect 24172 29892 24196 29894
rect 24252 29892 24276 29894
rect 24332 29892 24356 29894
rect 24412 29892 24418 29894
rect 24110 29872 24418 29892
rect 24032 29640 24084 29646
rect 24032 29582 24084 29588
rect 23664 28756 23716 28762
rect 23664 28698 23716 28704
rect 23572 28076 23624 28082
rect 23572 28018 23624 28024
rect 23388 27464 23440 27470
rect 23388 27406 23440 27412
rect 23296 27328 23348 27334
rect 23296 27270 23348 27276
rect 23204 26580 23256 26586
rect 23204 26522 23256 26528
rect 23216 26382 23244 26522
rect 23308 26382 23336 27270
rect 23388 26784 23440 26790
rect 23388 26726 23440 26732
rect 23204 26376 23256 26382
rect 23204 26318 23256 26324
rect 23296 26376 23348 26382
rect 23296 26318 23348 26324
rect 23308 26246 23336 26318
rect 23296 26240 23348 26246
rect 23296 26182 23348 26188
rect 23204 25832 23256 25838
rect 23204 25774 23256 25780
rect 23112 25356 23164 25362
rect 23112 25298 23164 25304
rect 23020 24404 23072 24410
rect 23020 24346 23072 24352
rect 22560 23044 22612 23050
rect 22560 22986 22612 22992
rect 22744 22976 22796 22982
rect 22744 22918 22796 22924
rect 22192 22432 22244 22438
rect 22192 22374 22244 22380
rect 22204 21554 22232 22374
rect 22756 22030 22784 22918
rect 22928 22636 22980 22642
rect 22928 22578 22980 22584
rect 22940 22234 22968 22578
rect 22928 22228 22980 22234
rect 22928 22170 22980 22176
rect 22744 22024 22796 22030
rect 22744 21966 22796 21972
rect 22192 21548 22244 21554
rect 22192 21490 22244 21496
rect 22284 21480 22336 21486
rect 22284 21422 22336 21428
rect 22296 20058 22324 21422
rect 23216 21010 23244 25774
rect 23308 25362 23336 26182
rect 23400 25906 23428 26726
rect 23480 26376 23532 26382
rect 23480 26318 23532 26324
rect 23388 25900 23440 25906
rect 23388 25842 23440 25848
rect 23296 25356 23348 25362
rect 23296 25298 23348 25304
rect 23492 25226 23520 26318
rect 23584 25906 23612 28018
rect 24044 28014 24072 29582
rect 24110 28860 24418 28880
rect 24110 28858 24116 28860
rect 24172 28858 24196 28860
rect 24252 28858 24276 28860
rect 24332 28858 24356 28860
rect 24412 28858 24418 28860
rect 24172 28806 24174 28858
rect 24354 28806 24356 28858
rect 24110 28804 24116 28806
rect 24172 28804 24196 28806
rect 24252 28804 24276 28806
rect 24332 28804 24356 28806
rect 24412 28804 24418 28806
rect 24110 28784 24418 28804
rect 24032 28008 24084 28014
rect 24032 27950 24084 27956
rect 23848 27464 23900 27470
rect 23848 27406 23900 27412
rect 23860 26586 23888 27406
rect 23848 26580 23900 26586
rect 23848 26522 23900 26528
rect 23756 26512 23808 26518
rect 23756 26454 23808 26460
rect 23664 26240 23716 26246
rect 23664 26182 23716 26188
rect 23676 25974 23704 26182
rect 23768 25974 23796 26454
rect 23664 25968 23716 25974
rect 23664 25910 23716 25916
rect 23756 25968 23808 25974
rect 23756 25910 23808 25916
rect 23572 25900 23624 25906
rect 23572 25842 23624 25848
rect 23584 25498 23612 25842
rect 23860 25786 23888 26522
rect 24044 26382 24072 27950
rect 24110 27772 24418 27792
rect 24110 27770 24116 27772
rect 24172 27770 24196 27772
rect 24252 27770 24276 27772
rect 24332 27770 24356 27772
rect 24412 27770 24418 27772
rect 24172 27718 24174 27770
rect 24354 27718 24356 27770
rect 24110 27716 24116 27718
rect 24172 27716 24196 27718
rect 24252 27716 24276 27718
rect 24332 27716 24356 27718
rect 24412 27716 24418 27718
rect 24110 27696 24418 27716
rect 24110 26684 24418 26704
rect 24110 26682 24116 26684
rect 24172 26682 24196 26684
rect 24252 26682 24276 26684
rect 24332 26682 24356 26684
rect 24412 26682 24418 26684
rect 24172 26630 24174 26682
rect 24354 26630 24356 26682
rect 24110 26628 24116 26630
rect 24172 26628 24196 26630
rect 24252 26628 24276 26630
rect 24332 26628 24356 26630
rect 24412 26628 24418 26630
rect 24110 26608 24418 26628
rect 24032 26376 24084 26382
rect 24032 26318 24084 26324
rect 23768 25758 23888 25786
rect 23572 25492 23624 25498
rect 23572 25434 23624 25440
rect 23768 25294 23796 25758
rect 24044 25294 24072 26318
rect 24492 26308 24544 26314
rect 24492 26250 24544 26256
rect 24504 25770 24532 26250
rect 24492 25764 24544 25770
rect 24492 25706 24544 25712
rect 24676 25764 24728 25770
rect 24676 25706 24728 25712
rect 24110 25596 24418 25616
rect 24110 25594 24116 25596
rect 24172 25594 24196 25596
rect 24252 25594 24276 25596
rect 24332 25594 24356 25596
rect 24412 25594 24418 25596
rect 24172 25542 24174 25594
rect 24354 25542 24356 25594
rect 24110 25540 24116 25542
rect 24172 25540 24196 25542
rect 24252 25540 24276 25542
rect 24332 25540 24356 25542
rect 24412 25540 24418 25542
rect 24110 25520 24418 25540
rect 23756 25288 23808 25294
rect 23756 25230 23808 25236
rect 24032 25288 24084 25294
rect 24032 25230 24084 25236
rect 23480 25220 23532 25226
rect 23480 25162 23532 25168
rect 23940 25152 23992 25158
rect 23940 25094 23992 25100
rect 23664 23180 23716 23186
rect 23664 23122 23716 23128
rect 23388 23112 23440 23118
rect 23388 23054 23440 23060
rect 23400 22778 23428 23054
rect 23480 22976 23532 22982
rect 23480 22918 23532 22924
rect 23492 22778 23520 22918
rect 23388 22772 23440 22778
rect 23388 22714 23440 22720
rect 23480 22772 23532 22778
rect 23480 22714 23532 22720
rect 23676 22098 23704 23122
rect 23664 22092 23716 22098
rect 23664 22034 23716 22040
rect 23676 21690 23704 22034
rect 23664 21684 23716 21690
rect 23664 21626 23716 21632
rect 23204 21004 23256 21010
rect 23204 20946 23256 20952
rect 23572 20936 23624 20942
rect 23572 20878 23624 20884
rect 22468 20800 22520 20806
rect 22468 20742 22520 20748
rect 22836 20800 22888 20806
rect 22836 20742 22888 20748
rect 22480 20398 22508 20742
rect 22848 20602 22876 20742
rect 22836 20596 22888 20602
rect 22836 20538 22888 20544
rect 22468 20392 22520 20398
rect 22468 20334 22520 20340
rect 22284 20052 22336 20058
rect 22284 19994 22336 20000
rect 22192 19984 22244 19990
rect 22192 19926 22244 19932
rect 22204 19786 22232 19926
rect 22192 19780 22244 19786
rect 22192 19722 22244 19728
rect 22480 19718 22508 20334
rect 22848 19922 22876 20538
rect 23480 20460 23532 20466
rect 23480 20402 23532 20408
rect 23388 20256 23440 20262
rect 23388 20198 23440 20204
rect 22836 19916 22888 19922
rect 22836 19858 22888 19864
rect 23400 19854 23428 20198
rect 23492 19922 23520 20402
rect 23584 20058 23612 20878
rect 23756 20800 23808 20806
rect 23756 20742 23808 20748
rect 23768 20534 23796 20742
rect 23756 20528 23808 20534
rect 23756 20470 23808 20476
rect 23572 20052 23624 20058
rect 23572 19994 23624 20000
rect 23480 19916 23532 19922
rect 23480 19858 23532 19864
rect 22744 19848 22796 19854
rect 22744 19790 22796 19796
rect 23388 19848 23440 19854
rect 23388 19790 23440 19796
rect 22468 19712 22520 19718
rect 22468 19654 22520 19660
rect 22376 18624 22428 18630
rect 22376 18566 22428 18572
rect 22100 18352 22152 18358
rect 22100 18294 22152 18300
rect 22008 18284 22060 18290
rect 22008 18226 22060 18232
rect 21088 18158 21140 18164
rect 20996 17672 21048 17678
rect 20996 17614 21048 17620
rect 20812 16652 20864 16658
rect 20812 16594 20864 16600
rect 20720 16108 20772 16114
rect 20720 16050 20772 16056
rect 20732 15706 20760 16050
rect 20720 15700 20772 15706
rect 20720 15642 20772 15648
rect 20628 15632 20680 15638
rect 20628 15574 20680 15580
rect 19984 15088 20036 15094
rect 19984 15030 20036 15036
rect 20536 15020 20588 15026
rect 20536 14962 20588 14968
rect 20260 14952 20312 14958
rect 20260 14894 20312 14900
rect 19984 14816 20036 14822
rect 19984 14758 20036 14764
rect 19996 14414 20024 14758
rect 19984 14408 20036 14414
rect 19984 14350 20036 14356
rect 20076 14272 20128 14278
rect 20076 14214 20128 14220
rect 20088 13326 20116 14214
rect 20076 13320 20128 13326
rect 20076 13262 20128 13268
rect 19892 11892 19944 11898
rect 19892 11834 19944 11840
rect 19340 11824 19392 11830
rect 19340 11766 19392 11772
rect 19984 11756 20036 11762
rect 19984 11698 20036 11704
rect 19340 11620 19392 11626
rect 19340 11562 19392 11568
rect 19248 11076 19300 11082
rect 19248 11018 19300 11024
rect 19352 11014 19380 11562
rect 19340 11008 19392 11014
rect 19340 10950 19392 10956
rect 19352 10810 19380 10950
rect 19478 10908 19786 10928
rect 19478 10906 19484 10908
rect 19540 10906 19564 10908
rect 19620 10906 19644 10908
rect 19700 10906 19724 10908
rect 19780 10906 19786 10908
rect 19540 10854 19542 10906
rect 19722 10854 19724 10906
rect 19478 10852 19484 10854
rect 19540 10852 19564 10854
rect 19620 10852 19644 10854
rect 19700 10852 19724 10854
rect 19780 10852 19786 10854
rect 19478 10832 19786 10852
rect 19996 10810 20024 11698
rect 19340 10804 19392 10810
rect 19340 10746 19392 10752
rect 19984 10804 20036 10810
rect 19984 10746 20036 10752
rect 20272 10606 20300 14894
rect 20548 14890 20576 14962
rect 20536 14884 20588 14890
rect 20536 14826 20588 14832
rect 20548 14074 20576 14826
rect 20824 14482 20852 16594
rect 20812 14476 20864 14482
rect 20812 14418 20864 14424
rect 20536 14068 20588 14074
rect 20536 14010 20588 14016
rect 20824 12850 20852 14418
rect 21008 14414 21036 17614
rect 21100 17338 21128 18158
rect 21192 18142 21312 18170
rect 22100 18216 22152 18222
rect 22100 18158 22152 18164
rect 21088 17332 21140 17338
rect 21088 17274 21140 17280
rect 21192 16726 21220 18142
rect 21272 18080 21324 18086
rect 21272 18022 21324 18028
rect 21180 16720 21232 16726
rect 21180 16662 21232 16668
rect 20996 14408 21048 14414
rect 20996 14350 21048 14356
rect 21008 14006 21036 14350
rect 20996 14000 21048 14006
rect 20996 13942 21048 13948
rect 21192 13462 21220 16662
rect 21284 14346 21312 18022
rect 21364 17536 21416 17542
rect 21364 17478 21416 17484
rect 21376 17134 21404 17478
rect 22112 17202 22140 18158
rect 22388 17610 22416 18566
rect 22756 18290 22784 19790
rect 22836 19780 22888 19786
rect 22836 19722 22888 19728
rect 22848 18358 22876 19722
rect 23664 19712 23716 19718
rect 23664 19654 23716 19660
rect 22836 18352 22888 18358
rect 22836 18294 22888 18300
rect 22744 18284 22796 18290
rect 22744 18226 22796 18232
rect 22376 17604 22428 17610
rect 22376 17546 22428 17552
rect 22192 17332 22244 17338
rect 22192 17274 22244 17280
rect 22100 17196 22152 17202
rect 22100 17138 22152 17144
rect 22204 17134 22232 17274
rect 22756 17270 22784 18226
rect 22848 17338 22876 18294
rect 23204 18216 23256 18222
rect 23204 18158 23256 18164
rect 23480 18216 23532 18222
rect 23480 18158 23532 18164
rect 23216 17882 23244 18158
rect 23204 17876 23256 17882
rect 23204 17818 23256 17824
rect 22836 17332 22888 17338
rect 22836 17274 22888 17280
rect 23216 17270 23244 17818
rect 22744 17264 22796 17270
rect 22744 17206 22796 17212
rect 23204 17264 23256 17270
rect 23204 17206 23256 17212
rect 21364 17128 21416 17134
rect 21364 17070 21416 17076
rect 22192 17128 22244 17134
rect 22192 17070 22244 17076
rect 22836 17128 22888 17134
rect 22836 17070 22888 17076
rect 21272 14340 21324 14346
rect 21272 14282 21324 14288
rect 21180 13456 21232 13462
rect 21180 13398 21232 13404
rect 21376 13394 21404 17070
rect 22848 15570 22876 17070
rect 22836 15564 22888 15570
rect 22836 15506 22888 15512
rect 22284 15088 22336 15094
rect 22284 15030 22336 15036
rect 22100 15020 22152 15026
rect 22100 14962 22152 14968
rect 21824 14952 21876 14958
rect 21824 14894 21876 14900
rect 21836 14414 21864 14894
rect 22112 14618 22140 14962
rect 22296 14890 22324 15030
rect 22284 14884 22336 14890
rect 22284 14826 22336 14832
rect 22848 14634 22876 15506
rect 23020 15360 23072 15366
rect 23020 15302 23072 15308
rect 22100 14612 22152 14618
rect 22100 14554 22152 14560
rect 22756 14606 22876 14634
rect 22756 14550 22784 14606
rect 22744 14544 22796 14550
rect 22744 14486 22796 14492
rect 23032 14414 23060 15302
rect 23492 15178 23520 18158
rect 23572 18080 23624 18086
rect 23572 18022 23624 18028
rect 23584 16590 23612 18022
rect 23676 17134 23704 19654
rect 23848 18284 23900 18290
rect 23848 18226 23900 18232
rect 23756 17604 23808 17610
rect 23756 17546 23808 17552
rect 23664 17128 23716 17134
rect 23664 17070 23716 17076
rect 23572 16584 23624 16590
rect 23572 16526 23624 16532
rect 23676 16402 23704 17070
rect 23768 16794 23796 17546
rect 23860 17338 23888 18226
rect 23848 17332 23900 17338
rect 23848 17274 23900 17280
rect 23756 16788 23808 16794
rect 23756 16730 23808 16736
rect 23584 16374 23704 16402
rect 23584 15502 23612 16374
rect 23572 15496 23624 15502
rect 23572 15438 23624 15444
rect 23400 15150 23520 15178
rect 23400 14414 23428 15150
rect 21824 14408 21876 14414
rect 21824 14350 21876 14356
rect 23020 14408 23072 14414
rect 23020 14350 23072 14356
rect 23388 14408 23440 14414
rect 23388 14350 23440 14356
rect 21364 13388 21416 13394
rect 21364 13330 21416 13336
rect 20996 13184 21048 13190
rect 20996 13126 21048 13132
rect 21008 12850 21036 13126
rect 20812 12844 20864 12850
rect 20812 12786 20864 12792
rect 20996 12844 21048 12850
rect 20996 12786 21048 12792
rect 21836 12782 21864 14350
rect 23400 13938 23428 14350
rect 23296 13932 23348 13938
rect 23296 13874 23348 13880
rect 23388 13932 23440 13938
rect 23388 13874 23440 13880
rect 23020 13864 23072 13870
rect 23020 13806 23072 13812
rect 22008 13320 22060 13326
rect 22008 13262 22060 13268
rect 21824 12776 21876 12782
rect 21824 12718 21876 12724
rect 21088 12640 21140 12646
rect 21088 12582 21140 12588
rect 20720 12300 20772 12306
rect 20720 12242 20772 12248
rect 20732 11218 20760 12242
rect 21100 12238 21128 12582
rect 21836 12306 21864 12718
rect 21824 12300 21876 12306
rect 21824 12242 21876 12248
rect 21088 12232 21140 12238
rect 21088 12174 21140 12180
rect 22020 11830 22048 13262
rect 22100 12844 22152 12850
rect 22100 12786 22152 12792
rect 22112 12442 22140 12786
rect 22100 12436 22152 12442
rect 22100 12378 22152 12384
rect 22836 12164 22888 12170
rect 22836 12106 22888 12112
rect 22848 11898 22876 12106
rect 22836 11892 22888 11898
rect 22836 11834 22888 11840
rect 22008 11824 22060 11830
rect 22008 11766 22060 11772
rect 23032 11762 23060 13806
rect 23204 13184 23256 13190
rect 23204 13126 23256 13132
rect 23216 12986 23244 13126
rect 23204 12980 23256 12986
rect 23204 12922 23256 12928
rect 23308 11898 23336 13874
rect 23400 13326 23428 13874
rect 23388 13320 23440 13326
rect 23388 13262 23440 13268
rect 23584 13258 23612 15438
rect 23664 15360 23716 15366
rect 23664 15302 23716 15308
rect 23676 15162 23704 15302
rect 23664 15156 23716 15162
rect 23664 15098 23716 15104
rect 23572 13252 23624 13258
rect 23572 13194 23624 13200
rect 23848 12844 23900 12850
rect 23848 12786 23900 12792
rect 23860 12442 23888 12786
rect 23848 12436 23900 12442
rect 23848 12378 23900 12384
rect 23296 11892 23348 11898
rect 23296 11834 23348 11840
rect 23860 11830 23888 12378
rect 23952 11898 23980 25094
rect 24044 24274 24072 25230
rect 24110 24508 24418 24528
rect 24110 24506 24116 24508
rect 24172 24506 24196 24508
rect 24252 24506 24276 24508
rect 24332 24506 24356 24508
rect 24412 24506 24418 24508
rect 24172 24454 24174 24506
rect 24354 24454 24356 24506
rect 24110 24452 24116 24454
rect 24172 24452 24196 24454
rect 24252 24452 24276 24454
rect 24332 24452 24356 24454
rect 24412 24452 24418 24454
rect 24110 24432 24418 24452
rect 24032 24268 24084 24274
rect 24032 24210 24084 24216
rect 24110 23420 24418 23440
rect 24110 23418 24116 23420
rect 24172 23418 24196 23420
rect 24252 23418 24276 23420
rect 24332 23418 24356 23420
rect 24412 23418 24418 23420
rect 24172 23366 24174 23418
rect 24354 23366 24356 23418
rect 24110 23364 24116 23366
rect 24172 23364 24196 23366
rect 24252 23364 24276 23366
rect 24332 23364 24356 23366
rect 24412 23364 24418 23366
rect 24110 23344 24418 23364
rect 24688 23118 24716 25706
rect 24872 23118 24900 30670
rect 24964 25974 24992 31726
rect 25136 30592 25188 30598
rect 25136 30534 25188 30540
rect 25148 30258 25176 30534
rect 25136 30252 25188 30258
rect 25136 30194 25188 30200
rect 25688 29572 25740 29578
rect 25688 29514 25740 29520
rect 25042 29336 25098 29345
rect 25042 29271 25098 29280
rect 24952 25968 25004 25974
rect 24952 25910 25004 25916
rect 24952 25696 25004 25702
rect 24952 25638 25004 25644
rect 24964 25226 24992 25638
rect 24952 25220 25004 25226
rect 24952 25162 25004 25168
rect 25056 24818 25084 29271
rect 25136 26240 25188 26246
rect 25136 26182 25188 26188
rect 25148 25906 25176 26182
rect 25136 25900 25188 25906
rect 25136 25842 25188 25848
rect 25044 24812 25096 24818
rect 25044 24754 25096 24760
rect 25042 24168 25098 24177
rect 25042 24103 25044 24112
rect 25096 24103 25098 24112
rect 25596 24132 25648 24138
rect 25044 24074 25096 24080
rect 25596 24074 25648 24080
rect 25056 23474 25084 24074
rect 25608 23730 25636 24074
rect 25596 23724 25648 23730
rect 25596 23666 25648 23672
rect 25412 23656 25464 23662
rect 25412 23598 25464 23604
rect 24964 23446 25084 23474
rect 24676 23112 24728 23118
rect 24676 23054 24728 23060
rect 24860 23112 24912 23118
rect 24860 23054 24912 23060
rect 24676 22772 24728 22778
rect 24676 22714 24728 22720
rect 24110 22332 24418 22352
rect 24110 22330 24116 22332
rect 24172 22330 24196 22332
rect 24252 22330 24276 22332
rect 24332 22330 24356 22332
rect 24412 22330 24418 22332
rect 24172 22278 24174 22330
rect 24354 22278 24356 22330
rect 24110 22276 24116 22278
rect 24172 22276 24196 22278
rect 24252 22276 24276 22278
rect 24332 22276 24356 22278
rect 24412 22276 24418 22278
rect 24110 22256 24418 22276
rect 24584 22024 24636 22030
rect 24584 21966 24636 21972
rect 24110 21244 24418 21264
rect 24110 21242 24116 21244
rect 24172 21242 24196 21244
rect 24252 21242 24276 21244
rect 24332 21242 24356 21244
rect 24412 21242 24418 21244
rect 24172 21190 24174 21242
rect 24354 21190 24356 21242
rect 24110 21188 24116 21190
rect 24172 21188 24196 21190
rect 24252 21188 24276 21190
rect 24332 21188 24356 21190
rect 24412 21188 24418 21190
rect 24110 21168 24418 21188
rect 24492 20800 24544 20806
rect 24492 20742 24544 20748
rect 24110 20156 24418 20176
rect 24110 20154 24116 20156
rect 24172 20154 24196 20156
rect 24252 20154 24276 20156
rect 24332 20154 24356 20156
rect 24412 20154 24418 20156
rect 24172 20102 24174 20154
rect 24354 20102 24356 20154
rect 24110 20100 24116 20102
rect 24172 20100 24196 20102
rect 24252 20100 24276 20102
rect 24332 20100 24356 20102
rect 24412 20100 24418 20102
rect 24110 20080 24418 20100
rect 24032 19780 24084 19786
rect 24032 19722 24084 19728
rect 24044 19310 24072 19722
rect 24504 19378 24532 20742
rect 24492 19372 24544 19378
rect 24492 19314 24544 19320
rect 24032 19304 24084 19310
rect 24032 19246 24084 19252
rect 24044 18222 24072 19246
rect 24110 19068 24418 19088
rect 24110 19066 24116 19068
rect 24172 19066 24196 19068
rect 24252 19066 24276 19068
rect 24332 19066 24356 19068
rect 24412 19066 24418 19068
rect 24172 19014 24174 19066
rect 24354 19014 24356 19066
rect 24110 19012 24116 19014
rect 24172 19012 24196 19014
rect 24252 19012 24276 19014
rect 24332 19012 24356 19014
rect 24412 19012 24418 19014
rect 24110 18992 24418 19012
rect 24032 18216 24084 18222
rect 24032 18158 24084 18164
rect 24110 17980 24418 18000
rect 24110 17978 24116 17980
rect 24172 17978 24196 17980
rect 24252 17978 24276 17980
rect 24332 17978 24356 17980
rect 24412 17978 24418 17980
rect 24172 17926 24174 17978
rect 24354 17926 24356 17978
rect 24110 17924 24116 17926
rect 24172 17924 24196 17926
rect 24252 17924 24276 17926
rect 24332 17924 24356 17926
rect 24412 17924 24418 17926
rect 24110 17904 24418 17924
rect 24110 16892 24418 16912
rect 24110 16890 24116 16892
rect 24172 16890 24196 16892
rect 24252 16890 24276 16892
rect 24332 16890 24356 16892
rect 24412 16890 24418 16892
rect 24172 16838 24174 16890
rect 24354 16838 24356 16890
rect 24110 16836 24116 16838
rect 24172 16836 24196 16838
rect 24252 16836 24276 16838
rect 24332 16836 24356 16838
rect 24412 16836 24418 16838
rect 24110 16816 24418 16836
rect 24110 15804 24418 15824
rect 24110 15802 24116 15804
rect 24172 15802 24196 15804
rect 24252 15802 24276 15804
rect 24332 15802 24356 15804
rect 24412 15802 24418 15804
rect 24172 15750 24174 15802
rect 24354 15750 24356 15802
rect 24110 15748 24116 15750
rect 24172 15748 24196 15750
rect 24252 15748 24276 15750
rect 24332 15748 24356 15750
rect 24412 15748 24418 15750
rect 24110 15728 24418 15748
rect 24596 15706 24624 21966
rect 24584 15700 24636 15706
rect 24584 15642 24636 15648
rect 24124 15428 24176 15434
rect 24124 15370 24176 15376
rect 24136 15162 24164 15370
rect 24124 15156 24176 15162
rect 24124 15098 24176 15104
rect 24110 14716 24418 14736
rect 24110 14714 24116 14716
rect 24172 14714 24196 14716
rect 24252 14714 24276 14716
rect 24332 14714 24356 14716
rect 24412 14714 24418 14716
rect 24172 14662 24174 14714
rect 24354 14662 24356 14714
rect 24110 14660 24116 14662
rect 24172 14660 24196 14662
rect 24252 14660 24276 14662
rect 24332 14660 24356 14662
rect 24412 14660 24418 14662
rect 24110 14640 24418 14660
rect 24688 14482 24716 22714
rect 24872 21418 24900 23054
rect 24860 21412 24912 21418
rect 24860 21354 24912 21360
rect 24964 20482 24992 23446
rect 25228 23248 25280 23254
rect 25228 23190 25280 23196
rect 25136 22976 25188 22982
rect 25136 22918 25188 22924
rect 25148 22778 25176 22918
rect 25136 22772 25188 22778
rect 25136 22714 25188 22720
rect 25044 22636 25096 22642
rect 25044 22578 25096 22584
rect 25056 22234 25084 22578
rect 25044 22228 25096 22234
rect 25044 22170 25096 22176
rect 25148 22094 25176 22714
rect 24872 20454 24992 20482
rect 25056 22066 25176 22094
rect 24872 18902 24900 20454
rect 24952 20392 25004 20398
rect 24952 20334 25004 20340
rect 24860 18896 24912 18902
rect 24860 18838 24912 18844
rect 24872 17610 24900 18838
rect 24964 18222 24992 20334
rect 24952 18216 25004 18222
rect 24952 18158 25004 18164
rect 24860 17604 24912 17610
rect 24860 17546 24912 17552
rect 24860 15496 24912 15502
rect 24860 15438 24912 15444
rect 24768 15156 24820 15162
rect 24768 15098 24820 15104
rect 24492 14476 24544 14482
rect 24492 14418 24544 14424
rect 24676 14476 24728 14482
rect 24676 14418 24728 14424
rect 24110 13628 24418 13648
rect 24110 13626 24116 13628
rect 24172 13626 24196 13628
rect 24252 13626 24276 13628
rect 24332 13626 24356 13628
rect 24412 13626 24418 13628
rect 24172 13574 24174 13626
rect 24354 13574 24356 13626
rect 24110 13572 24116 13574
rect 24172 13572 24196 13574
rect 24252 13572 24276 13574
rect 24332 13572 24356 13574
rect 24412 13572 24418 13574
rect 24110 13552 24418 13572
rect 24032 13252 24084 13258
rect 24032 13194 24084 13200
rect 23940 11892 23992 11898
rect 23940 11834 23992 11840
rect 23848 11824 23900 11830
rect 23848 11766 23900 11772
rect 20904 11756 20956 11762
rect 20904 11698 20956 11704
rect 23020 11756 23072 11762
rect 23020 11698 23072 11704
rect 20720 11212 20772 11218
rect 20720 11154 20772 11160
rect 20916 10810 20944 11698
rect 24044 11694 24072 13194
rect 24504 12782 24532 14418
rect 24780 14414 24808 15098
rect 24872 15065 24900 15438
rect 24858 15056 24914 15065
rect 24858 14991 24914 15000
rect 24860 14816 24912 14822
rect 24860 14758 24912 14764
rect 24768 14408 24820 14414
rect 24768 14350 24820 14356
rect 24676 13320 24728 13326
rect 24676 13262 24728 13268
rect 24688 12986 24716 13262
rect 24676 12980 24728 12986
rect 24676 12922 24728 12928
rect 24492 12776 24544 12782
rect 24492 12718 24544 12724
rect 24110 12540 24418 12560
rect 24110 12538 24116 12540
rect 24172 12538 24196 12540
rect 24252 12538 24276 12540
rect 24332 12538 24356 12540
rect 24412 12538 24418 12540
rect 24172 12486 24174 12538
rect 24354 12486 24356 12538
rect 24110 12484 24116 12486
rect 24172 12484 24196 12486
rect 24252 12484 24276 12486
rect 24332 12484 24356 12486
rect 24412 12484 24418 12486
rect 24110 12464 24418 12484
rect 24872 11778 24900 14758
rect 24964 14550 24992 18158
rect 24952 14544 25004 14550
rect 24952 14486 25004 14492
rect 24952 12164 25004 12170
rect 24952 12106 25004 12112
rect 24964 11898 24992 12106
rect 24952 11892 25004 11898
rect 24952 11834 25004 11840
rect 24872 11750 24992 11778
rect 25056 11762 25084 22066
rect 25240 22030 25268 23190
rect 25228 22024 25280 22030
rect 25228 21966 25280 21972
rect 25320 22024 25372 22030
rect 25320 21966 25372 21972
rect 25332 21010 25360 21966
rect 25320 21004 25372 21010
rect 25320 20946 25372 20952
rect 25136 20800 25188 20806
rect 25136 20742 25188 20748
rect 25148 20058 25176 20742
rect 25424 20346 25452 23598
rect 25608 23118 25636 23666
rect 25596 23112 25648 23118
rect 25596 23054 25648 23060
rect 25504 22160 25556 22166
rect 25504 22102 25556 22108
rect 25516 21010 25544 22102
rect 25504 21004 25556 21010
rect 25504 20946 25556 20952
rect 25700 20398 25728 29514
rect 25778 26616 25834 26625
rect 25778 26551 25834 26560
rect 25332 20318 25452 20346
rect 25688 20392 25740 20398
rect 25688 20334 25740 20340
rect 25136 20052 25188 20058
rect 25136 19994 25188 20000
rect 25148 19938 25176 19994
rect 25148 19910 25268 19938
rect 25136 19780 25188 19786
rect 25136 19722 25188 19728
rect 25148 19514 25176 19722
rect 25136 19508 25188 19514
rect 25136 19450 25188 19456
rect 25240 18426 25268 19910
rect 25228 18420 25280 18426
rect 25228 18362 25280 18368
rect 25332 15994 25360 20318
rect 25412 20256 25464 20262
rect 25412 20198 25464 20204
rect 25240 15966 25360 15994
rect 25240 15609 25268 15966
rect 25226 15600 25282 15609
rect 25226 15535 25282 15544
rect 25136 14952 25188 14958
rect 25136 14894 25188 14900
rect 25148 14618 25176 14894
rect 25240 14822 25268 15535
rect 25320 15428 25372 15434
rect 25320 15370 25372 15376
rect 25332 15094 25360 15370
rect 25320 15088 25372 15094
rect 25320 15030 25372 15036
rect 25228 14816 25280 14822
rect 25228 14758 25280 14764
rect 25136 14612 25188 14618
rect 25136 14554 25188 14560
rect 25148 14074 25176 14554
rect 25136 14068 25188 14074
rect 25136 14010 25188 14016
rect 25424 13938 25452 20198
rect 25596 18284 25648 18290
rect 25596 18226 25648 18232
rect 25504 18080 25556 18086
rect 25504 18022 25556 18028
rect 25516 16590 25544 18022
rect 25608 17542 25636 18226
rect 25596 17536 25648 17542
rect 25596 17478 25648 17484
rect 25608 17202 25636 17478
rect 25596 17196 25648 17202
rect 25596 17138 25648 17144
rect 25792 16590 25820 26551
rect 25884 23186 25912 35566
rect 25962 32736 26018 32745
rect 25962 32671 26018 32680
rect 25976 32366 26004 32671
rect 25964 32360 26016 32366
rect 25964 32302 26016 32308
rect 25964 24744 26016 24750
rect 25964 24686 26016 24692
rect 25976 24585 26004 24686
rect 25962 24576 26018 24585
rect 25962 24511 26018 24520
rect 25872 23180 25924 23186
rect 25872 23122 25924 23128
rect 25964 22500 26016 22506
rect 25964 22442 26016 22448
rect 25976 21622 26004 22442
rect 25964 21616 26016 21622
rect 25964 21558 26016 21564
rect 26068 17814 26096 42191
rect 26424 42016 26476 42022
rect 26424 41958 26476 41964
rect 26436 41138 26464 41958
rect 26424 41132 26476 41138
rect 26424 41074 26476 41080
rect 26332 39840 26384 39846
rect 26332 39782 26384 39788
rect 26344 39506 26372 39782
rect 26332 39500 26384 39506
rect 26332 39442 26384 39448
rect 26516 39364 26568 39370
rect 26516 39306 26568 39312
rect 26528 39098 26556 39306
rect 26516 39092 26568 39098
rect 26516 39034 26568 39040
rect 26332 38752 26384 38758
rect 26332 38694 26384 38700
rect 26344 38418 26372 38694
rect 26332 38412 26384 38418
rect 26332 38354 26384 38360
rect 26792 37256 26844 37262
rect 26792 37198 26844 37204
rect 26608 37120 26660 37126
rect 26608 37062 26660 37068
rect 26332 35488 26384 35494
rect 26332 35430 26384 35436
rect 26344 34610 26372 35430
rect 26620 35086 26648 37062
rect 26804 36825 26832 37198
rect 26790 36816 26846 36825
rect 26790 36751 26846 36760
rect 26792 36168 26844 36174
rect 26792 36110 26844 36116
rect 26608 35080 26660 35086
rect 26608 35022 26660 35028
rect 26332 34604 26384 34610
rect 26332 34546 26384 34552
rect 26240 33312 26292 33318
rect 26240 33254 26292 33260
rect 26332 33312 26384 33318
rect 26332 33254 26384 33260
rect 26252 32366 26280 33254
rect 26344 32978 26372 33254
rect 26332 32972 26384 32978
rect 26332 32914 26384 32920
rect 26240 32360 26292 32366
rect 26240 32302 26292 32308
rect 26148 30728 26200 30734
rect 26148 30670 26200 30676
rect 26160 30054 26188 30670
rect 26148 30048 26200 30054
rect 26148 29990 26200 29996
rect 26516 30048 26568 30054
rect 26516 29990 26568 29996
rect 26160 29578 26188 29990
rect 26528 29714 26556 29990
rect 26516 29708 26568 29714
rect 26516 29650 26568 29656
rect 26148 29572 26200 29578
rect 26148 29514 26200 29520
rect 26424 26376 26476 26382
rect 26424 26318 26476 26324
rect 26436 24818 26464 26318
rect 26804 24818 26832 36110
rect 26896 26058 26924 45766
rect 26988 33522 27016 46038
rect 27528 45892 27580 45898
rect 27528 45834 27580 45840
rect 27436 45824 27488 45830
rect 27436 45766 27488 45772
rect 27448 45490 27476 45766
rect 27540 45558 27568 45834
rect 27528 45552 27580 45558
rect 27528 45494 27580 45500
rect 27436 45484 27488 45490
rect 27436 45426 27488 45432
rect 27436 45008 27488 45014
rect 27436 44950 27488 44956
rect 27526 44976 27582 44985
rect 27448 44402 27476 44950
rect 27908 44946 27936 46310
rect 27526 44911 27528 44920
rect 27580 44911 27582 44920
rect 27896 44940 27948 44946
rect 27528 44882 27580 44888
rect 27896 44882 27948 44888
rect 27620 44804 27672 44810
rect 27620 44746 27672 44752
rect 27632 44538 27660 44746
rect 27620 44532 27672 44538
rect 27620 44474 27672 44480
rect 27436 44396 27488 44402
rect 27436 44338 27488 44344
rect 27068 43716 27120 43722
rect 27068 43658 27120 43664
rect 27080 43450 27108 43658
rect 27068 43444 27120 43450
rect 27068 43386 27120 43392
rect 27068 42016 27120 42022
rect 27068 41958 27120 41964
rect 27080 41682 27108 41958
rect 27068 41676 27120 41682
rect 27068 41618 27120 41624
rect 27344 41132 27396 41138
rect 27344 41074 27396 41080
rect 27356 40118 27384 41074
rect 27344 40112 27396 40118
rect 27344 40054 27396 40060
rect 27252 35692 27304 35698
rect 27252 35634 27304 35640
rect 27264 35290 27292 35634
rect 27252 35284 27304 35290
rect 27252 35226 27304 35232
rect 27160 33924 27212 33930
rect 27160 33866 27212 33872
rect 27172 33658 27200 33866
rect 27160 33652 27212 33658
rect 27160 33594 27212 33600
rect 26976 33516 27028 33522
rect 26976 33458 27028 33464
rect 26988 33402 27016 33458
rect 26988 33374 27108 33402
rect 26976 33040 27028 33046
rect 26976 32982 27028 32988
rect 26988 32434 27016 32982
rect 26976 32428 27028 32434
rect 26976 32370 27028 32376
rect 26988 30258 27016 32370
rect 26976 30252 27028 30258
rect 26976 30194 27028 30200
rect 26896 26030 27016 26058
rect 26884 25968 26936 25974
rect 26884 25910 26936 25916
rect 26424 24812 26476 24818
rect 26424 24754 26476 24760
rect 26792 24812 26844 24818
rect 26792 24754 26844 24760
rect 26240 22432 26292 22438
rect 26240 22374 26292 22380
rect 26516 22432 26568 22438
rect 26516 22374 26568 22380
rect 26252 22166 26280 22374
rect 26240 22160 26292 22166
rect 26240 22102 26292 22108
rect 26148 21480 26200 21486
rect 26148 21422 26200 21428
rect 26160 21185 26188 21422
rect 26146 21176 26202 21185
rect 26146 21111 26202 21120
rect 26252 20754 26280 22102
rect 26528 22098 26556 22374
rect 26516 22092 26568 22098
rect 26896 22094 26924 25910
rect 26988 23322 27016 26030
rect 27080 23662 27108 33374
rect 27252 32224 27304 32230
rect 27252 32166 27304 32172
rect 27264 31890 27292 32166
rect 27252 31884 27304 31890
rect 27252 31826 27304 31832
rect 27356 31754 27384 40054
rect 27448 34950 27476 44338
rect 28000 43858 28028 49286
rect 28326 49200 28438 50000
rect 28970 49200 29082 50000
rect 29614 49200 29726 50000
rect 28368 47122 28396 49200
rect 28356 47116 28408 47122
rect 28356 47058 28408 47064
rect 28172 47048 28224 47054
rect 28172 46990 28224 46996
rect 28814 47016 28870 47025
rect 28080 46912 28132 46918
rect 28080 46854 28132 46860
rect 27988 43852 28040 43858
rect 27988 43794 28040 43800
rect 27712 42560 27764 42566
rect 27712 42502 27764 42508
rect 27724 42226 27752 42502
rect 27712 42220 27764 42226
rect 27712 42162 27764 42168
rect 27526 40896 27582 40905
rect 27526 40831 27582 40840
rect 27540 40594 27568 40831
rect 27528 40588 27580 40594
rect 27528 40530 27580 40536
rect 27620 40384 27672 40390
rect 27620 40326 27672 40332
rect 27632 36786 27660 40326
rect 27724 40050 27752 42162
rect 27804 42016 27856 42022
rect 27804 41958 27856 41964
rect 27816 41546 27844 41958
rect 27804 41540 27856 41546
rect 27804 41482 27856 41488
rect 27988 40452 28040 40458
rect 27988 40394 28040 40400
rect 28000 40186 28028 40394
rect 27988 40180 28040 40186
rect 27988 40122 28040 40128
rect 27712 40044 27764 40050
rect 27712 39986 27764 39992
rect 27804 38956 27856 38962
rect 27804 38898 27856 38904
rect 27712 38276 27764 38282
rect 27712 38218 27764 38224
rect 27724 38010 27752 38218
rect 27712 38004 27764 38010
rect 27712 37946 27764 37952
rect 27712 37868 27764 37874
rect 27712 37810 27764 37816
rect 27620 36780 27672 36786
rect 27620 36722 27672 36728
rect 27528 36236 27580 36242
rect 27528 36178 27580 36184
rect 27540 36145 27568 36178
rect 27526 36136 27582 36145
rect 27526 36071 27582 36080
rect 27436 34944 27488 34950
rect 27436 34886 27488 34892
rect 27436 34672 27488 34678
rect 27434 34640 27436 34649
rect 27488 34640 27490 34649
rect 27434 34575 27490 34584
rect 27526 34096 27582 34105
rect 27526 34031 27528 34040
rect 27580 34031 27582 34040
rect 27528 34002 27580 34008
rect 27632 33590 27660 36722
rect 27724 35630 27752 37810
rect 27712 35624 27764 35630
rect 27712 35566 27764 35572
rect 27712 35080 27764 35086
rect 27712 35022 27764 35028
rect 27724 34610 27752 35022
rect 27816 35018 27844 38898
rect 27896 37324 27948 37330
rect 27896 37266 27948 37272
rect 27908 36310 27936 37266
rect 27988 36576 28040 36582
rect 27988 36518 28040 36524
rect 27896 36304 27948 36310
rect 27896 36246 27948 36252
rect 28000 36242 28028 36518
rect 27988 36236 28040 36242
rect 27988 36178 28040 36184
rect 27804 35012 27856 35018
rect 27804 34954 27856 34960
rect 27712 34604 27764 34610
rect 27712 34546 27764 34552
rect 27620 33584 27672 33590
rect 27620 33526 27672 33532
rect 27724 33522 27752 34546
rect 27896 33584 27948 33590
rect 27896 33526 27948 33532
rect 27712 33516 27764 33522
rect 27712 33458 27764 33464
rect 27436 31816 27488 31822
rect 27436 31758 27488 31764
rect 27264 31726 27384 31754
rect 27264 28082 27292 31726
rect 27342 30016 27398 30025
rect 27342 29951 27398 29960
rect 27356 29170 27384 29951
rect 27344 29164 27396 29170
rect 27344 29106 27396 29112
rect 27344 28484 27396 28490
rect 27344 28426 27396 28432
rect 27356 28218 27384 28426
rect 27344 28212 27396 28218
rect 27344 28154 27396 28160
rect 27252 28076 27304 28082
rect 27252 28018 27304 28024
rect 27448 26874 27476 31758
rect 27908 31754 27936 33526
rect 28092 32978 28120 46854
rect 28184 46034 28212 46990
rect 28814 46951 28870 46960
rect 28172 46028 28224 46034
rect 28172 45970 28224 45976
rect 28264 43308 28316 43314
rect 28264 43250 28316 43256
rect 28170 42936 28226 42945
rect 28170 42871 28226 42880
rect 28184 41682 28212 42871
rect 28172 41676 28224 41682
rect 28172 41618 28224 41624
rect 28172 40928 28224 40934
rect 28172 40870 28224 40876
rect 28184 40594 28212 40870
rect 28172 40588 28224 40594
rect 28172 40530 28224 40536
rect 28170 40216 28226 40225
rect 28170 40151 28226 40160
rect 28184 39506 28212 40151
rect 28172 39500 28224 39506
rect 28172 39442 28224 39448
rect 28276 38962 28304 43250
rect 28828 42770 28856 46951
rect 28816 42764 28868 42770
rect 28816 42706 28868 42712
rect 28722 39536 28778 39545
rect 28722 39471 28778 39480
rect 28264 38956 28316 38962
rect 28264 38898 28316 38904
rect 28736 38418 28764 39471
rect 28724 38412 28776 38418
rect 28724 38354 28776 38360
rect 28172 37324 28224 37330
rect 28172 37266 28224 37272
rect 28184 34066 28212 37266
rect 28816 35012 28868 35018
rect 28816 34954 28868 34960
rect 28172 34060 28224 34066
rect 28172 34002 28224 34008
rect 28080 32972 28132 32978
rect 28080 32914 28132 32920
rect 28448 32428 28500 32434
rect 28448 32370 28500 32376
rect 28172 31816 28224 31822
rect 28172 31758 28224 31764
rect 27816 31726 27936 31754
rect 27816 31346 27844 31726
rect 27804 31340 27856 31346
rect 27804 31282 27856 31288
rect 27528 30796 27580 30802
rect 27528 30738 27580 30744
rect 27540 30705 27568 30738
rect 27526 30696 27582 30705
rect 27526 30631 27582 30640
rect 27816 30258 27844 31282
rect 27988 31136 28040 31142
rect 27988 31078 28040 31084
rect 28000 30802 28028 31078
rect 28184 30802 28212 31758
rect 27988 30796 28040 30802
rect 27988 30738 28040 30744
rect 28172 30796 28224 30802
rect 28172 30738 28224 30744
rect 27620 30252 27672 30258
rect 27620 30194 27672 30200
rect 27804 30252 27856 30258
rect 27804 30194 27856 30200
rect 27526 28656 27582 28665
rect 27526 28591 27528 28600
rect 27580 28591 27582 28600
rect 27528 28562 27580 28568
rect 27528 27532 27580 27538
rect 27528 27474 27580 27480
rect 27540 27305 27568 27474
rect 27526 27296 27582 27305
rect 27526 27231 27582 27240
rect 27172 26846 27476 26874
rect 27068 23656 27120 23662
rect 27068 23598 27120 23604
rect 26976 23316 27028 23322
rect 26976 23258 27028 23264
rect 26988 23118 27016 23258
rect 26976 23112 27028 23118
rect 26976 23054 27028 23060
rect 26516 22034 26568 22040
rect 26804 22066 26924 22094
rect 26516 21344 26568 21350
rect 26516 21286 26568 21292
rect 26528 21010 26556 21286
rect 26516 21004 26568 21010
rect 26516 20946 26568 20952
rect 26160 20726 26280 20754
rect 26160 20602 26188 20726
rect 26148 20596 26200 20602
rect 26148 20538 26200 20544
rect 26516 20256 26568 20262
rect 26516 20198 26568 20204
rect 26528 19922 26556 20198
rect 26516 19916 26568 19922
rect 26516 19858 26568 19864
rect 26332 19848 26384 19854
rect 26332 19790 26384 19796
rect 26344 19378 26372 19790
rect 26332 19372 26384 19378
rect 26332 19314 26384 19320
rect 26516 18080 26568 18086
rect 26516 18022 26568 18028
rect 26056 17808 26108 17814
rect 26056 17750 26108 17756
rect 26528 17746 26556 18022
rect 26516 17740 26568 17746
rect 26516 17682 26568 17688
rect 26332 17672 26384 17678
rect 26332 17614 26384 17620
rect 26344 17338 26372 17614
rect 26332 17332 26384 17338
rect 26332 17274 26384 17280
rect 25872 17196 25924 17202
rect 25872 17138 25924 17144
rect 26240 17196 26292 17202
rect 26240 17138 26292 17144
rect 25504 16584 25556 16590
rect 25504 16526 25556 16532
rect 25688 16584 25740 16590
rect 25688 16526 25740 16532
rect 25780 16584 25832 16590
rect 25780 16526 25832 16532
rect 25412 13932 25464 13938
rect 25412 13874 25464 13880
rect 25228 13320 25280 13326
rect 25228 13262 25280 13268
rect 25240 11830 25268 13262
rect 25424 12850 25452 13874
rect 25516 13870 25544 16526
rect 25700 16130 25728 16526
rect 25884 16182 25912 17138
rect 25872 16176 25924 16182
rect 25700 16114 25820 16130
rect 25872 16118 25924 16124
rect 26252 16114 26280 17138
rect 26332 17128 26384 17134
rect 26332 17070 26384 17076
rect 26344 16998 26372 17070
rect 26332 16992 26384 16998
rect 26332 16934 26384 16940
rect 26344 16726 26372 16934
rect 26332 16720 26384 16726
rect 26332 16662 26384 16668
rect 25700 16108 25832 16114
rect 25700 16102 25780 16108
rect 25780 16050 25832 16056
rect 26240 16108 26292 16114
rect 26240 16050 26292 16056
rect 25688 15564 25740 15570
rect 25688 15506 25740 15512
rect 25596 15088 25648 15094
rect 25596 15030 25648 15036
rect 25608 14414 25636 15030
rect 25596 14408 25648 14414
rect 25596 14350 25648 14356
rect 25608 14074 25636 14350
rect 25596 14068 25648 14074
rect 25596 14010 25648 14016
rect 25504 13864 25556 13870
rect 25504 13806 25556 13812
rect 25516 13326 25544 13806
rect 25700 13802 25728 15506
rect 25792 14958 25820 16050
rect 25872 16040 25924 16046
rect 25872 15982 25924 15988
rect 25884 15366 25912 15982
rect 26056 15972 26108 15978
rect 26056 15914 26108 15920
rect 26068 15570 26096 15914
rect 26148 15904 26200 15910
rect 26148 15846 26200 15852
rect 26056 15564 26108 15570
rect 26056 15506 26108 15512
rect 25872 15360 25924 15366
rect 25872 15302 25924 15308
rect 25780 14952 25832 14958
rect 25780 14894 25832 14900
rect 25884 14414 25912 15302
rect 25872 14408 25924 14414
rect 25872 14350 25924 14356
rect 25780 14272 25832 14278
rect 25780 14214 25832 14220
rect 25688 13796 25740 13802
rect 25688 13738 25740 13744
rect 25700 13530 25728 13738
rect 25792 13530 25820 14214
rect 25884 14006 25912 14350
rect 25872 14000 25924 14006
rect 25872 13942 25924 13948
rect 25688 13524 25740 13530
rect 25688 13466 25740 13472
rect 25780 13524 25832 13530
rect 25780 13466 25832 13472
rect 25504 13320 25556 13326
rect 25504 13262 25556 13268
rect 25412 12844 25464 12850
rect 25412 12786 25464 12792
rect 25688 12844 25740 12850
rect 25688 12786 25740 12792
rect 25700 11830 25728 12786
rect 25792 12434 25820 13466
rect 25884 12850 25912 13942
rect 25964 13728 26016 13734
rect 25964 13670 26016 13676
rect 25976 13394 26004 13670
rect 25964 13388 26016 13394
rect 25964 13330 26016 13336
rect 25872 12844 25924 12850
rect 25872 12786 25924 12792
rect 25976 12782 26004 13330
rect 25964 12776 26016 12782
rect 25964 12718 26016 12724
rect 25792 12406 25912 12434
rect 25884 12102 25912 12406
rect 26160 12306 26188 15846
rect 26252 15162 26280 16050
rect 26344 15434 26372 16662
rect 26608 15904 26660 15910
rect 26608 15846 26660 15852
rect 26332 15428 26384 15434
rect 26332 15370 26384 15376
rect 26516 15428 26568 15434
rect 26516 15370 26568 15376
rect 26240 15156 26292 15162
rect 26240 15098 26292 15104
rect 26344 14958 26372 15370
rect 26424 15360 26476 15366
rect 26424 15302 26476 15308
rect 26436 15026 26464 15302
rect 26528 15162 26556 15370
rect 26516 15156 26568 15162
rect 26516 15098 26568 15104
rect 26424 15020 26476 15026
rect 26424 14962 26476 14968
rect 26332 14952 26384 14958
rect 26332 14894 26384 14900
rect 26240 13320 26292 13326
rect 26240 13262 26292 13268
rect 26148 12300 26200 12306
rect 26148 12242 26200 12248
rect 25872 12096 25924 12102
rect 25872 12038 25924 12044
rect 25228 11824 25280 11830
rect 25228 11766 25280 11772
rect 25688 11824 25740 11830
rect 25688 11766 25740 11772
rect 24032 11688 24084 11694
rect 24032 11630 24084 11636
rect 21364 11552 21416 11558
rect 21364 11494 21416 11500
rect 21376 11150 21404 11494
rect 24110 11452 24418 11472
rect 24110 11450 24116 11452
rect 24172 11450 24196 11452
rect 24252 11450 24276 11452
rect 24332 11450 24356 11452
rect 24412 11450 24418 11452
rect 24172 11398 24174 11450
rect 24354 11398 24356 11450
rect 24110 11396 24116 11398
rect 24172 11396 24196 11398
rect 24252 11396 24276 11398
rect 24332 11396 24356 11398
rect 24412 11396 24418 11398
rect 24110 11376 24418 11396
rect 21364 11144 21416 11150
rect 21364 11086 21416 11092
rect 20904 10804 20956 10810
rect 20904 10746 20956 10752
rect 20260 10600 20312 10606
rect 20260 10542 20312 10548
rect 20444 10600 20496 10606
rect 20444 10542 20496 10548
rect 20272 10130 20300 10542
rect 20260 10124 20312 10130
rect 20260 10066 20312 10072
rect 19478 9820 19786 9840
rect 19478 9818 19484 9820
rect 19540 9818 19564 9820
rect 19620 9818 19644 9820
rect 19700 9818 19724 9820
rect 19780 9818 19786 9820
rect 19540 9766 19542 9818
rect 19722 9766 19724 9818
rect 19478 9764 19484 9766
rect 19540 9764 19564 9766
rect 19620 9764 19644 9766
rect 19700 9764 19724 9766
rect 19780 9764 19786 9766
rect 19478 9744 19786 9764
rect 19478 8732 19786 8752
rect 19478 8730 19484 8732
rect 19540 8730 19564 8732
rect 19620 8730 19644 8732
rect 19700 8730 19724 8732
rect 19780 8730 19786 8732
rect 19540 8678 19542 8730
rect 19722 8678 19724 8730
rect 19478 8676 19484 8678
rect 19540 8676 19564 8678
rect 19620 8676 19644 8678
rect 19700 8676 19724 8678
rect 19780 8676 19786 8678
rect 19478 8656 19786 8676
rect 18694 7984 18750 7993
rect 18694 7919 18750 7928
rect 18708 7886 18736 7919
rect 18696 7880 18748 7886
rect 18696 7822 18748 7828
rect 19478 7644 19786 7664
rect 19478 7642 19484 7644
rect 19540 7642 19564 7644
rect 19620 7642 19644 7644
rect 19700 7642 19724 7644
rect 19780 7642 19786 7644
rect 19540 7590 19542 7642
rect 19722 7590 19724 7642
rect 19478 7588 19484 7590
rect 19540 7588 19564 7590
rect 19620 7588 19644 7590
rect 19700 7588 19724 7590
rect 19780 7588 19786 7590
rect 19478 7568 19786 7588
rect 19478 6556 19786 6576
rect 19478 6554 19484 6556
rect 19540 6554 19564 6556
rect 19620 6554 19644 6556
rect 19700 6554 19724 6556
rect 19780 6554 19786 6556
rect 19540 6502 19542 6554
rect 19722 6502 19724 6554
rect 19478 6500 19484 6502
rect 19540 6500 19564 6502
rect 19620 6500 19644 6502
rect 19700 6500 19724 6502
rect 19780 6500 19786 6502
rect 19478 6480 19786 6500
rect 18604 5704 18656 5710
rect 18604 5646 18656 5652
rect 18616 5234 18644 5646
rect 19478 5468 19786 5488
rect 19478 5466 19484 5468
rect 19540 5466 19564 5468
rect 19620 5466 19644 5468
rect 19700 5466 19724 5468
rect 19780 5466 19786 5468
rect 19540 5414 19542 5466
rect 19722 5414 19724 5466
rect 19478 5412 19484 5414
rect 19540 5412 19564 5414
rect 19620 5412 19644 5414
rect 19700 5412 19724 5414
rect 19780 5412 19786 5414
rect 19478 5392 19786 5412
rect 18604 5228 18656 5234
rect 18604 5170 18656 5176
rect 19340 5160 19392 5166
rect 19340 5102 19392 5108
rect 19352 4264 19380 5102
rect 19478 4380 19786 4400
rect 19478 4378 19484 4380
rect 19540 4378 19564 4380
rect 19620 4378 19644 4380
rect 19700 4378 19724 4380
rect 19780 4378 19786 4380
rect 19540 4326 19542 4378
rect 19722 4326 19724 4378
rect 19478 4324 19484 4326
rect 19540 4324 19564 4326
rect 19620 4324 19644 4326
rect 19700 4324 19724 4326
rect 19780 4324 19786 4326
rect 19478 4304 19786 4324
rect 19352 4236 19472 4264
rect 18052 4072 18104 4078
rect 18052 4014 18104 4020
rect 18236 4072 18288 4078
rect 18236 4014 18288 4020
rect 16856 2644 16908 2650
rect 16856 2586 16908 2592
rect 17500 2644 17552 2650
rect 17500 2586 17552 2592
rect 17408 2440 17460 2446
rect 17408 2382 17460 2388
rect 17420 800 17448 2382
rect 18064 800 18092 4014
rect 19294 3596 19346 3602
rect 19444 3584 19472 4236
rect 19616 4072 19668 4078
rect 19616 4014 19668 4020
rect 19892 4072 19944 4078
rect 19892 4014 19944 4020
rect 19346 3556 19472 3584
rect 19294 3538 19346 3544
rect 19628 3534 19656 4014
rect 19904 3738 19932 4014
rect 19984 3936 20036 3942
rect 19984 3878 20036 3884
rect 19892 3732 19944 3738
rect 19892 3674 19944 3680
rect 19616 3528 19668 3534
rect 19616 3470 19668 3476
rect 19340 3392 19392 3398
rect 19340 3334 19392 3340
rect 19352 3126 19380 3334
rect 19478 3292 19786 3312
rect 19478 3290 19484 3292
rect 19540 3290 19564 3292
rect 19620 3290 19644 3292
rect 19700 3290 19724 3292
rect 19780 3290 19786 3292
rect 19540 3238 19542 3290
rect 19722 3238 19724 3290
rect 19478 3236 19484 3238
rect 19540 3236 19564 3238
rect 19620 3236 19644 3238
rect 19700 3236 19724 3238
rect 19780 3236 19786 3238
rect 19478 3216 19786 3236
rect 19996 3194 20024 3878
rect 19984 3188 20036 3194
rect 19984 3130 20036 3136
rect 19340 3120 19392 3126
rect 19340 3062 19392 3068
rect 19432 2984 19484 2990
rect 19432 2926 19484 2932
rect 19984 2984 20036 2990
rect 19984 2926 20036 2932
rect 19444 2650 19472 2926
rect 19432 2644 19484 2650
rect 19432 2586 19484 2592
rect 19478 2204 19786 2224
rect 19478 2202 19484 2204
rect 19540 2202 19564 2204
rect 19620 2202 19644 2204
rect 19700 2202 19724 2204
rect 19780 2202 19786 2204
rect 19540 2150 19542 2202
rect 19722 2150 19724 2202
rect 19478 2148 19484 2150
rect 19540 2148 19564 2150
rect 19620 2148 19644 2150
rect 19700 2148 19724 2150
rect 19780 2148 19786 2150
rect 19478 2128 19786 2148
rect 19996 800 20024 2926
rect 20456 2650 20484 10542
rect 24110 10364 24418 10384
rect 24110 10362 24116 10364
rect 24172 10362 24196 10364
rect 24252 10362 24276 10364
rect 24332 10362 24356 10364
rect 24412 10362 24418 10364
rect 24172 10310 24174 10362
rect 24354 10310 24356 10362
rect 24110 10308 24116 10310
rect 24172 10308 24196 10310
rect 24252 10308 24276 10310
rect 24332 10308 24356 10310
rect 24412 10308 24418 10310
rect 24110 10288 24418 10308
rect 24860 9512 24912 9518
rect 24860 9454 24912 9460
rect 24110 9276 24418 9296
rect 24110 9274 24116 9276
rect 24172 9274 24196 9276
rect 24252 9274 24276 9276
rect 24332 9274 24356 9276
rect 24412 9274 24418 9276
rect 24172 9222 24174 9274
rect 24354 9222 24356 9274
rect 24110 9220 24116 9222
rect 24172 9220 24196 9222
rect 24252 9220 24276 9222
rect 24332 9220 24356 9222
rect 24412 9220 24418 9222
rect 24110 9200 24418 9220
rect 24584 8968 24636 8974
rect 24584 8910 24636 8916
rect 24110 8188 24418 8208
rect 24110 8186 24116 8188
rect 24172 8186 24196 8188
rect 24252 8186 24276 8188
rect 24332 8186 24356 8188
rect 24412 8186 24418 8188
rect 24172 8134 24174 8186
rect 24354 8134 24356 8186
rect 24110 8132 24116 8134
rect 24172 8132 24196 8134
rect 24252 8132 24276 8134
rect 24332 8132 24356 8134
rect 24412 8132 24418 8134
rect 24110 8112 24418 8132
rect 24596 7410 24624 8910
rect 24584 7404 24636 7410
rect 24584 7346 24636 7352
rect 24110 7100 24418 7120
rect 24110 7098 24116 7100
rect 24172 7098 24196 7100
rect 24252 7098 24276 7100
rect 24332 7098 24356 7100
rect 24412 7098 24418 7100
rect 24172 7046 24174 7098
rect 24354 7046 24356 7098
rect 24110 7044 24116 7046
rect 24172 7044 24196 7046
rect 24252 7044 24276 7046
rect 24332 7044 24356 7046
rect 24412 7044 24418 7046
rect 24110 7024 24418 7044
rect 24872 6866 24900 9454
rect 24964 6914 24992 11750
rect 25044 11756 25096 11762
rect 25044 11698 25096 11704
rect 25056 10062 25084 11698
rect 26252 11354 26280 13262
rect 26332 12368 26384 12374
rect 26332 12310 26384 12316
rect 26240 11348 26292 11354
rect 26240 11290 26292 11296
rect 25964 10600 26016 10606
rect 25964 10542 26016 10548
rect 26240 10600 26292 10606
rect 26240 10542 26292 10548
rect 25976 10305 26004 10542
rect 25962 10296 26018 10305
rect 25962 10231 26018 10240
rect 25320 10124 25372 10130
rect 25320 10066 25372 10072
rect 25044 10056 25096 10062
rect 25044 9998 25096 10004
rect 25056 9926 25084 9998
rect 25044 9920 25096 9926
rect 25044 9862 25096 9868
rect 25056 8974 25084 9862
rect 25228 9512 25280 9518
rect 25228 9454 25280 9460
rect 25240 9178 25268 9454
rect 25228 9172 25280 9178
rect 25228 9114 25280 9120
rect 25044 8968 25096 8974
rect 25044 8910 25096 8916
rect 24964 6886 25084 6914
rect 24860 6860 24912 6866
rect 24860 6802 24912 6808
rect 24110 6012 24418 6032
rect 24110 6010 24116 6012
rect 24172 6010 24196 6012
rect 24252 6010 24276 6012
rect 24332 6010 24356 6012
rect 24412 6010 24418 6012
rect 24172 5958 24174 6010
rect 24354 5958 24356 6010
rect 24110 5956 24116 5958
rect 24172 5956 24196 5958
rect 24252 5956 24276 5958
rect 24332 5956 24356 5958
rect 24412 5956 24418 5958
rect 24110 5936 24418 5956
rect 22744 5704 22796 5710
rect 22744 5646 22796 5652
rect 22756 5234 22784 5646
rect 22744 5228 22796 5234
rect 22744 5170 22796 5176
rect 21364 4684 21416 4690
rect 21364 4626 21416 4632
rect 20720 4616 20772 4622
rect 20720 4558 20772 4564
rect 20628 4140 20680 4146
rect 20628 4082 20680 4088
rect 20640 3670 20668 4082
rect 20732 4078 20760 4558
rect 20904 4548 20956 4554
rect 20904 4490 20956 4496
rect 20916 4282 20944 4490
rect 20904 4276 20956 4282
rect 20904 4218 20956 4224
rect 20720 4072 20772 4078
rect 20720 4014 20772 4020
rect 20628 3664 20680 3670
rect 20628 3606 20680 3612
rect 21272 3528 21324 3534
rect 21272 3470 21324 3476
rect 21284 3058 21312 3470
rect 21272 3052 21324 3058
rect 21272 2994 21324 3000
rect 20444 2644 20496 2650
rect 20444 2586 20496 2592
rect 21376 2258 21404 4626
rect 22756 4146 22784 5170
rect 22836 5024 22888 5030
rect 22836 4966 22888 4972
rect 22744 4140 22796 4146
rect 22744 4082 22796 4088
rect 21916 3596 21968 3602
rect 21916 3538 21968 3544
rect 21284 2230 21404 2258
rect 21284 800 21312 2230
rect 21928 800 21956 3538
rect 22848 3058 22876 4966
rect 24110 4924 24418 4944
rect 24110 4922 24116 4924
rect 24172 4922 24196 4924
rect 24252 4922 24276 4924
rect 24332 4922 24356 4924
rect 24412 4922 24418 4924
rect 24172 4870 24174 4922
rect 24354 4870 24356 4922
rect 24110 4868 24116 4870
rect 24172 4868 24196 4870
rect 24252 4868 24276 4870
rect 24332 4868 24356 4870
rect 24412 4868 24418 4870
rect 24110 4848 24418 4868
rect 24110 3836 24418 3856
rect 24110 3834 24116 3836
rect 24172 3834 24196 3836
rect 24252 3834 24276 3836
rect 24332 3834 24356 3836
rect 24412 3834 24418 3836
rect 24172 3782 24174 3834
rect 24354 3782 24356 3834
rect 24110 3780 24116 3782
rect 24172 3780 24196 3782
rect 24252 3780 24276 3782
rect 24332 3780 24356 3782
rect 24412 3780 24418 3782
rect 24110 3760 24418 3780
rect 25056 3641 25084 6886
rect 25042 3632 25098 3641
rect 25042 3567 25098 3576
rect 24032 3528 24084 3534
rect 24032 3470 24084 3476
rect 24044 3058 24072 3470
rect 22836 3052 22888 3058
rect 22836 2994 22888 3000
rect 24032 3052 24084 3058
rect 24032 2994 24084 3000
rect 25136 2984 25188 2990
rect 25136 2926 25188 2932
rect 24110 2748 24418 2768
rect 24110 2746 24116 2748
rect 24172 2746 24196 2748
rect 24252 2746 24276 2748
rect 24332 2746 24356 2748
rect 24412 2746 24418 2748
rect 24172 2694 24174 2746
rect 24354 2694 24356 2746
rect 24110 2692 24116 2694
rect 24172 2692 24196 2694
rect 24252 2692 24276 2694
rect 24332 2692 24356 2694
rect 24412 2692 24418 2694
rect 24110 2672 24418 2692
rect 25148 800 25176 2926
rect 25332 2582 25360 10066
rect 26252 9722 26280 10542
rect 26240 9716 26292 9722
rect 26240 9658 26292 9664
rect 25504 9376 25556 9382
rect 25504 9318 25556 9324
rect 25516 7478 25544 9318
rect 26344 9042 26372 12310
rect 26436 12170 26464 14962
rect 26516 14816 26568 14822
rect 26516 14758 26568 14764
rect 26424 12164 26476 12170
rect 26424 12106 26476 12112
rect 26436 11898 26464 12106
rect 26424 11892 26476 11898
rect 26424 11834 26476 11840
rect 26528 9586 26556 14758
rect 26620 14278 26648 15846
rect 26608 14272 26660 14278
rect 26608 14214 26660 14220
rect 26516 9580 26568 9586
rect 26516 9522 26568 9528
rect 26332 9036 26384 9042
rect 26332 8978 26384 8984
rect 26146 8936 26202 8945
rect 26146 8871 26202 8880
rect 25964 8424 26016 8430
rect 25964 8366 26016 8372
rect 25976 8265 26004 8366
rect 25962 8256 26018 8265
rect 25962 8191 26018 8200
rect 25504 7472 25556 7478
rect 25504 7414 25556 7420
rect 26160 7342 26188 8871
rect 26240 8424 26292 8430
rect 26240 8366 26292 8372
rect 26424 8424 26476 8430
rect 26424 8366 26476 8372
rect 26252 8090 26280 8366
rect 26240 8084 26292 8090
rect 26240 8026 26292 8032
rect 26436 7410 26464 8366
rect 26424 7404 26476 7410
rect 26424 7346 26476 7352
rect 26148 7336 26200 7342
rect 26148 7278 26200 7284
rect 26332 6112 26384 6118
rect 26332 6054 26384 6060
rect 26344 5778 26372 6054
rect 26332 5772 26384 5778
rect 26332 5714 26384 5720
rect 26516 5636 26568 5642
rect 26516 5578 26568 5584
rect 26528 5370 26556 5578
rect 26516 5364 26568 5370
rect 26516 5306 26568 5312
rect 26804 4010 26832 22066
rect 27172 17270 27200 26846
rect 27528 25356 27580 25362
rect 27528 25298 27580 25304
rect 27540 25265 27568 25298
rect 27526 25256 27582 25265
rect 27526 25191 27582 25200
rect 27436 24608 27488 24614
rect 27436 24550 27488 24556
rect 27448 24138 27476 24550
rect 27528 24268 27580 24274
rect 27528 24210 27580 24216
rect 27436 24132 27488 24138
rect 27436 24074 27488 24080
rect 27448 23798 27476 24074
rect 27540 23905 27568 24210
rect 27526 23896 27582 23905
rect 27632 23866 27660 30194
rect 27988 28960 28040 28966
rect 27988 28902 28040 28908
rect 28000 28626 28028 28902
rect 27988 28620 28040 28626
rect 27988 28562 28040 28568
rect 28172 27872 28224 27878
rect 28172 27814 28224 27820
rect 28184 27538 28212 27814
rect 28172 27532 28224 27538
rect 28172 27474 28224 27480
rect 27712 27396 27764 27402
rect 27712 27338 27764 27344
rect 27724 27130 27752 27338
rect 27712 27124 27764 27130
rect 27712 27066 27764 27072
rect 27896 26988 27948 26994
rect 27896 26930 27948 26936
rect 27526 23831 27582 23840
rect 27620 23860 27672 23866
rect 27620 23802 27672 23808
rect 27436 23792 27488 23798
rect 27436 23734 27488 23740
rect 27344 23112 27396 23118
rect 27344 23054 27396 23060
rect 27356 20466 27384 23054
rect 27344 20460 27396 20466
rect 27344 20402 27396 20408
rect 27356 20369 27384 20402
rect 27342 20360 27398 20369
rect 27342 20295 27398 20304
rect 27342 19816 27398 19825
rect 27342 19751 27398 19760
rect 27356 18834 27384 19751
rect 27436 19168 27488 19174
rect 27436 19110 27488 19116
rect 27448 18834 27476 19110
rect 27344 18828 27396 18834
rect 27344 18770 27396 18776
rect 27436 18828 27488 18834
rect 27436 18770 27488 18776
rect 27632 18290 27660 23802
rect 27712 23248 27764 23254
rect 27712 23190 27764 23196
rect 27724 23050 27752 23190
rect 27712 23044 27764 23050
rect 27712 22986 27764 22992
rect 27724 22642 27752 22986
rect 27712 22636 27764 22642
rect 27712 22578 27764 22584
rect 27724 21554 27752 22578
rect 27712 21548 27764 21554
rect 27712 21490 27764 21496
rect 27804 18692 27856 18698
rect 27804 18634 27856 18640
rect 27816 18426 27844 18634
rect 27804 18420 27856 18426
rect 27804 18362 27856 18368
rect 27252 18284 27304 18290
rect 27252 18226 27304 18232
rect 27620 18284 27672 18290
rect 27620 18226 27672 18232
rect 27160 17264 27212 17270
rect 27160 17206 27212 17212
rect 27068 17196 27120 17202
rect 27068 17138 27120 17144
rect 26976 16788 27028 16794
rect 26976 16730 27028 16736
rect 26988 16046 27016 16730
rect 27080 16454 27108 17138
rect 27264 17082 27292 18226
rect 27528 17604 27580 17610
rect 27528 17546 27580 17552
rect 27436 17264 27488 17270
rect 27172 17054 27292 17082
rect 27356 17212 27436 17218
rect 27356 17206 27488 17212
rect 27356 17190 27476 17206
rect 27356 17066 27384 17190
rect 27344 17060 27396 17066
rect 27068 16448 27120 16454
rect 27068 16390 27120 16396
rect 26976 16040 27028 16046
rect 26976 15982 27028 15988
rect 26884 14884 26936 14890
rect 26884 14826 26936 14832
rect 26896 12714 26924 14826
rect 26988 13462 27016 15982
rect 26976 13456 27028 13462
rect 26976 13398 27028 13404
rect 26884 12708 26936 12714
rect 26884 12650 26936 12656
rect 26896 12238 26924 12650
rect 26976 12640 27028 12646
rect 26976 12582 27028 12588
rect 26884 12232 26936 12238
rect 26884 12174 26936 12180
rect 26988 10130 27016 12582
rect 26976 10124 27028 10130
rect 26976 10066 27028 10072
rect 27172 8498 27200 17054
rect 27344 17002 27396 17008
rect 27356 16250 27384 17002
rect 27344 16244 27396 16250
rect 27344 16186 27396 16192
rect 27252 14952 27304 14958
rect 27356 14940 27384 16186
rect 27304 14912 27384 14940
rect 27436 14952 27488 14958
rect 27252 14894 27304 14900
rect 27436 14894 27488 14900
rect 27264 14006 27292 14894
rect 27344 14816 27396 14822
rect 27344 14758 27396 14764
rect 27252 14000 27304 14006
rect 27252 13942 27304 13948
rect 27252 13864 27304 13870
rect 27252 13806 27304 13812
rect 27264 12238 27292 13806
rect 27356 12306 27384 14758
rect 27448 14618 27476 14894
rect 27540 14890 27568 17546
rect 27620 17196 27672 17202
rect 27620 17138 27672 17144
rect 27528 14884 27580 14890
rect 27528 14826 27580 14832
rect 27436 14612 27488 14618
rect 27436 14554 27488 14560
rect 27528 14476 27580 14482
rect 27528 14418 27580 14424
rect 27540 14385 27568 14418
rect 27526 14376 27582 14385
rect 27526 14311 27582 14320
rect 27528 13388 27580 13394
rect 27528 13330 27580 13336
rect 27540 12345 27568 13330
rect 27526 12336 27582 12345
rect 27344 12300 27396 12306
rect 27526 12271 27582 12280
rect 27344 12242 27396 12248
rect 27252 12232 27304 12238
rect 27252 12174 27304 12180
rect 27528 11212 27580 11218
rect 27528 11154 27580 11160
rect 27540 10985 27568 11154
rect 27526 10976 27582 10985
rect 27526 10911 27582 10920
rect 27632 10674 27660 17138
rect 27908 14498 27936 26930
rect 28172 26376 28224 26382
rect 28172 26318 28224 26324
rect 27988 25696 28040 25702
rect 27988 25638 28040 25644
rect 28000 25362 28028 25638
rect 28184 25362 28212 26318
rect 27988 25356 28040 25362
rect 27988 25298 28040 25304
rect 28172 25356 28224 25362
rect 28172 25298 28224 25304
rect 28264 24676 28316 24682
rect 28264 24618 28316 24624
rect 28172 24200 28224 24206
rect 28172 24142 28224 24148
rect 27988 24132 28040 24138
rect 27988 24074 28040 24080
rect 28000 23322 28028 24074
rect 27988 23316 28040 23322
rect 27988 23258 28040 23264
rect 28184 22094 28212 24142
rect 28092 22066 28212 22094
rect 28092 20466 28120 22066
rect 28170 21856 28226 21865
rect 28170 21791 28226 21800
rect 28184 21010 28212 21791
rect 28172 21004 28224 21010
rect 28172 20946 28224 20952
rect 28170 20496 28226 20505
rect 28080 20460 28132 20466
rect 28170 20431 28226 20440
rect 28080 20402 28132 20408
rect 28184 19922 28212 20431
rect 28172 19916 28224 19922
rect 28172 19858 28224 19864
rect 28172 19168 28224 19174
rect 28172 19110 28224 19116
rect 27988 16992 28040 16998
rect 27988 16934 28040 16940
rect 28000 16658 28028 16934
rect 28184 16658 28212 19110
rect 27988 16652 28040 16658
rect 27988 16594 28040 16600
rect 28172 16652 28224 16658
rect 28172 16594 28224 16600
rect 28078 16416 28134 16425
rect 28078 16351 28134 16360
rect 28092 16182 28120 16351
rect 28080 16176 28132 16182
rect 28080 16118 28132 16124
rect 27988 15904 28040 15910
rect 27988 15846 28040 15852
rect 28000 15706 28028 15846
rect 28170 15736 28226 15745
rect 27988 15700 28040 15706
rect 28170 15671 28226 15680
rect 27988 15642 28040 15648
rect 28184 15570 28212 15671
rect 28172 15564 28224 15570
rect 28172 15506 28224 15512
rect 27908 14470 28028 14498
rect 27896 14340 27948 14346
rect 27896 14282 27948 14288
rect 27908 14074 27936 14282
rect 27896 14068 27948 14074
rect 27896 14010 27948 14016
rect 27802 13968 27858 13977
rect 27802 13903 27804 13912
rect 27856 13903 27858 13912
rect 27804 13874 27856 13880
rect 27712 12844 27764 12850
rect 27712 12786 27764 12792
rect 27724 12442 27752 12786
rect 27712 12436 27764 12442
rect 27712 12378 27764 12384
rect 27712 12300 27764 12306
rect 27712 12242 27764 12248
rect 27620 10668 27672 10674
rect 27620 10610 27672 10616
rect 27528 9920 27580 9926
rect 27528 9862 27580 9868
rect 27540 9042 27568 9862
rect 27528 9036 27580 9042
rect 27528 8978 27580 8984
rect 27160 8492 27212 8498
rect 27160 8434 27212 8440
rect 27528 7948 27580 7954
rect 27528 7890 27580 7896
rect 27540 7585 27568 7890
rect 27526 7576 27582 7585
rect 27526 7511 27582 7520
rect 27526 6896 27582 6905
rect 27526 6831 27528 6840
rect 27580 6831 27582 6840
rect 27528 6802 27580 6808
rect 27632 6322 27660 10610
rect 27620 6316 27672 6322
rect 27620 6258 27672 6264
rect 27632 5846 27660 6258
rect 27620 5840 27672 5846
rect 27620 5782 27672 5788
rect 27436 4684 27488 4690
rect 27436 4626 27488 4632
rect 26792 4004 26844 4010
rect 26792 3946 26844 3952
rect 26424 3936 26476 3942
rect 26424 3878 26476 3884
rect 26976 3936 27028 3942
rect 26976 3878 27028 3884
rect 26240 2848 26292 2854
rect 25962 2816 26018 2825
rect 26240 2790 26292 2796
rect 25962 2751 26018 2760
rect 25320 2576 25372 2582
rect 25320 2518 25372 2524
rect 25976 2514 26004 2751
rect 26252 2514 26280 2790
rect 26436 2514 26464 3878
rect 26988 3602 27016 3878
rect 26976 3596 27028 3602
rect 26976 3538 27028 3544
rect 27448 3505 27476 4626
rect 27528 3596 27580 3602
rect 27528 3538 27580 3544
rect 27434 3496 27490 3505
rect 27068 3460 27120 3466
rect 27434 3431 27490 3440
rect 27068 3402 27120 3408
rect 26976 3392 27028 3398
rect 26976 3334 27028 3340
rect 26988 3058 27016 3334
rect 27080 3194 27108 3402
rect 27068 3188 27120 3194
rect 27068 3130 27120 3136
rect 26976 3052 27028 3058
rect 26976 2994 27028 3000
rect 25964 2508 26016 2514
rect 25964 2450 26016 2456
rect 26240 2508 26292 2514
rect 26240 2450 26292 2456
rect 26424 2508 26476 2514
rect 26424 2450 26476 2456
rect 27068 2440 27120 2446
rect 27068 2382 27120 2388
rect 27080 800 27108 2382
rect 27540 1465 27568 3538
rect 27724 3058 27752 12242
rect 27816 6848 27844 13874
rect 28000 12866 28028 14470
rect 28172 14408 28224 14414
rect 28172 14350 28224 14356
rect 28080 13252 28132 13258
rect 28080 13194 28132 13200
rect 28092 12986 28120 13194
rect 28080 12980 28132 12986
rect 28080 12922 28132 12928
rect 28000 12850 28120 12866
rect 27988 12844 28120 12850
rect 28040 12838 28120 12844
rect 27988 12786 28040 12792
rect 28000 12755 28028 12786
rect 27896 11552 27948 11558
rect 27896 11494 27948 11500
rect 27908 11218 27936 11494
rect 27896 11212 27948 11218
rect 27896 11154 27948 11160
rect 27988 11076 28040 11082
rect 27988 11018 28040 11024
rect 28000 10810 28028 11018
rect 27988 10804 28040 10810
rect 27988 10746 28040 10752
rect 27896 8356 27948 8362
rect 27896 8298 27948 8304
rect 27908 7818 27936 8298
rect 27988 8288 28040 8294
rect 27988 8230 28040 8236
rect 28000 7954 28028 8230
rect 27988 7948 28040 7954
rect 27988 7890 28040 7896
rect 27896 7812 27948 7818
rect 27896 7754 27948 7760
rect 27816 6820 27936 6848
rect 27804 6724 27856 6730
rect 27804 6666 27856 6672
rect 27816 6458 27844 6666
rect 27804 6452 27856 6458
rect 27804 6394 27856 6400
rect 27908 5234 27936 6820
rect 27896 5228 27948 5234
rect 27896 5170 27948 5176
rect 28092 3126 28120 12838
rect 28184 11762 28212 14350
rect 28172 11756 28224 11762
rect 28172 11698 28224 11704
rect 28276 9518 28304 24618
rect 28460 23254 28488 32370
rect 28630 32056 28686 32065
rect 28630 31991 28686 32000
rect 28540 30048 28592 30054
rect 28540 29990 28592 29996
rect 28448 23248 28500 23254
rect 28448 23190 28500 23196
rect 28356 23112 28408 23118
rect 28356 23054 28408 23060
rect 28368 10198 28396 23054
rect 28448 18284 28500 18290
rect 28448 18226 28500 18232
rect 28356 10192 28408 10198
rect 28356 10134 28408 10140
rect 28264 9512 28316 9518
rect 28264 9454 28316 9460
rect 28172 7200 28224 7206
rect 28172 7142 28224 7148
rect 28184 6866 28212 7142
rect 28172 6860 28224 6866
rect 28172 6802 28224 6808
rect 28172 5636 28224 5642
rect 28172 5578 28224 5584
rect 28184 5545 28212 5578
rect 28170 5536 28226 5545
rect 28170 5471 28226 5480
rect 28172 4616 28224 4622
rect 28172 4558 28224 4564
rect 28184 4146 28212 4558
rect 28172 4140 28224 4146
rect 28172 4082 28224 4088
rect 28460 3670 28488 18226
rect 28552 4690 28580 29990
rect 28644 22098 28672 31991
rect 28722 31376 28778 31385
rect 28722 31311 28778 31320
rect 28736 29714 28764 31311
rect 28724 29708 28776 29714
rect 28724 29650 28776 29656
rect 28632 22092 28684 22098
rect 28828 22094 28856 34954
rect 28632 22034 28684 22040
rect 28736 22066 28856 22094
rect 28736 18290 28764 22066
rect 28724 18284 28776 18290
rect 28724 18226 28776 18232
rect 29000 8900 29052 8906
rect 29000 8842 29052 8848
rect 28540 4684 28592 4690
rect 28540 4626 28592 4632
rect 28448 3664 28500 3670
rect 28448 3606 28500 3612
rect 28080 3120 28132 3126
rect 28080 3062 28132 3068
rect 27712 3052 27764 3058
rect 27712 2994 27764 3000
rect 29012 2145 29040 8842
rect 28998 2136 29054 2145
rect 28998 2071 29054 2080
rect 27526 1456 27582 1465
rect 27526 1391 27582 1400
rect -10 0 102 800
rect 634 0 746 800
rect 1278 0 1390 800
rect 1922 0 2034 800
rect 2566 0 2678 800
rect 3210 0 3322 800
rect 3854 0 3966 800
rect 4498 0 4610 800
rect 5786 0 5898 800
rect 6430 0 6542 800
rect 7074 0 7186 800
rect 7718 0 7830 800
rect 8362 0 8474 800
rect 9006 0 9118 800
rect 9650 0 9762 800
rect 10938 0 11050 800
rect 11582 0 11694 800
rect 12226 0 12338 800
rect 12870 0 12982 800
rect 13514 0 13626 800
rect 14158 0 14270 800
rect 14802 0 14914 800
rect 16090 0 16202 800
rect 16734 0 16846 800
rect 17378 0 17490 800
rect 18022 0 18134 800
rect 18666 0 18778 800
rect 19310 0 19422 800
rect 19954 0 20066 800
rect 21242 0 21354 800
rect 21886 0 21998 800
rect 22530 0 22642 800
rect 23174 0 23286 800
rect 23818 0 23930 800
rect 24462 0 24574 800
rect 25106 0 25218 800
rect 26394 0 26506 800
rect 27038 0 27150 800
rect 27682 0 27794 800
rect 28326 0 28438 800
rect 28970 0 29082 800
rect 29614 0 29726 800
<< via2 >>
rect 4066 49680 4122 49736
rect 1398 42200 1454 42256
rect 2870 44240 2926 44296
rect 5588 47354 5644 47356
rect 5668 47354 5724 47356
rect 5748 47354 5804 47356
rect 5828 47354 5884 47356
rect 5588 47302 5634 47354
rect 5634 47302 5644 47354
rect 5668 47302 5698 47354
rect 5698 47302 5710 47354
rect 5710 47302 5724 47354
rect 5748 47302 5762 47354
rect 5762 47302 5774 47354
rect 5774 47302 5804 47354
rect 5828 47302 5838 47354
rect 5838 47302 5884 47354
rect 5588 47300 5644 47302
rect 5668 47300 5724 47302
rect 5748 47300 5804 47302
rect 5828 47300 5884 47302
rect 5588 46266 5644 46268
rect 5668 46266 5724 46268
rect 5748 46266 5804 46268
rect 5828 46266 5884 46268
rect 5588 46214 5634 46266
rect 5634 46214 5644 46266
rect 5668 46214 5698 46266
rect 5698 46214 5710 46266
rect 5710 46214 5724 46266
rect 5748 46214 5762 46266
rect 5762 46214 5774 46266
rect 5774 46214 5804 46266
rect 5828 46214 5838 46266
rect 5838 46214 5884 46266
rect 5588 46212 5644 46214
rect 5668 46212 5724 46214
rect 5748 46212 5804 46214
rect 5828 46212 5884 46214
rect 3238 44920 3294 44976
rect 2778 41520 2834 41576
rect 2778 38800 2834 38856
rect 1398 37440 1454 37496
rect 1858 36780 1914 36816
rect 1858 36760 1860 36780
rect 1860 36760 1912 36780
rect 1912 36760 1914 36780
rect 1398 29960 1454 30016
rect 1398 27920 1454 27976
rect 1398 25200 1454 25256
rect 1766 34720 1822 34776
rect 1858 32000 1914 32056
rect 1858 19080 1914 19136
rect 2778 36080 2834 36136
rect 2778 25880 2834 25936
rect 3330 33360 3386 33416
rect 2962 19760 3018 19816
rect 2410 18400 2466 18456
rect 2778 17740 2834 17776
rect 2778 17720 2780 17740
rect 2780 17720 2832 17740
rect 2832 17720 2834 17740
rect 1858 14320 1914 14376
rect 1950 13640 2006 13696
rect 1950 11636 1952 11656
rect 1952 11636 2004 11656
rect 2004 11636 2006 11656
rect 1950 11600 2006 11636
rect 2778 15680 2834 15736
rect 1858 8880 1914 8936
rect 1398 4120 1454 4176
rect 3330 12280 3386 12336
rect 2870 7520 2926 7576
rect 2778 2760 2834 2816
rect 3422 8236 3424 8256
rect 3424 8236 3476 8256
rect 3476 8236 3478 8256
rect 3422 8200 3478 8236
rect 3422 6160 3478 6216
rect 3330 4800 3386 4856
rect 3974 15544 4030 15600
rect 5588 45178 5644 45180
rect 5668 45178 5724 45180
rect 5748 45178 5804 45180
rect 5828 45178 5884 45180
rect 5588 45126 5634 45178
rect 5634 45126 5644 45178
rect 5668 45126 5698 45178
rect 5698 45126 5710 45178
rect 5710 45126 5724 45178
rect 5748 45126 5762 45178
rect 5762 45126 5774 45178
rect 5774 45126 5804 45178
rect 5828 45126 5838 45178
rect 5838 45126 5884 45178
rect 5588 45124 5644 45126
rect 5668 45124 5724 45126
rect 5748 45124 5804 45126
rect 5828 45124 5884 45126
rect 5588 44090 5644 44092
rect 5668 44090 5724 44092
rect 5748 44090 5804 44092
rect 5828 44090 5884 44092
rect 5588 44038 5634 44090
rect 5634 44038 5644 44090
rect 5668 44038 5698 44090
rect 5698 44038 5710 44090
rect 5710 44038 5724 44090
rect 5748 44038 5762 44090
rect 5762 44038 5774 44090
rect 5774 44038 5804 44090
rect 5828 44038 5838 44090
rect 5838 44038 5884 44090
rect 5588 44036 5644 44038
rect 5668 44036 5724 44038
rect 5748 44036 5804 44038
rect 5828 44036 5884 44038
rect 5588 43002 5644 43004
rect 5668 43002 5724 43004
rect 5748 43002 5804 43004
rect 5828 43002 5884 43004
rect 5588 42950 5634 43002
rect 5634 42950 5644 43002
rect 5668 42950 5698 43002
rect 5698 42950 5710 43002
rect 5710 42950 5724 43002
rect 5748 42950 5762 43002
rect 5762 42950 5774 43002
rect 5774 42950 5804 43002
rect 5828 42950 5838 43002
rect 5838 42950 5884 43002
rect 5588 42948 5644 42950
rect 5668 42948 5724 42950
rect 5748 42948 5804 42950
rect 5828 42948 5884 42950
rect 5588 41914 5644 41916
rect 5668 41914 5724 41916
rect 5748 41914 5804 41916
rect 5828 41914 5884 41916
rect 5588 41862 5634 41914
rect 5634 41862 5644 41914
rect 5668 41862 5698 41914
rect 5698 41862 5710 41914
rect 5710 41862 5724 41914
rect 5748 41862 5762 41914
rect 5762 41862 5774 41914
rect 5774 41862 5804 41914
rect 5828 41862 5838 41914
rect 5838 41862 5884 41914
rect 5588 41860 5644 41862
rect 5668 41860 5724 41862
rect 5748 41860 5804 41862
rect 5828 41860 5884 41862
rect 5588 40826 5644 40828
rect 5668 40826 5724 40828
rect 5748 40826 5804 40828
rect 5828 40826 5884 40828
rect 5588 40774 5634 40826
rect 5634 40774 5644 40826
rect 5668 40774 5698 40826
rect 5698 40774 5710 40826
rect 5710 40774 5724 40826
rect 5748 40774 5762 40826
rect 5762 40774 5774 40826
rect 5774 40774 5804 40826
rect 5828 40774 5838 40826
rect 5838 40774 5884 40826
rect 5588 40772 5644 40774
rect 5668 40772 5724 40774
rect 5748 40772 5804 40774
rect 5828 40772 5884 40774
rect 5588 39738 5644 39740
rect 5668 39738 5724 39740
rect 5748 39738 5804 39740
rect 5828 39738 5884 39740
rect 5588 39686 5634 39738
rect 5634 39686 5644 39738
rect 5668 39686 5698 39738
rect 5698 39686 5710 39738
rect 5710 39686 5724 39738
rect 5748 39686 5762 39738
rect 5762 39686 5774 39738
rect 5774 39686 5804 39738
rect 5828 39686 5838 39738
rect 5838 39686 5884 39738
rect 5588 39684 5644 39686
rect 5668 39684 5724 39686
rect 5748 39684 5804 39686
rect 5828 39684 5884 39686
rect 5588 38650 5644 38652
rect 5668 38650 5724 38652
rect 5748 38650 5804 38652
rect 5828 38650 5884 38652
rect 5588 38598 5634 38650
rect 5634 38598 5644 38650
rect 5668 38598 5698 38650
rect 5698 38598 5710 38650
rect 5710 38598 5724 38650
rect 5748 38598 5762 38650
rect 5762 38598 5774 38650
rect 5774 38598 5804 38650
rect 5828 38598 5838 38650
rect 5838 38598 5884 38650
rect 5588 38596 5644 38598
rect 5668 38596 5724 38598
rect 5748 38596 5804 38598
rect 5828 38596 5884 38598
rect 5588 37562 5644 37564
rect 5668 37562 5724 37564
rect 5748 37562 5804 37564
rect 5828 37562 5884 37564
rect 5588 37510 5634 37562
rect 5634 37510 5644 37562
rect 5668 37510 5698 37562
rect 5698 37510 5710 37562
rect 5710 37510 5724 37562
rect 5748 37510 5762 37562
rect 5762 37510 5774 37562
rect 5774 37510 5804 37562
rect 5828 37510 5838 37562
rect 5838 37510 5884 37562
rect 5588 37508 5644 37510
rect 5668 37508 5724 37510
rect 5748 37508 5804 37510
rect 5828 37508 5884 37510
rect 5588 36474 5644 36476
rect 5668 36474 5724 36476
rect 5748 36474 5804 36476
rect 5828 36474 5884 36476
rect 5588 36422 5634 36474
rect 5634 36422 5644 36474
rect 5668 36422 5698 36474
rect 5698 36422 5710 36474
rect 5710 36422 5724 36474
rect 5748 36422 5762 36474
rect 5762 36422 5774 36474
rect 5774 36422 5804 36474
rect 5828 36422 5838 36474
rect 5838 36422 5884 36474
rect 5588 36420 5644 36422
rect 5668 36420 5724 36422
rect 5748 36420 5804 36422
rect 5828 36420 5884 36422
rect 5588 35386 5644 35388
rect 5668 35386 5724 35388
rect 5748 35386 5804 35388
rect 5828 35386 5884 35388
rect 5588 35334 5634 35386
rect 5634 35334 5644 35386
rect 5668 35334 5698 35386
rect 5698 35334 5710 35386
rect 5710 35334 5724 35386
rect 5748 35334 5762 35386
rect 5762 35334 5774 35386
rect 5774 35334 5804 35386
rect 5828 35334 5838 35386
rect 5838 35334 5884 35386
rect 5588 35332 5644 35334
rect 5668 35332 5724 35334
rect 5748 35332 5804 35334
rect 5828 35332 5884 35334
rect 5588 34298 5644 34300
rect 5668 34298 5724 34300
rect 5748 34298 5804 34300
rect 5828 34298 5884 34300
rect 5588 34246 5634 34298
rect 5634 34246 5644 34298
rect 5668 34246 5698 34298
rect 5698 34246 5710 34298
rect 5710 34246 5724 34298
rect 5748 34246 5762 34298
rect 5762 34246 5774 34298
rect 5774 34246 5804 34298
rect 5828 34246 5838 34298
rect 5838 34246 5884 34298
rect 5588 34244 5644 34246
rect 5668 34244 5724 34246
rect 5748 34244 5804 34246
rect 5828 34244 5884 34246
rect 5588 33210 5644 33212
rect 5668 33210 5724 33212
rect 5748 33210 5804 33212
rect 5828 33210 5884 33212
rect 5588 33158 5634 33210
rect 5634 33158 5644 33210
rect 5668 33158 5698 33210
rect 5698 33158 5710 33210
rect 5710 33158 5724 33210
rect 5748 33158 5762 33210
rect 5762 33158 5774 33210
rect 5774 33158 5804 33210
rect 5828 33158 5838 33210
rect 5838 33158 5884 33210
rect 5588 33156 5644 33158
rect 5668 33156 5724 33158
rect 5748 33156 5804 33158
rect 5828 33156 5884 33158
rect 5588 32122 5644 32124
rect 5668 32122 5724 32124
rect 5748 32122 5804 32124
rect 5828 32122 5884 32124
rect 5588 32070 5634 32122
rect 5634 32070 5644 32122
rect 5668 32070 5698 32122
rect 5698 32070 5710 32122
rect 5710 32070 5724 32122
rect 5748 32070 5762 32122
rect 5762 32070 5774 32122
rect 5774 32070 5804 32122
rect 5828 32070 5838 32122
rect 5838 32070 5884 32122
rect 5588 32068 5644 32070
rect 5668 32068 5724 32070
rect 5748 32068 5804 32070
rect 5828 32068 5884 32070
rect 5588 31034 5644 31036
rect 5668 31034 5724 31036
rect 5748 31034 5804 31036
rect 5828 31034 5884 31036
rect 5588 30982 5634 31034
rect 5634 30982 5644 31034
rect 5668 30982 5698 31034
rect 5698 30982 5710 31034
rect 5710 30982 5724 31034
rect 5748 30982 5762 31034
rect 5762 30982 5774 31034
rect 5774 30982 5804 31034
rect 5828 30982 5838 31034
rect 5838 30982 5884 31034
rect 5588 30980 5644 30982
rect 5668 30980 5724 30982
rect 5748 30980 5804 30982
rect 5828 30980 5884 30982
rect 5588 29946 5644 29948
rect 5668 29946 5724 29948
rect 5748 29946 5804 29948
rect 5828 29946 5884 29948
rect 5588 29894 5634 29946
rect 5634 29894 5644 29946
rect 5668 29894 5698 29946
rect 5698 29894 5710 29946
rect 5710 29894 5724 29946
rect 5748 29894 5762 29946
rect 5762 29894 5774 29946
rect 5774 29894 5804 29946
rect 5828 29894 5838 29946
rect 5838 29894 5884 29946
rect 5588 29892 5644 29894
rect 5668 29892 5724 29894
rect 5748 29892 5804 29894
rect 5828 29892 5884 29894
rect 5588 28858 5644 28860
rect 5668 28858 5724 28860
rect 5748 28858 5804 28860
rect 5828 28858 5884 28860
rect 5588 28806 5634 28858
rect 5634 28806 5644 28858
rect 5668 28806 5698 28858
rect 5698 28806 5710 28858
rect 5710 28806 5724 28858
rect 5748 28806 5762 28858
rect 5762 28806 5774 28858
rect 5774 28806 5804 28858
rect 5828 28806 5838 28858
rect 5838 28806 5884 28858
rect 5588 28804 5644 28806
rect 5668 28804 5724 28806
rect 5748 28804 5804 28806
rect 5828 28804 5884 28806
rect 5588 27770 5644 27772
rect 5668 27770 5724 27772
rect 5748 27770 5804 27772
rect 5828 27770 5884 27772
rect 5588 27718 5634 27770
rect 5634 27718 5644 27770
rect 5668 27718 5698 27770
rect 5698 27718 5710 27770
rect 5710 27718 5724 27770
rect 5748 27718 5762 27770
rect 5762 27718 5774 27770
rect 5774 27718 5804 27770
rect 5828 27718 5838 27770
rect 5838 27718 5884 27770
rect 5588 27716 5644 27718
rect 5668 27716 5724 27718
rect 5748 27716 5804 27718
rect 5828 27716 5884 27718
rect 5588 26682 5644 26684
rect 5668 26682 5724 26684
rect 5748 26682 5804 26684
rect 5828 26682 5884 26684
rect 5588 26630 5634 26682
rect 5634 26630 5644 26682
rect 5668 26630 5698 26682
rect 5698 26630 5710 26682
rect 5710 26630 5724 26682
rect 5748 26630 5762 26682
rect 5762 26630 5774 26682
rect 5774 26630 5804 26682
rect 5828 26630 5838 26682
rect 5838 26630 5884 26682
rect 5588 26628 5644 26630
rect 5668 26628 5724 26630
rect 5748 26628 5804 26630
rect 5828 26628 5884 26630
rect 5588 25594 5644 25596
rect 5668 25594 5724 25596
rect 5748 25594 5804 25596
rect 5828 25594 5884 25596
rect 5588 25542 5634 25594
rect 5634 25542 5644 25594
rect 5668 25542 5698 25594
rect 5698 25542 5710 25594
rect 5710 25542 5724 25594
rect 5748 25542 5762 25594
rect 5762 25542 5774 25594
rect 5774 25542 5804 25594
rect 5828 25542 5838 25594
rect 5838 25542 5884 25594
rect 5588 25540 5644 25542
rect 5668 25540 5724 25542
rect 5748 25540 5804 25542
rect 5828 25540 5884 25542
rect 5588 24506 5644 24508
rect 5668 24506 5724 24508
rect 5748 24506 5804 24508
rect 5828 24506 5884 24508
rect 5588 24454 5634 24506
rect 5634 24454 5644 24506
rect 5668 24454 5698 24506
rect 5698 24454 5710 24506
rect 5710 24454 5724 24506
rect 5748 24454 5762 24506
rect 5762 24454 5774 24506
rect 5774 24454 5804 24506
rect 5828 24454 5838 24506
rect 5838 24454 5884 24506
rect 5588 24452 5644 24454
rect 5668 24452 5724 24454
rect 5748 24452 5804 24454
rect 5828 24452 5884 24454
rect 3698 3440 3754 3496
rect 5262 3984 5318 4040
rect 5588 23418 5644 23420
rect 5668 23418 5724 23420
rect 5748 23418 5804 23420
rect 5828 23418 5884 23420
rect 5588 23366 5634 23418
rect 5634 23366 5644 23418
rect 5668 23366 5698 23418
rect 5698 23366 5710 23418
rect 5710 23366 5724 23418
rect 5748 23366 5762 23418
rect 5762 23366 5774 23418
rect 5774 23366 5804 23418
rect 5828 23366 5838 23418
rect 5838 23366 5884 23418
rect 5588 23364 5644 23366
rect 5668 23364 5724 23366
rect 5748 23364 5804 23366
rect 5828 23364 5884 23366
rect 5588 22330 5644 22332
rect 5668 22330 5724 22332
rect 5748 22330 5804 22332
rect 5828 22330 5884 22332
rect 5588 22278 5634 22330
rect 5634 22278 5644 22330
rect 5668 22278 5698 22330
rect 5698 22278 5710 22330
rect 5710 22278 5724 22330
rect 5748 22278 5762 22330
rect 5762 22278 5774 22330
rect 5774 22278 5804 22330
rect 5828 22278 5838 22330
rect 5838 22278 5884 22330
rect 5588 22276 5644 22278
rect 5668 22276 5724 22278
rect 5748 22276 5804 22278
rect 5828 22276 5884 22278
rect 5588 21242 5644 21244
rect 5668 21242 5724 21244
rect 5748 21242 5804 21244
rect 5828 21242 5884 21244
rect 5588 21190 5634 21242
rect 5634 21190 5644 21242
rect 5668 21190 5698 21242
rect 5698 21190 5710 21242
rect 5710 21190 5724 21242
rect 5748 21190 5762 21242
rect 5762 21190 5774 21242
rect 5774 21190 5804 21242
rect 5828 21190 5838 21242
rect 5838 21190 5884 21242
rect 5588 21188 5644 21190
rect 5668 21188 5724 21190
rect 5748 21188 5804 21190
rect 5828 21188 5884 21190
rect 5588 20154 5644 20156
rect 5668 20154 5724 20156
rect 5748 20154 5804 20156
rect 5828 20154 5884 20156
rect 5588 20102 5634 20154
rect 5634 20102 5644 20154
rect 5668 20102 5698 20154
rect 5698 20102 5710 20154
rect 5710 20102 5724 20154
rect 5748 20102 5762 20154
rect 5762 20102 5774 20154
rect 5774 20102 5804 20154
rect 5828 20102 5838 20154
rect 5838 20102 5884 20154
rect 5588 20100 5644 20102
rect 5668 20100 5724 20102
rect 5748 20100 5804 20102
rect 5828 20100 5884 20102
rect 5588 19066 5644 19068
rect 5668 19066 5724 19068
rect 5748 19066 5804 19068
rect 5828 19066 5884 19068
rect 5588 19014 5634 19066
rect 5634 19014 5644 19066
rect 5668 19014 5698 19066
rect 5698 19014 5710 19066
rect 5710 19014 5724 19066
rect 5748 19014 5762 19066
rect 5762 19014 5774 19066
rect 5774 19014 5804 19066
rect 5828 19014 5838 19066
rect 5838 19014 5884 19066
rect 5588 19012 5644 19014
rect 5668 19012 5724 19014
rect 5748 19012 5804 19014
rect 5828 19012 5884 19014
rect 5588 17978 5644 17980
rect 5668 17978 5724 17980
rect 5748 17978 5804 17980
rect 5828 17978 5884 17980
rect 5588 17926 5634 17978
rect 5634 17926 5644 17978
rect 5668 17926 5698 17978
rect 5698 17926 5710 17978
rect 5710 17926 5724 17978
rect 5748 17926 5762 17978
rect 5762 17926 5774 17978
rect 5774 17926 5804 17978
rect 5828 17926 5838 17978
rect 5838 17926 5884 17978
rect 5588 17924 5644 17926
rect 5668 17924 5724 17926
rect 5748 17924 5804 17926
rect 5828 17924 5884 17926
rect 5588 16890 5644 16892
rect 5668 16890 5724 16892
rect 5748 16890 5804 16892
rect 5828 16890 5884 16892
rect 5588 16838 5634 16890
rect 5634 16838 5644 16890
rect 5668 16838 5698 16890
rect 5698 16838 5710 16890
rect 5710 16838 5724 16890
rect 5748 16838 5762 16890
rect 5762 16838 5774 16890
rect 5774 16838 5804 16890
rect 5828 16838 5838 16890
rect 5838 16838 5884 16890
rect 5588 16836 5644 16838
rect 5668 16836 5724 16838
rect 5748 16836 5804 16838
rect 5828 16836 5884 16838
rect 10220 46810 10276 46812
rect 10300 46810 10356 46812
rect 10380 46810 10436 46812
rect 10460 46810 10516 46812
rect 10220 46758 10266 46810
rect 10266 46758 10276 46810
rect 10300 46758 10330 46810
rect 10330 46758 10342 46810
rect 10342 46758 10356 46810
rect 10380 46758 10394 46810
rect 10394 46758 10406 46810
rect 10406 46758 10436 46810
rect 10460 46758 10470 46810
rect 10470 46758 10516 46810
rect 10220 46756 10276 46758
rect 10300 46756 10356 46758
rect 10380 46756 10436 46758
rect 10460 46756 10516 46758
rect 10220 45722 10276 45724
rect 10300 45722 10356 45724
rect 10380 45722 10436 45724
rect 10460 45722 10516 45724
rect 10220 45670 10266 45722
rect 10266 45670 10276 45722
rect 10300 45670 10330 45722
rect 10330 45670 10342 45722
rect 10342 45670 10356 45722
rect 10380 45670 10394 45722
rect 10394 45670 10406 45722
rect 10406 45670 10436 45722
rect 10460 45670 10470 45722
rect 10470 45670 10516 45722
rect 10220 45668 10276 45670
rect 10300 45668 10356 45670
rect 10380 45668 10436 45670
rect 10460 45668 10516 45670
rect 14852 47354 14908 47356
rect 14932 47354 14988 47356
rect 15012 47354 15068 47356
rect 15092 47354 15148 47356
rect 14852 47302 14898 47354
rect 14898 47302 14908 47354
rect 14932 47302 14962 47354
rect 14962 47302 14974 47354
rect 14974 47302 14988 47354
rect 15012 47302 15026 47354
rect 15026 47302 15038 47354
rect 15038 47302 15068 47354
rect 15092 47302 15102 47354
rect 15102 47302 15148 47354
rect 14852 47300 14908 47302
rect 14932 47300 14988 47302
rect 15012 47300 15068 47302
rect 15092 47300 15148 47302
rect 14852 46266 14908 46268
rect 14932 46266 14988 46268
rect 15012 46266 15068 46268
rect 15092 46266 15148 46268
rect 14852 46214 14898 46266
rect 14898 46214 14908 46266
rect 14932 46214 14962 46266
rect 14962 46214 14974 46266
rect 14974 46214 14988 46266
rect 15012 46214 15026 46266
rect 15026 46214 15038 46266
rect 15038 46214 15068 46266
rect 15092 46214 15102 46266
rect 15102 46214 15148 46266
rect 14852 46212 14908 46214
rect 14932 46212 14988 46214
rect 15012 46212 15068 46214
rect 15092 46212 15148 46214
rect 14852 45178 14908 45180
rect 14932 45178 14988 45180
rect 15012 45178 15068 45180
rect 15092 45178 15148 45180
rect 14852 45126 14898 45178
rect 14898 45126 14908 45178
rect 14932 45126 14962 45178
rect 14962 45126 14974 45178
rect 14974 45126 14988 45178
rect 15012 45126 15026 45178
rect 15026 45126 15038 45178
rect 15038 45126 15068 45178
rect 15092 45126 15102 45178
rect 15102 45126 15148 45178
rect 14852 45124 14908 45126
rect 14932 45124 14988 45126
rect 15012 45124 15068 45126
rect 15092 45124 15148 45126
rect 10220 44634 10276 44636
rect 10300 44634 10356 44636
rect 10380 44634 10436 44636
rect 10460 44634 10516 44636
rect 10220 44582 10266 44634
rect 10266 44582 10276 44634
rect 10300 44582 10330 44634
rect 10330 44582 10342 44634
rect 10342 44582 10356 44634
rect 10380 44582 10394 44634
rect 10394 44582 10406 44634
rect 10406 44582 10436 44634
rect 10460 44582 10470 44634
rect 10470 44582 10516 44634
rect 10220 44580 10276 44582
rect 10300 44580 10356 44582
rect 10380 44580 10436 44582
rect 10460 44580 10516 44582
rect 10220 43546 10276 43548
rect 10300 43546 10356 43548
rect 10380 43546 10436 43548
rect 10460 43546 10516 43548
rect 10220 43494 10266 43546
rect 10266 43494 10276 43546
rect 10300 43494 10330 43546
rect 10330 43494 10342 43546
rect 10342 43494 10356 43546
rect 10380 43494 10394 43546
rect 10394 43494 10406 43546
rect 10406 43494 10436 43546
rect 10460 43494 10470 43546
rect 10470 43494 10516 43546
rect 10220 43492 10276 43494
rect 10300 43492 10356 43494
rect 10380 43492 10436 43494
rect 10460 43492 10516 43494
rect 10220 42458 10276 42460
rect 10300 42458 10356 42460
rect 10380 42458 10436 42460
rect 10460 42458 10516 42460
rect 10220 42406 10266 42458
rect 10266 42406 10276 42458
rect 10300 42406 10330 42458
rect 10330 42406 10342 42458
rect 10342 42406 10356 42458
rect 10380 42406 10394 42458
rect 10394 42406 10406 42458
rect 10406 42406 10436 42458
rect 10460 42406 10470 42458
rect 10470 42406 10516 42458
rect 10220 42404 10276 42406
rect 10300 42404 10356 42406
rect 10380 42404 10436 42406
rect 10460 42404 10516 42406
rect 10220 41370 10276 41372
rect 10300 41370 10356 41372
rect 10380 41370 10436 41372
rect 10460 41370 10516 41372
rect 10220 41318 10266 41370
rect 10266 41318 10276 41370
rect 10300 41318 10330 41370
rect 10330 41318 10342 41370
rect 10342 41318 10356 41370
rect 10380 41318 10394 41370
rect 10394 41318 10406 41370
rect 10406 41318 10436 41370
rect 10460 41318 10470 41370
rect 10470 41318 10516 41370
rect 10220 41316 10276 41318
rect 10300 41316 10356 41318
rect 10380 41316 10436 41318
rect 10460 41316 10516 41318
rect 10220 40282 10276 40284
rect 10300 40282 10356 40284
rect 10380 40282 10436 40284
rect 10460 40282 10516 40284
rect 10220 40230 10266 40282
rect 10266 40230 10276 40282
rect 10300 40230 10330 40282
rect 10330 40230 10342 40282
rect 10342 40230 10356 40282
rect 10380 40230 10394 40282
rect 10394 40230 10406 40282
rect 10406 40230 10436 40282
rect 10460 40230 10470 40282
rect 10470 40230 10516 40282
rect 10220 40228 10276 40230
rect 10300 40228 10356 40230
rect 10380 40228 10436 40230
rect 10460 40228 10516 40230
rect 10220 39194 10276 39196
rect 10300 39194 10356 39196
rect 10380 39194 10436 39196
rect 10460 39194 10516 39196
rect 10220 39142 10266 39194
rect 10266 39142 10276 39194
rect 10300 39142 10330 39194
rect 10330 39142 10342 39194
rect 10342 39142 10356 39194
rect 10380 39142 10394 39194
rect 10394 39142 10406 39194
rect 10406 39142 10436 39194
rect 10460 39142 10470 39194
rect 10470 39142 10516 39194
rect 10220 39140 10276 39142
rect 10300 39140 10356 39142
rect 10380 39140 10436 39142
rect 10460 39140 10516 39142
rect 10220 38106 10276 38108
rect 10300 38106 10356 38108
rect 10380 38106 10436 38108
rect 10460 38106 10516 38108
rect 10220 38054 10266 38106
rect 10266 38054 10276 38106
rect 10300 38054 10330 38106
rect 10330 38054 10342 38106
rect 10342 38054 10356 38106
rect 10380 38054 10394 38106
rect 10394 38054 10406 38106
rect 10406 38054 10436 38106
rect 10460 38054 10470 38106
rect 10470 38054 10516 38106
rect 10220 38052 10276 38054
rect 10300 38052 10356 38054
rect 10380 38052 10436 38054
rect 10460 38052 10516 38054
rect 10220 37018 10276 37020
rect 10300 37018 10356 37020
rect 10380 37018 10436 37020
rect 10460 37018 10516 37020
rect 10220 36966 10266 37018
rect 10266 36966 10276 37018
rect 10300 36966 10330 37018
rect 10330 36966 10342 37018
rect 10342 36966 10356 37018
rect 10380 36966 10394 37018
rect 10394 36966 10406 37018
rect 10406 36966 10436 37018
rect 10460 36966 10470 37018
rect 10470 36966 10516 37018
rect 10220 36964 10276 36966
rect 10300 36964 10356 36966
rect 10380 36964 10436 36966
rect 10460 36964 10516 36966
rect 10220 35930 10276 35932
rect 10300 35930 10356 35932
rect 10380 35930 10436 35932
rect 10460 35930 10516 35932
rect 10220 35878 10266 35930
rect 10266 35878 10276 35930
rect 10300 35878 10330 35930
rect 10330 35878 10342 35930
rect 10342 35878 10356 35930
rect 10380 35878 10394 35930
rect 10394 35878 10406 35930
rect 10406 35878 10436 35930
rect 10460 35878 10470 35930
rect 10470 35878 10516 35930
rect 10220 35876 10276 35878
rect 10300 35876 10356 35878
rect 10380 35876 10436 35878
rect 10460 35876 10516 35878
rect 14852 44090 14908 44092
rect 14932 44090 14988 44092
rect 15012 44090 15068 44092
rect 15092 44090 15148 44092
rect 14852 44038 14898 44090
rect 14898 44038 14908 44090
rect 14932 44038 14962 44090
rect 14962 44038 14974 44090
rect 14974 44038 14988 44090
rect 15012 44038 15026 44090
rect 15026 44038 15038 44090
rect 15038 44038 15068 44090
rect 15092 44038 15102 44090
rect 15102 44038 15148 44090
rect 14852 44036 14908 44038
rect 14932 44036 14988 44038
rect 15012 44036 15068 44038
rect 15092 44036 15148 44038
rect 14852 43002 14908 43004
rect 14932 43002 14988 43004
rect 15012 43002 15068 43004
rect 15092 43002 15148 43004
rect 14852 42950 14898 43002
rect 14898 42950 14908 43002
rect 14932 42950 14962 43002
rect 14962 42950 14974 43002
rect 14974 42950 14988 43002
rect 15012 42950 15026 43002
rect 15026 42950 15038 43002
rect 15038 42950 15068 43002
rect 15092 42950 15102 43002
rect 15102 42950 15148 43002
rect 14852 42948 14908 42950
rect 14932 42948 14988 42950
rect 15012 42948 15068 42950
rect 15092 42948 15148 42950
rect 14852 41914 14908 41916
rect 14932 41914 14988 41916
rect 15012 41914 15068 41916
rect 15092 41914 15148 41916
rect 14852 41862 14898 41914
rect 14898 41862 14908 41914
rect 14932 41862 14962 41914
rect 14962 41862 14974 41914
rect 14974 41862 14988 41914
rect 15012 41862 15026 41914
rect 15026 41862 15038 41914
rect 15038 41862 15068 41914
rect 15092 41862 15102 41914
rect 15102 41862 15148 41914
rect 14852 41860 14908 41862
rect 14932 41860 14988 41862
rect 15012 41860 15068 41862
rect 15092 41860 15148 41862
rect 14852 40826 14908 40828
rect 14932 40826 14988 40828
rect 15012 40826 15068 40828
rect 15092 40826 15148 40828
rect 14852 40774 14898 40826
rect 14898 40774 14908 40826
rect 14932 40774 14962 40826
rect 14962 40774 14974 40826
rect 14974 40774 14988 40826
rect 15012 40774 15026 40826
rect 15026 40774 15038 40826
rect 15038 40774 15068 40826
rect 15092 40774 15102 40826
rect 15102 40774 15148 40826
rect 14852 40772 14908 40774
rect 14932 40772 14988 40774
rect 15012 40772 15068 40774
rect 15092 40772 15148 40774
rect 14852 39738 14908 39740
rect 14932 39738 14988 39740
rect 15012 39738 15068 39740
rect 15092 39738 15148 39740
rect 14852 39686 14898 39738
rect 14898 39686 14908 39738
rect 14932 39686 14962 39738
rect 14962 39686 14974 39738
rect 14974 39686 14988 39738
rect 15012 39686 15026 39738
rect 15026 39686 15038 39738
rect 15038 39686 15068 39738
rect 15092 39686 15102 39738
rect 15102 39686 15148 39738
rect 14852 39684 14908 39686
rect 14932 39684 14988 39686
rect 15012 39684 15068 39686
rect 15092 39684 15148 39686
rect 14852 38650 14908 38652
rect 14932 38650 14988 38652
rect 15012 38650 15068 38652
rect 15092 38650 15148 38652
rect 14852 38598 14898 38650
rect 14898 38598 14908 38650
rect 14932 38598 14962 38650
rect 14962 38598 14974 38650
rect 14974 38598 14988 38650
rect 15012 38598 15026 38650
rect 15026 38598 15038 38650
rect 15038 38598 15068 38650
rect 15092 38598 15102 38650
rect 15102 38598 15148 38650
rect 14852 38596 14908 38598
rect 14932 38596 14988 38598
rect 15012 38596 15068 38598
rect 15092 38596 15148 38598
rect 14852 37562 14908 37564
rect 14932 37562 14988 37564
rect 15012 37562 15068 37564
rect 15092 37562 15148 37564
rect 14852 37510 14898 37562
rect 14898 37510 14908 37562
rect 14932 37510 14962 37562
rect 14962 37510 14974 37562
rect 14974 37510 14988 37562
rect 15012 37510 15026 37562
rect 15026 37510 15038 37562
rect 15038 37510 15068 37562
rect 15092 37510 15102 37562
rect 15102 37510 15148 37562
rect 14852 37508 14908 37510
rect 14932 37508 14988 37510
rect 15012 37508 15068 37510
rect 15092 37508 15148 37510
rect 14852 36474 14908 36476
rect 14932 36474 14988 36476
rect 15012 36474 15068 36476
rect 15092 36474 15148 36476
rect 14852 36422 14898 36474
rect 14898 36422 14908 36474
rect 14932 36422 14962 36474
rect 14962 36422 14974 36474
rect 14974 36422 14988 36474
rect 15012 36422 15026 36474
rect 15026 36422 15038 36474
rect 15038 36422 15068 36474
rect 15092 36422 15102 36474
rect 15102 36422 15148 36474
rect 14852 36420 14908 36422
rect 14932 36420 14988 36422
rect 15012 36420 15068 36422
rect 15092 36420 15148 36422
rect 14852 35386 14908 35388
rect 14932 35386 14988 35388
rect 15012 35386 15068 35388
rect 15092 35386 15148 35388
rect 14852 35334 14898 35386
rect 14898 35334 14908 35386
rect 14932 35334 14962 35386
rect 14962 35334 14974 35386
rect 14974 35334 14988 35386
rect 15012 35334 15026 35386
rect 15026 35334 15038 35386
rect 15038 35334 15068 35386
rect 15092 35334 15102 35386
rect 15102 35334 15148 35386
rect 14852 35332 14908 35334
rect 14932 35332 14988 35334
rect 15012 35332 15068 35334
rect 15092 35332 15148 35334
rect 10598 35128 10654 35184
rect 10220 34842 10276 34844
rect 10300 34842 10356 34844
rect 10380 34842 10436 34844
rect 10460 34842 10516 34844
rect 10220 34790 10266 34842
rect 10266 34790 10276 34842
rect 10300 34790 10330 34842
rect 10330 34790 10342 34842
rect 10342 34790 10356 34842
rect 10380 34790 10394 34842
rect 10394 34790 10406 34842
rect 10406 34790 10436 34842
rect 10460 34790 10470 34842
rect 10470 34790 10516 34842
rect 10220 34788 10276 34790
rect 10300 34788 10356 34790
rect 10380 34788 10436 34790
rect 10460 34788 10516 34790
rect 14852 34298 14908 34300
rect 14932 34298 14988 34300
rect 15012 34298 15068 34300
rect 15092 34298 15148 34300
rect 14852 34246 14898 34298
rect 14898 34246 14908 34298
rect 14932 34246 14962 34298
rect 14962 34246 14974 34298
rect 14974 34246 14988 34298
rect 15012 34246 15026 34298
rect 15026 34246 15038 34298
rect 15038 34246 15068 34298
rect 15092 34246 15102 34298
rect 15102 34246 15148 34298
rect 14852 34244 14908 34246
rect 14932 34244 14988 34246
rect 15012 34244 15068 34246
rect 15092 34244 15148 34246
rect 10220 33754 10276 33756
rect 10300 33754 10356 33756
rect 10380 33754 10436 33756
rect 10460 33754 10516 33756
rect 10220 33702 10266 33754
rect 10266 33702 10276 33754
rect 10300 33702 10330 33754
rect 10330 33702 10342 33754
rect 10342 33702 10356 33754
rect 10380 33702 10394 33754
rect 10394 33702 10406 33754
rect 10406 33702 10436 33754
rect 10460 33702 10470 33754
rect 10470 33702 10516 33754
rect 10220 33700 10276 33702
rect 10300 33700 10356 33702
rect 10380 33700 10436 33702
rect 10460 33700 10516 33702
rect 14852 33210 14908 33212
rect 14932 33210 14988 33212
rect 15012 33210 15068 33212
rect 15092 33210 15148 33212
rect 14852 33158 14898 33210
rect 14898 33158 14908 33210
rect 14932 33158 14962 33210
rect 14962 33158 14974 33210
rect 14974 33158 14988 33210
rect 15012 33158 15026 33210
rect 15026 33158 15038 33210
rect 15038 33158 15068 33210
rect 15092 33158 15102 33210
rect 15102 33158 15148 33210
rect 14852 33156 14908 33158
rect 14932 33156 14988 33158
rect 15012 33156 15068 33158
rect 15092 33156 15148 33158
rect 10220 32666 10276 32668
rect 10300 32666 10356 32668
rect 10380 32666 10436 32668
rect 10460 32666 10516 32668
rect 10220 32614 10266 32666
rect 10266 32614 10276 32666
rect 10300 32614 10330 32666
rect 10330 32614 10342 32666
rect 10342 32614 10356 32666
rect 10380 32614 10394 32666
rect 10394 32614 10406 32666
rect 10406 32614 10436 32666
rect 10460 32614 10470 32666
rect 10470 32614 10516 32666
rect 10220 32612 10276 32614
rect 10300 32612 10356 32614
rect 10380 32612 10436 32614
rect 10460 32612 10516 32614
rect 14852 32122 14908 32124
rect 14932 32122 14988 32124
rect 15012 32122 15068 32124
rect 15092 32122 15148 32124
rect 14852 32070 14898 32122
rect 14898 32070 14908 32122
rect 14932 32070 14962 32122
rect 14962 32070 14974 32122
rect 14974 32070 14988 32122
rect 15012 32070 15026 32122
rect 15026 32070 15038 32122
rect 15038 32070 15068 32122
rect 15092 32070 15102 32122
rect 15102 32070 15148 32122
rect 14852 32068 14908 32070
rect 14932 32068 14988 32070
rect 15012 32068 15068 32070
rect 15092 32068 15148 32070
rect 19484 46810 19540 46812
rect 19564 46810 19620 46812
rect 19644 46810 19700 46812
rect 19724 46810 19780 46812
rect 19484 46758 19530 46810
rect 19530 46758 19540 46810
rect 19564 46758 19594 46810
rect 19594 46758 19606 46810
rect 19606 46758 19620 46810
rect 19644 46758 19658 46810
rect 19658 46758 19670 46810
rect 19670 46758 19700 46810
rect 19724 46758 19734 46810
rect 19734 46758 19780 46810
rect 19484 46756 19540 46758
rect 19564 46756 19620 46758
rect 19644 46756 19700 46758
rect 19724 46756 19780 46758
rect 19484 45722 19540 45724
rect 19564 45722 19620 45724
rect 19644 45722 19700 45724
rect 19724 45722 19780 45724
rect 19484 45670 19530 45722
rect 19530 45670 19540 45722
rect 19564 45670 19594 45722
rect 19594 45670 19606 45722
rect 19606 45670 19620 45722
rect 19644 45670 19658 45722
rect 19658 45670 19670 45722
rect 19670 45670 19700 45722
rect 19724 45670 19734 45722
rect 19734 45670 19780 45722
rect 19484 45668 19540 45670
rect 19564 45668 19620 45670
rect 19644 45668 19700 45670
rect 19724 45668 19780 45670
rect 19484 44634 19540 44636
rect 19564 44634 19620 44636
rect 19644 44634 19700 44636
rect 19724 44634 19780 44636
rect 19484 44582 19530 44634
rect 19530 44582 19540 44634
rect 19564 44582 19594 44634
rect 19594 44582 19606 44634
rect 19606 44582 19620 44634
rect 19644 44582 19658 44634
rect 19658 44582 19670 44634
rect 19670 44582 19700 44634
rect 19724 44582 19734 44634
rect 19734 44582 19780 44634
rect 19484 44580 19540 44582
rect 19564 44580 19620 44582
rect 19644 44580 19700 44582
rect 19724 44580 19780 44582
rect 19484 43546 19540 43548
rect 19564 43546 19620 43548
rect 19644 43546 19700 43548
rect 19724 43546 19780 43548
rect 19484 43494 19530 43546
rect 19530 43494 19540 43546
rect 19564 43494 19594 43546
rect 19594 43494 19606 43546
rect 19606 43494 19620 43546
rect 19644 43494 19658 43546
rect 19658 43494 19670 43546
rect 19670 43494 19700 43546
rect 19724 43494 19734 43546
rect 19734 43494 19780 43546
rect 19484 43492 19540 43494
rect 19564 43492 19620 43494
rect 19644 43492 19700 43494
rect 19724 43492 19780 43494
rect 19484 42458 19540 42460
rect 19564 42458 19620 42460
rect 19644 42458 19700 42460
rect 19724 42458 19780 42460
rect 19484 42406 19530 42458
rect 19530 42406 19540 42458
rect 19564 42406 19594 42458
rect 19594 42406 19606 42458
rect 19606 42406 19620 42458
rect 19644 42406 19658 42458
rect 19658 42406 19670 42458
rect 19670 42406 19700 42458
rect 19724 42406 19734 42458
rect 19734 42406 19780 42458
rect 19484 42404 19540 42406
rect 19564 42404 19620 42406
rect 19644 42404 19700 42406
rect 19724 42404 19780 42406
rect 19484 41370 19540 41372
rect 19564 41370 19620 41372
rect 19644 41370 19700 41372
rect 19724 41370 19780 41372
rect 19484 41318 19530 41370
rect 19530 41318 19540 41370
rect 19564 41318 19594 41370
rect 19594 41318 19606 41370
rect 19606 41318 19620 41370
rect 19644 41318 19658 41370
rect 19658 41318 19670 41370
rect 19670 41318 19700 41370
rect 19724 41318 19734 41370
rect 19734 41318 19780 41370
rect 19484 41316 19540 41318
rect 19564 41316 19620 41318
rect 19644 41316 19700 41318
rect 19724 41316 19780 41318
rect 19484 40282 19540 40284
rect 19564 40282 19620 40284
rect 19644 40282 19700 40284
rect 19724 40282 19780 40284
rect 19484 40230 19530 40282
rect 19530 40230 19540 40282
rect 19564 40230 19594 40282
rect 19594 40230 19606 40282
rect 19606 40230 19620 40282
rect 19644 40230 19658 40282
rect 19658 40230 19670 40282
rect 19670 40230 19700 40282
rect 19724 40230 19734 40282
rect 19734 40230 19780 40282
rect 19484 40228 19540 40230
rect 19564 40228 19620 40230
rect 19644 40228 19700 40230
rect 19724 40228 19780 40230
rect 19484 39194 19540 39196
rect 19564 39194 19620 39196
rect 19644 39194 19700 39196
rect 19724 39194 19780 39196
rect 19484 39142 19530 39194
rect 19530 39142 19540 39194
rect 19564 39142 19594 39194
rect 19594 39142 19606 39194
rect 19606 39142 19620 39194
rect 19644 39142 19658 39194
rect 19658 39142 19670 39194
rect 19670 39142 19700 39194
rect 19724 39142 19734 39194
rect 19734 39142 19780 39194
rect 19484 39140 19540 39142
rect 19564 39140 19620 39142
rect 19644 39140 19700 39142
rect 19724 39140 19780 39142
rect 10220 31578 10276 31580
rect 10300 31578 10356 31580
rect 10380 31578 10436 31580
rect 10460 31578 10516 31580
rect 10220 31526 10266 31578
rect 10266 31526 10276 31578
rect 10300 31526 10330 31578
rect 10330 31526 10342 31578
rect 10342 31526 10356 31578
rect 10380 31526 10394 31578
rect 10394 31526 10406 31578
rect 10406 31526 10436 31578
rect 10460 31526 10470 31578
rect 10470 31526 10516 31578
rect 10220 31524 10276 31526
rect 10300 31524 10356 31526
rect 10380 31524 10436 31526
rect 10460 31524 10516 31526
rect 14852 31034 14908 31036
rect 14932 31034 14988 31036
rect 15012 31034 15068 31036
rect 15092 31034 15148 31036
rect 14852 30982 14898 31034
rect 14898 30982 14908 31034
rect 14932 30982 14962 31034
rect 14962 30982 14974 31034
rect 14974 30982 14988 31034
rect 15012 30982 15026 31034
rect 15026 30982 15038 31034
rect 15038 30982 15068 31034
rect 15092 30982 15102 31034
rect 15102 30982 15148 31034
rect 14852 30980 14908 30982
rect 14932 30980 14988 30982
rect 15012 30980 15068 30982
rect 15092 30980 15148 30982
rect 10220 30490 10276 30492
rect 10300 30490 10356 30492
rect 10380 30490 10436 30492
rect 10460 30490 10516 30492
rect 10220 30438 10266 30490
rect 10266 30438 10276 30490
rect 10300 30438 10330 30490
rect 10330 30438 10342 30490
rect 10342 30438 10356 30490
rect 10380 30438 10394 30490
rect 10394 30438 10406 30490
rect 10406 30438 10436 30490
rect 10460 30438 10470 30490
rect 10470 30438 10516 30490
rect 10220 30436 10276 30438
rect 10300 30436 10356 30438
rect 10380 30436 10436 30438
rect 10460 30436 10516 30438
rect 10220 29402 10276 29404
rect 10300 29402 10356 29404
rect 10380 29402 10436 29404
rect 10460 29402 10516 29404
rect 10220 29350 10266 29402
rect 10266 29350 10276 29402
rect 10300 29350 10330 29402
rect 10330 29350 10342 29402
rect 10342 29350 10356 29402
rect 10380 29350 10394 29402
rect 10394 29350 10406 29402
rect 10406 29350 10436 29402
rect 10460 29350 10470 29402
rect 10470 29350 10516 29402
rect 10220 29348 10276 29350
rect 10300 29348 10356 29350
rect 10380 29348 10436 29350
rect 10460 29348 10516 29350
rect 10220 28314 10276 28316
rect 10300 28314 10356 28316
rect 10380 28314 10436 28316
rect 10460 28314 10516 28316
rect 10220 28262 10266 28314
rect 10266 28262 10276 28314
rect 10300 28262 10330 28314
rect 10330 28262 10342 28314
rect 10342 28262 10356 28314
rect 10380 28262 10394 28314
rect 10394 28262 10406 28314
rect 10406 28262 10436 28314
rect 10460 28262 10470 28314
rect 10470 28262 10516 28314
rect 10220 28260 10276 28262
rect 10300 28260 10356 28262
rect 10380 28260 10436 28262
rect 10460 28260 10516 28262
rect 10220 27226 10276 27228
rect 10300 27226 10356 27228
rect 10380 27226 10436 27228
rect 10460 27226 10516 27228
rect 10220 27174 10266 27226
rect 10266 27174 10276 27226
rect 10300 27174 10330 27226
rect 10330 27174 10342 27226
rect 10342 27174 10356 27226
rect 10380 27174 10394 27226
rect 10394 27174 10406 27226
rect 10406 27174 10436 27226
rect 10460 27174 10470 27226
rect 10470 27174 10516 27226
rect 10220 27172 10276 27174
rect 10300 27172 10356 27174
rect 10380 27172 10436 27174
rect 10460 27172 10516 27174
rect 10220 26138 10276 26140
rect 10300 26138 10356 26140
rect 10380 26138 10436 26140
rect 10460 26138 10516 26140
rect 10220 26086 10266 26138
rect 10266 26086 10276 26138
rect 10300 26086 10330 26138
rect 10330 26086 10342 26138
rect 10342 26086 10356 26138
rect 10380 26086 10394 26138
rect 10394 26086 10406 26138
rect 10406 26086 10436 26138
rect 10460 26086 10470 26138
rect 10470 26086 10516 26138
rect 10220 26084 10276 26086
rect 10300 26084 10356 26086
rect 10380 26084 10436 26086
rect 10460 26084 10516 26086
rect 10220 25050 10276 25052
rect 10300 25050 10356 25052
rect 10380 25050 10436 25052
rect 10460 25050 10516 25052
rect 10220 24998 10266 25050
rect 10266 24998 10276 25050
rect 10300 24998 10330 25050
rect 10330 24998 10342 25050
rect 10342 24998 10356 25050
rect 10380 24998 10394 25050
rect 10394 24998 10406 25050
rect 10406 24998 10436 25050
rect 10460 24998 10470 25050
rect 10470 24998 10516 25050
rect 10220 24996 10276 24998
rect 10300 24996 10356 24998
rect 10380 24996 10436 24998
rect 10460 24996 10516 24998
rect 10220 23962 10276 23964
rect 10300 23962 10356 23964
rect 10380 23962 10436 23964
rect 10460 23962 10516 23964
rect 10220 23910 10266 23962
rect 10266 23910 10276 23962
rect 10300 23910 10330 23962
rect 10330 23910 10342 23962
rect 10342 23910 10356 23962
rect 10380 23910 10394 23962
rect 10394 23910 10406 23962
rect 10406 23910 10436 23962
rect 10460 23910 10470 23962
rect 10470 23910 10516 23962
rect 10220 23908 10276 23910
rect 10300 23908 10356 23910
rect 10380 23908 10436 23910
rect 10460 23908 10516 23910
rect 5588 15802 5644 15804
rect 5668 15802 5724 15804
rect 5748 15802 5804 15804
rect 5828 15802 5884 15804
rect 5588 15750 5634 15802
rect 5634 15750 5644 15802
rect 5668 15750 5698 15802
rect 5698 15750 5710 15802
rect 5710 15750 5724 15802
rect 5748 15750 5762 15802
rect 5762 15750 5774 15802
rect 5774 15750 5804 15802
rect 5828 15750 5838 15802
rect 5838 15750 5884 15802
rect 5588 15748 5644 15750
rect 5668 15748 5724 15750
rect 5748 15748 5804 15750
rect 5828 15748 5884 15750
rect 5588 14714 5644 14716
rect 5668 14714 5724 14716
rect 5748 14714 5804 14716
rect 5828 14714 5884 14716
rect 5588 14662 5634 14714
rect 5634 14662 5644 14714
rect 5668 14662 5698 14714
rect 5698 14662 5710 14714
rect 5710 14662 5724 14714
rect 5748 14662 5762 14714
rect 5762 14662 5774 14714
rect 5774 14662 5804 14714
rect 5828 14662 5838 14714
rect 5838 14662 5884 14714
rect 5588 14660 5644 14662
rect 5668 14660 5724 14662
rect 5748 14660 5804 14662
rect 5828 14660 5884 14662
rect 5588 13626 5644 13628
rect 5668 13626 5724 13628
rect 5748 13626 5804 13628
rect 5828 13626 5884 13628
rect 5588 13574 5634 13626
rect 5634 13574 5644 13626
rect 5668 13574 5698 13626
rect 5698 13574 5710 13626
rect 5710 13574 5724 13626
rect 5748 13574 5762 13626
rect 5762 13574 5774 13626
rect 5774 13574 5804 13626
rect 5828 13574 5838 13626
rect 5838 13574 5884 13626
rect 5588 13572 5644 13574
rect 5668 13572 5724 13574
rect 5748 13572 5804 13574
rect 5828 13572 5884 13574
rect 5588 12538 5644 12540
rect 5668 12538 5724 12540
rect 5748 12538 5804 12540
rect 5828 12538 5884 12540
rect 5588 12486 5634 12538
rect 5634 12486 5644 12538
rect 5668 12486 5698 12538
rect 5698 12486 5710 12538
rect 5710 12486 5724 12538
rect 5748 12486 5762 12538
rect 5762 12486 5774 12538
rect 5774 12486 5804 12538
rect 5828 12486 5838 12538
rect 5838 12486 5884 12538
rect 5588 12484 5644 12486
rect 5668 12484 5724 12486
rect 5748 12484 5804 12486
rect 5828 12484 5884 12486
rect 5588 11450 5644 11452
rect 5668 11450 5724 11452
rect 5748 11450 5804 11452
rect 5828 11450 5884 11452
rect 5588 11398 5634 11450
rect 5634 11398 5644 11450
rect 5668 11398 5698 11450
rect 5698 11398 5710 11450
rect 5710 11398 5724 11450
rect 5748 11398 5762 11450
rect 5762 11398 5774 11450
rect 5774 11398 5804 11450
rect 5828 11398 5838 11450
rect 5838 11398 5884 11450
rect 5588 11396 5644 11398
rect 5668 11396 5724 11398
rect 5748 11396 5804 11398
rect 5828 11396 5884 11398
rect 5588 10362 5644 10364
rect 5668 10362 5724 10364
rect 5748 10362 5804 10364
rect 5828 10362 5884 10364
rect 5588 10310 5634 10362
rect 5634 10310 5644 10362
rect 5668 10310 5698 10362
rect 5698 10310 5710 10362
rect 5710 10310 5724 10362
rect 5748 10310 5762 10362
rect 5762 10310 5774 10362
rect 5774 10310 5804 10362
rect 5828 10310 5838 10362
rect 5838 10310 5884 10362
rect 5588 10308 5644 10310
rect 5668 10308 5724 10310
rect 5748 10308 5804 10310
rect 5828 10308 5884 10310
rect 5588 9274 5644 9276
rect 5668 9274 5724 9276
rect 5748 9274 5804 9276
rect 5828 9274 5884 9276
rect 5588 9222 5634 9274
rect 5634 9222 5644 9274
rect 5668 9222 5698 9274
rect 5698 9222 5710 9274
rect 5710 9222 5724 9274
rect 5748 9222 5762 9274
rect 5762 9222 5774 9274
rect 5774 9222 5804 9274
rect 5828 9222 5838 9274
rect 5838 9222 5884 9274
rect 5588 9220 5644 9222
rect 5668 9220 5724 9222
rect 5748 9220 5804 9222
rect 5828 9220 5884 9222
rect 5588 8186 5644 8188
rect 5668 8186 5724 8188
rect 5748 8186 5804 8188
rect 5828 8186 5884 8188
rect 5588 8134 5634 8186
rect 5634 8134 5644 8186
rect 5668 8134 5698 8186
rect 5698 8134 5710 8186
rect 5710 8134 5724 8186
rect 5748 8134 5762 8186
rect 5762 8134 5774 8186
rect 5774 8134 5804 8186
rect 5828 8134 5838 8186
rect 5838 8134 5884 8186
rect 5588 8132 5644 8134
rect 5668 8132 5724 8134
rect 5748 8132 5804 8134
rect 5828 8132 5884 8134
rect 5588 7098 5644 7100
rect 5668 7098 5724 7100
rect 5748 7098 5804 7100
rect 5828 7098 5884 7100
rect 5588 7046 5634 7098
rect 5634 7046 5644 7098
rect 5668 7046 5698 7098
rect 5698 7046 5710 7098
rect 5710 7046 5724 7098
rect 5748 7046 5762 7098
rect 5762 7046 5774 7098
rect 5774 7046 5804 7098
rect 5828 7046 5838 7098
rect 5838 7046 5884 7098
rect 5588 7044 5644 7046
rect 5668 7044 5724 7046
rect 5748 7044 5804 7046
rect 5828 7044 5884 7046
rect 5588 6010 5644 6012
rect 5668 6010 5724 6012
rect 5748 6010 5804 6012
rect 5828 6010 5884 6012
rect 5588 5958 5634 6010
rect 5634 5958 5644 6010
rect 5668 5958 5698 6010
rect 5698 5958 5710 6010
rect 5710 5958 5724 6010
rect 5748 5958 5762 6010
rect 5762 5958 5774 6010
rect 5774 5958 5804 6010
rect 5828 5958 5838 6010
rect 5838 5958 5884 6010
rect 5588 5956 5644 5958
rect 5668 5956 5724 5958
rect 5748 5956 5804 5958
rect 5828 5956 5884 5958
rect 5588 4922 5644 4924
rect 5668 4922 5724 4924
rect 5748 4922 5804 4924
rect 5828 4922 5884 4924
rect 5588 4870 5634 4922
rect 5634 4870 5644 4922
rect 5668 4870 5698 4922
rect 5698 4870 5710 4922
rect 5710 4870 5724 4922
rect 5748 4870 5762 4922
rect 5762 4870 5774 4922
rect 5774 4870 5804 4922
rect 5828 4870 5838 4922
rect 5838 4870 5884 4922
rect 5588 4868 5644 4870
rect 5668 4868 5724 4870
rect 5748 4868 5804 4870
rect 5828 4868 5884 4870
rect 5588 3834 5644 3836
rect 5668 3834 5724 3836
rect 5748 3834 5804 3836
rect 5828 3834 5884 3836
rect 5588 3782 5634 3834
rect 5634 3782 5644 3834
rect 5668 3782 5698 3834
rect 5698 3782 5710 3834
rect 5710 3782 5724 3834
rect 5748 3782 5762 3834
rect 5762 3782 5774 3834
rect 5774 3782 5804 3834
rect 5828 3782 5838 3834
rect 5838 3782 5884 3834
rect 5588 3780 5644 3782
rect 5668 3780 5724 3782
rect 5748 3780 5804 3782
rect 5828 3780 5884 3782
rect 3422 2080 3478 2136
rect 3330 1400 3386 1456
rect 5588 2746 5644 2748
rect 5668 2746 5724 2748
rect 5748 2746 5804 2748
rect 5828 2746 5884 2748
rect 5588 2694 5634 2746
rect 5634 2694 5644 2746
rect 5668 2694 5698 2746
rect 5698 2694 5710 2746
rect 5710 2694 5724 2746
rect 5748 2694 5762 2746
rect 5762 2694 5774 2746
rect 5774 2694 5804 2746
rect 5828 2694 5838 2746
rect 5838 2694 5884 2746
rect 5588 2692 5644 2694
rect 5668 2692 5724 2694
rect 5748 2692 5804 2694
rect 5828 2692 5884 2694
rect 10220 22874 10276 22876
rect 10300 22874 10356 22876
rect 10380 22874 10436 22876
rect 10460 22874 10516 22876
rect 10220 22822 10266 22874
rect 10266 22822 10276 22874
rect 10300 22822 10330 22874
rect 10330 22822 10342 22874
rect 10342 22822 10356 22874
rect 10380 22822 10394 22874
rect 10394 22822 10406 22874
rect 10406 22822 10436 22874
rect 10460 22822 10470 22874
rect 10470 22822 10516 22874
rect 10220 22820 10276 22822
rect 10300 22820 10356 22822
rect 10380 22820 10436 22822
rect 10460 22820 10516 22822
rect 10220 21786 10276 21788
rect 10300 21786 10356 21788
rect 10380 21786 10436 21788
rect 10460 21786 10516 21788
rect 10220 21734 10266 21786
rect 10266 21734 10276 21786
rect 10300 21734 10330 21786
rect 10330 21734 10342 21786
rect 10342 21734 10356 21786
rect 10380 21734 10394 21786
rect 10394 21734 10406 21786
rect 10406 21734 10436 21786
rect 10460 21734 10470 21786
rect 10470 21734 10516 21786
rect 10220 21732 10276 21734
rect 10300 21732 10356 21734
rect 10380 21732 10436 21734
rect 10460 21732 10516 21734
rect 10220 20698 10276 20700
rect 10300 20698 10356 20700
rect 10380 20698 10436 20700
rect 10460 20698 10516 20700
rect 10220 20646 10266 20698
rect 10266 20646 10276 20698
rect 10300 20646 10330 20698
rect 10330 20646 10342 20698
rect 10342 20646 10356 20698
rect 10380 20646 10394 20698
rect 10394 20646 10406 20698
rect 10406 20646 10436 20698
rect 10460 20646 10470 20698
rect 10470 20646 10516 20698
rect 10220 20644 10276 20646
rect 10300 20644 10356 20646
rect 10380 20644 10436 20646
rect 10460 20644 10516 20646
rect 10220 19610 10276 19612
rect 10300 19610 10356 19612
rect 10380 19610 10436 19612
rect 10460 19610 10516 19612
rect 10220 19558 10266 19610
rect 10266 19558 10276 19610
rect 10300 19558 10330 19610
rect 10330 19558 10342 19610
rect 10342 19558 10356 19610
rect 10380 19558 10394 19610
rect 10394 19558 10406 19610
rect 10406 19558 10436 19610
rect 10460 19558 10470 19610
rect 10470 19558 10516 19610
rect 10220 19556 10276 19558
rect 10300 19556 10356 19558
rect 10380 19556 10436 19558
rect 10460 19556 10516 19558
rect 10220 18522 10276 18524
rect 10300 18522 10356 18524
rect 10380 18522 10436 18524
rect 10460 18522 10516 18524
rect 10220 18470 10266 18522
rect 10266 18470 10276 18522
rect 10300 18470 10330 18522
rect 10330 18470 10342 18522
rect 10342 18470 10356 18522
rect 10380 18470 10394 18522
rect 10394 18470 10406 18522
rect 10406 18470 10436 18522
rect 10460 18470 10470 18522
rect 10470 18470 10516 18522
rect 10220 18468 10276 18470
rect 10300 18468 10356 18470
rect 10380 18468 10436 18470
rect 10460 18468 10516 18470
rect 14852 29946 14908 29948
rect 14932 29946 14988 29948
rect 15012 29946 15068 29948
rect 15092 29946 15148 29948
rect 14852 29894 14898 29946
rect 14898 29894 14908 29946
rect 14932 29894 14962 29946
rect 14962 29894 14974 29946
rect 14974 29894 14988 29946
rect 15012 29894 15026 29946
rect 15026 29894 15038 29946
rect 15038 29894 15068 29946
rect 15092 29894 15102 29946
rect 15102 29894 15148 29946
rect 14852 29892 14908 29894
rect 14932 29892 14988 29894
rect 15012 29892 15068 29894
rect 15092 29892 15148 29894
rect 14852 28858 14908 28860
rect 14932 28858 14988 28860
rect 15012 28858 15068 28860
rect 15092 28858 15148 28860
rect 14852 28806 14898 28858
rect 14898 28806 14908 28858
rect 14932 28806 14962 28858
rect 14962 28806 14974 28858
rect 14974 28806 14988 28858
rect 15012 28806 15026 28858
rect 15026 28806 15038 28858
rect 15038 28806 15068 28858
rect 15092 28806 15102 28858
rect 15102 28806 15148 28858
rect 14852 28804 14908 28806
rect 14932 28804 14988 28806
rect 15012 28804 15068 28806
rect 15092 28804 15148 28806
rect 14852 27770 14908 27772
rect 14932 27770 14988 27772
rect 15012 27770 15068 27772
rect 15092 27770 15148 27772
rect 14852 27718 14898 27770
rect 14898 27718 14908 27770
rect 14932 27718 14962 27770
rect 14962 27718 14974 27770
rect 14974 27718 14988 27770
rect 15012 27718 15026 27770
rect 15026 27718 15038 27770
rect 15038 27718 15068 27770
rect 15092 27718 15102 27770
rect 15102 27718 15148 27770
rect 14852 27716 14908 27718
rect 14932 27716 14988 27718
rect 15012 27716 15068 27718
rect 15092 27716 15148 27718
rect 14852 26682 14908 26684
rect 14932 26682 14988 26684
rect 15012 26682 15068 26684
rect 15092 26682 15148 26684
rect 14852 26630 14898 26682
rect 14898 26630 14908 26682
rect 14932 26630 14962 26682
rect 14962 26630 14974 26682
rect 14974 26630 14988 26682
rect 15012 26630 15026 26682
rect 15026 26630 15038 26682
rect 15038 26630 15068 26682
rect 15092 26630 15102 26682
rect 15102 26630 15148 26682
rect 14852 26628 14908 26630
rect 14932 26628 14988 26630
rect 15012 26628 15068 26630
rect 15092 26628 15148 26630
rect 14852 25594 14908 25596
rect 14932 25594 14988 25596
rect 15012 25594 15068 25596
rect 15092 25594 15148 25596
rect 14852 25542 14898 25594
rect 14898 25542 14908 25594
rect 14932 25542 14962 25594
rect 14962 25542 14974 25594
rect 14974 25542 14988 25594
rect 15012 25542 15026 25594
rect 15026 25542 15038 25594
rect 15038 25542 15068 25594
rect 15092 25542 15102 25594
rect 15102 25542 15148 25594
rect 14852 25540 14908 25542
rect 14932 25540 14988 25542
rect 15012 25540 15068 25542
rect 15092 25540 15148 25542
rect 14852 24506 14908 24508
rect 14932 24506 14988 24508
rect 15012 24506 15068 24508
rect 15092 24506 15148 24508
rect 14852 24454 14898 24506
rect 14898 24454 14908 24506
rect 14932 24454 14962 24506
rect 14962 24454 14974 24506
rect 14974 24454 14988 24506
rect 15012 24454 15026 24506
rect 15026 24454 15038 24506
rect 15038 24454 15068 24506
rect 15092 24454 15102 24506
rect 15102 24454 15148 24506
rect 14852 24452 14908 24454
rect 14932 24452 14988 24454
rect 15012 24452 15068 24454
rect 15092 24452 15148 24454
rect 14852 23418 14908 23420
rect 14932 23418 14988 23420
rect 15012 23418 15068 23420
rect 15092 23418 15148 23420
rect 14852 23366 14898 23418
rect 14898 23366 14908 23418
rect 14932 23366 14962 23418
rect 14962 23366 14974 23418
rect 14974 23366 14988 23418
rect 15012 23366 15026 23418
rect 15026 23366 15038 23418
rect 15038 23366 15068 23418
rect 15092 23366 15102 23418
rect 15102 23366 15148 23418
rect 14852 23364 14908 23366
rect 14932 23364 14988 23366
rect 15012 23364 15068 23366
rect 15092 23364 15148 23366
rect 14852 22330 14908 22332
rect 14932 22330 14988 22332
rect 15012 22330 15068 22332
rect 15092 22330 15148 22332
rect 14852 22278 14898 22330
rect 14898 22278 14908 22330
rect 14932 22278 14962 22330
rect 14962 22278 14974 22330
rect 14974 22278 14988 22330
rect 15012 22278 15026 22330
rect 15026 22278 15038 22330
rect 15038 22278 15068 22330
rect 15092 22278 15102 22330
rect 15102 22278 15148 22330
rect 14852 22276 14908 22278
rect 14932 22276 14988 22278
rect 15012 22276 15068 22278
rect 15092 22276 15148 22278
rect 10220 17434 10276 17436
rect 10300 17434 10356 17436
rect 10380 17434 10436 17436
rect 10460 17434 10516 17436
rect 10220 17382 10266 17434
rect 10266 17382 10276 17434
rect 10300 17382 10330 17434
rect 10330 17382 10342 17434
rect 10342 17382 10356 17434
rect 10380 17382 10394 17434
rect 10394 17382 10406 17434
rect 10406 17382 10436 17434
rect 10460 17382 10470 17434
rect 10470 17382 10516 17434
rect 10220 17380 10276 17382
rect 10300 17380 10356 17382
rect 10380 17380 10436 17382
rect 10460 17380 10516 17382
rect 10220 16346 10276 16348
rect 10300 16346 10356 16348
rect 10380 16346 10436 16348
rect 10460 16346 10516 16348
rect 10220 16294 10266 16346
rect 10266 16294 10276 16346
rect 10300 16294 10330 16346
rect 10330 16294 10342 16346
rect 10342 16294 10356 16346
rect 10380 16294 10394 16346
rect 10394 16294 10406 16346
rect 10406 16294 10436 16346
rect 10460 16294 10470 16346
rect 10470 16294 10516 16346
rect 10220 16292 10276 16294
rect 10300 16292 10356 16294
rect 10380 16292 10436 16294
rect 10460 16292 10516 16294
rect 10220 15258 10276 15260
rect 10300 15258 10356 15260
rect 10380 15258 10436 15260
rect 10460 15258 10516 15260
rect 10220 15206 10266 15258
rect 10266 15206 10276 15258
rect 10300 15206 10330 15258
rect 10330 15206 10342 15258
rect 10342 15206 10356 15258
rect 10380 15206 10394 15258
rect 10394 15206 10406 15258
rect 10406 15206 10436 15258
rect 10460 15206 10470 15258
rect 10470 15206 10516 15258
rect 10220 15204 10276 15206
rect 10300 15204 10356 15206
rect 10380 15204 10436 15206
rect 10460 15204 10516 15206
rect 10220 14170 10276 14172
rect 10300 14170 10356 14172
rect 10380 14170 10436 14172
rect 10460 14170 10516 14172
rect 10220 14118 10266 14170
rect 10266 14118 10276 14170
rect 10300 14118 10330 14170
rect 10330 14118 10342 14170
rect 10342 14118 10356 14170
rect 10380 14118 10394 14170
rect 10394 14118 10406 14170
rect 10406 14118 10436 14170
rect 10460 14118 10470 14170
rect 10470 14118 10516 14170
rect 10220 14116 10276 14118
rect 10300 14116 10356 14118
rect 10380 14116 10436 14118
rect 10460 14116 10516 14118
rect 10220 13082 10276 13084
rect 10300 13082 10356 13084
rect 10380 13082 10436 13084
rect 10460 13082 10516 13084
rect 10220 13030 10266 13082
rect 10266 13030 10276 13082
rect 10300 13030 10330 13082
rect 10330 13030 10342 13082
rect 10342 13030 10356 13082
rect 10380 13030 10394 13082
rect 10394 13030 10406 13082
rect 10406 13030 10436 13082
rect 10460 13030 10470 13082
rect 10470 13030 10516 13082
rect 10220 13028 10276 13030
rect 10300 13028 10356 13030
rect 10380 13028 10436 13030
rect 10460 13028 10516 13030
rect 10220 11994 10276 11996
rect 10300 11994 10356 11996
rect 10380 11994 10436 11996
rect 10460 11994 10516 11996
rect 10220 11942 10266 11994
rect 10266 11942 10276 11994
rect 10300 11942 10330 11994
rect 10330 11942 10342 11994
rect 10342 11942 10356 11994
rect 10380 11942 10394 11994
rect 10394 11942 10406 11994
rect 10406 11942 10436 11994
rect 10460 11942 10470 11994
rect 10470 11942 10516 11994
rect 10220 11940 10276 11942
rect 10300 11940 10356 11942
rect 10380 11940 10436 11942
rect 10460 11940 10516 11942
rect 14852 21242 14908 21244
rect 14932 21242 14988 21244
rect 15012 21242 15068 21244
rect 15092 21242 15148 21244
rect 14852 21190 14898 21242
rect 14898 21190 14908 21242
rect 14932 21190 14962 21242
rect 14962 21190 14974 21242
rect 14974 21190 14988 21242
rect 15012 21190 15026 21242
rect 15026 21190 15038 21242
rect 15038 21190 15068 21242
rect 15092 21190 15102 21242
rect 15102 21190 15148 21242
rect 14852 21188 14908 21190
rect 14932 21188 14988 21190
rect 15012 21188 15068 21190
rect 15092 21188 15148 21190
rect 14852 20154 14908 20156
rect 14932 20154 14988 20156
rect 15012 20154 15068 20156
rect 15092 20154 15148 20156
rect 14852 20102 14898 20154
rect 14898 20102 14908 20154
rect 14932 20102 14962 20154
rect 14962 20102 14974 20154
rect 14974 20102 14988 20154
rect 15012 20102 15026 20154
rect 15026 20102 15038 20154
rect 15038 20102 15068 20154
rect 15092 20102 15102 20154
rect 15102 20102 15148 20154
rect 14852 20100 14908 20102
rect 14932 20100 14988 20102
rect 15012 20100 15068 20102
rect 15092 20100 15148 20102
rect 14852 19066 14908 19068
rect 14932 19066 14988 19068
rect 15012 19066 15068 19068
rect 15092 19066 15148 19068
rect 14852 19014 14898 19066
rect 14898 19014 14908 19066
rect 14932 19014 14962 19066
rect 14962 19014 14974 19066
rect 14974 19014 14988 19066
rect 15012 19014 15026 19066
rect 15026 19014 15038 19066
rect 15038 19014 15068 19066
rect 15092 19014 15102 19066
rect 15102 19014 15148 19066
rect 14852 19012 14908 19014
rect 14932 19012 14988 19014
rect 15012 19012 15068 19014
rect 15092 19012 15148 19014
rect 14852 17978 14908 17980
rect 14932 17978 14988 17980
rect 15012 17978 15068 17980
rect 15092 17978 15148 17980
rect 14852 17926 14898 17978
rect 14898 17926 14908 17978
rect 14932 17926 14962 17978
rect 14962 17926 14974 17978
rect 14974 17926 14988 17978
rect 15012 17926 15026 17978
rect 15026 17926 15038 17978
rect 15038 17926 15068 17978
rect 15092 17926 15102 17978
rect 15102 17926 15148 17978
rect 14852 17924 14908 17926
rect 14932 17924 14988 17926
rect 15012 17924 15068 17926
rect 15092 17924 15148 17926
rect 14852 16890 14908 16892
rect 14932 16890 14988 16892
rect 15012 16890 15068 16892
rect 15092 16890 15148 16892
rect 14852 16838 14898 16890
rect 14898 16838 14908 16890
rect 14932 16838 14962 16890
rect 14962 16838 14974 16890
rect 14974 16838 14988 16890
rect 15012 16838 15026 16890
rect 15026 16838 15038 16890
rect 15038 16838 15068 16890
rect 15092 16838 15102 16890
rect 15102 16838 15148 16890
rect 14852 16836 14908 16838
rect 14932 16836 14988 16838
rect 15012 16836 15068 16838
rect 15092 16836 15148 16838
rect 14852 15802 14908 15804
rect 14932 15802 14988 15804
rect 15012 15802 15068 15804
rect 15092 15802 15148 15804
rect 14852 15750 14898 15802
rect 14898 15750 14908 15802
rect 14932 15750 14962 15802
rect 14962 15750 14974 15802
rect 14974 15750 14988 15802
rect 15012 15750 15026 15802
rect 15026 15750 15038 15802
rect 15038 15750 15068 15802
rect 15092 15750 15102 15802
rect 15102 15750 15148 15802
rect 14852 15748 14908 15750
rect 14932 15748 14988 15750
rect 15012 15748 15068 15750
rect 15092 15748 15148 15750
rect 14852 14714 14908 14716
rect 14932 14714 14988 14716
rect 15012 14714 15068 14716
rect 15092 14714 15148 14716
rect 14852 14662 14898 14714
rect 14898 14662 14908 14714
rect 14932 14662 14962 14714
rect 14962 14662 14974 14714
rect 14974 14662 14988 14714
rect 15012 14662 15026 14714
rect 15026 14662 15038 14714
rect 15038 14662 15068 14714
rect 15092 14662 15102 14714
rect 15102 14662 15148 14714
rect 14852 14660 14908 14662
rect 14932 14660 14988 14662
rect 15012 14660 15068 14662
rect 15092 14660 15148 14662
rect 14852 13626 14908 13628
rect 14932 13626 14988 13628
rect 15012 13626 15068 13628
rect 15092 13626 15148 13628
rect 14852 13574 14898 13626
rect 14898 13574 14908 13626
rect 14932 13574 14962 13626
rect 14962 13574 14974 13626
rect 14974 13574 14988 13626
rect 15012 13574 15026 13626
rect 15026 13574 15038 13626
rect 15038 13574 15068 13626
rect 15092 13574 15102 13626
rect 15102 13574 15148 13626
rect 14852 13572 14908 13574
rect 14932 13572 14988 13574
rect 15012 13572 15068 13574
rect 15092 13572 15148 13574
rect 14852 12538 14908 12540
rect 14932 12538 14988 12540
rect 15012 12538 15068 12540
rect 15092 12538 15148 12540
rect 14852 12486 14898 12538
rect 14898 12486 14908 12538
rect 14932 12486 14962 12538
rect 14962 12486 14974 12538
rect 14974 12486 14988 12538
rect 15012 12486 15026 12538
rect 15026 12486 15038 12538
rect 15038 12486 15068 12538
rect 15092 12486 15102 12538
rect 15102 12486 15148 12538
rect 14852 12484 14908 12486
rect 14932 12484 14988 12486
rect 15012 12484 15068 12486
rect 15092 12484 15148 12486
rect 14852 11450 14908 11452
rect 14932 11450 14988 11452
rect 15012 11450 15068 11452
rect 15092 11450 15148 11452
rect 14852 11398 14898 11450
rect 14898 11398 14908 11450
rect 14932 11398 14962 11450
rect 14962 11398 14974 11450
rect 14974 11398 14988 11450
rect 15012 11398 15026 11450
rect 15026 11398 15038 11450
rect 15038 11398 15068 11450
rect 15092 11398 15102 11450
rect 15102 11398 15148 11450
rect 14852 11396 14908 11398
rect 14932 11396 14988 11398
rect 15012 11396 15068 11398
rect 15092 11396 15148 11398
rect 10220 10906 10276 10908
rect 10300 10906 10356 10908
rect 10380 10906 10436 10908
rect 10460 10906 10516 10908
rect 10220 10854 10266 10906
rect 10266 10854 10276 10906
rect 10300 10854 10330 10906
rect 10330 10854 10342 10906
rect 10342 10854 10356 10906
rect 10380 10854 10394 10906
rect 10394 10854 10406 10906
rect 10406 10854 10436 10906
rect 10460 10854 10470 10906
rect 10470 10854 10516 10906
rect 10220 10852 10276 10854
rect 10300 10852 10356 10854
rect 10380 10852 10436 10854
rect 10460 10852 10516 10854
rect 14852 10362 14908 10364
rect 14932 10362 14988 10364
rect 15012 10362 15068 10364
rect 15092 10362 15148 10364
rect 14852 10310 14898 10362
rect 14898 10310 14908 10362
rect 14932 10310 14962 10362
rect 14962 10310 14974 10362
rect 14974 10310 14988 10362
rect 15012 10310 15026 10362
rect 15026 10310 15038 10362
rect 15038 10310 15068 10362
rect 15092 10310 15102 10362
rect 15102 10310 15148 10362
rect 14852 10308 14908 10310
rect 14932 10308 14988 10310
rect 15012 10308 15068 10310
rect 15092 10308 15148 10310
rect 10220 9818 10276 9820
rect 10300 9818 10356 9820
rect 10380 9818 10436 9820
rect 10460 9818 10516 9820
rect 10220 9766 10266 9818
rect 10266 9766 10276 9818
rect 10300 9766 10330 9818
rect 10330 9766 10342 9818
rect 10342 9766 10356 9818
rect 10380 9766 10394 9818
rect 10394 9766 10406 9818
rect 10406 9766 10436 9818
rect 10460 9766 10470 9818
rect 10470 9766 10516 9818
rect 10220 9764 10276 9766
rect 10300 9764 10356 9766
rect 10380 9764 10436 9766
rect 10460 9764 10516 9766
rect 14852 9274 14908 9276
rect 14932 9274 14988 9276
rect 15012 9274 15068 9276
rect 15092 9274 15148 9276
rect 14852 9222 14898 9274
rect 14898 9222 14908 9274
rect 14932 9222 14962 9274
rect 14962 9222 14974 9274
rect 14974 9222 14988 9274
rect 15012 9222 15026 9274
rect 15026 9222 15038 9274
rect 15038 9222 15068 9274
rect 15092 9222 15102 9274
rect 15102 9222 15148 9274
rect 14852 9220 14908 9222
rect 14932 9220 14988 9222
rect 15012 9220 15068 9222
rect 15092 9220 15148 9222
rect 10220 8730 10276 8732
rect 10300 8730 10356 8732
rect 10380 8730 10436 8732
rect 10460 8730 10516 8732
rect 10220 8678 10266 8730
rect 10266 8678 10276 8730
rect 10300 8678 10330 8730
rect 10330 8678 10342 8730
rect 10342 8678 10356 8730
rect 10380 8678 10394 8730
rect 10394 8678 10406 8730
rect 10406 8678 10436 8730
rect 10460 8678 10470 8730
rect 10470 8678 10516 8730
rect 10220 8676 10276 8678
rect 10300 8676 10356 8678
rect 10380 8676 10436 8678
rect 10460 8676 10516 8678
rect 14852 8186 14908 8188
rect 14932 8186 14988 8188
rect 15012 8186 15068 8188
rect 15092 8186 15148 8188
rect 14852 8134 14898 8186
rect 14898 8134 14908 8186
rect 14932 8134 14962 8186
rect 14962 8134 14974 8186
rect 14974 8134 14988 8186
rect 15012 8134 15026 8186
rect 15026 8134 15038 8186
rect 15038 8134 15068 8186
rect 15092 8134 15102 8186
rect 15102 8134 15148 8186
rect 14852 8132 14908 8134
rect 14932 8132 14988 8134
rect 15012 8132 15068 8134
rect 15092 8132 15148 8134
rect 10220 7642 10276 7644
rect 10300 7642 10356 7644
rect 10380 7642 10436 7644
rect 10460 7642 10516 7644
rect 10220 7590 10266 7642
rect 10266 7590 10276 7642
rect 10300 7590 10330 7642
rect 10330 7590 10342 7642
rect 10342 7590 10356 7642
rect 10380 7590 10394 7642
rect 10394 7590 10406 7642
rect 10406 7590 10436 7642
rect 10460 7590 10470 7642
rect 10470 7590 10516 7642
rect 10220 7588 10276 7590
rect 10300 7588 10356 7590
rect 10380 7588 10436 7590
rect 10460 7588 10516 7590
rect 14852 7098 14908 7100
rect 14932 7098 14988 7100
rect 15012 7098 15068 7100
rect 15092 7098 15148 7100
rect 14852 7046 14898 7098
rect 14898 7046 14908 7098
rect 14932 7046 14962 7098
rect 14962 7046 14974 7098
rect 14974 7046 14988 7098
rect 15012 7046 15026 7098
rect 15026 7046 15038 7098
rect 15038 7046 15068 7098
rect 15092 7046 15102 7098
rect 15102 7046 15148 7098
rect 14852 7044 14908 7046
rect 14932 7044 14988 7046
rect 15012 7044 15068 7046
rect 15092 7044 15148 7046
rect 10220 6554 10276 6556
rect 10300 6554 10356 6556
rect 10380 6554 10436 6556
rect 10460 6554 10516 6556
rect 10220 6502 10266 6554
rect 10266 6502 10276 6554
rect 10300 6502 10330 6554
rect 10330 6502 10342 6554
rect 10342 6502 10356 6554
rect 10380 6502 10394 6554
rect 10394 6502 10406 6554
rect 10406 6502 10436 6554
rect 10460 6502 10470 6554
rect 10470 6502 10516 6554
rect 10220 6500 10276 6502
rect 10300 6500 10356 6502
rect 10380 6500 10436 6502
rect 10460 6500 10516 6502
rect 14852 6010 14908 6012
rect 14932 6010 14988 6012
rect 15012 6010 15068 6012
rect 15092 6010 15148 6012
rect 14852 5958 14898 6010
rect 14898 5958 14908 6010
rect 14932 5958 14962 6010
rect 14962 5958 14974 6010
rect 14974 5958 14988 6010
rect 15012 5958 15026 6010
rect 15026 5958 15038 6010
rect 15038 5958 15068 6010
rect 15092 5958 15102 6010
rect 15102 5958 15148 6010
rect 14852 5956 14908 5958
rect 14932 5956 14988 5958
rect 15012 5956 15068 5958
rect 15092 5956 15148 5958
rect 10220 5466 10276 5468
rect 10300 5466 10356 5468
rect 10380 5466 10436 5468
rect 10460 5466 10516 5468
rect 10220 5414 10266 5466
rect 10266 5414 10276 5466
rect 10300 5414 10330 5466
rect 10330 5414 10342 5466
rect 10342 5414 10356 5466
rect 10380 5414 10394 5466
rect 10394 5414 10406 5466
rect 10406 5414 10436 5466
rect 10460 5414 10470 5466
rect 10470 5414 10516 5466
rect 10220 5412 10276 5414
rect 10300 5412 10356 5414
rect 10380 5412 10436 5414
rect 10460 5412 10516 5414
rect 14852 4922 14908 4924
rect 14932 4922 14988 4924
rect 15012 4922 15068 4924
rect 15092 4922 15148 4924
rect 14852 4870 14898 4922
rect 14898 4870 14908 4922
rect 14932 4870 14962 4922
rect 14962 4870 14974 4922
rect 14974 4870 14988 4922
rect 15012 4870 15026 4922
rect 15026 4870 15038 4922
rect 15038 4870 15068 4922
rect 15092 4870 15102 4922
rect 15102 4870 15148 4922
rect 14852 4868 14908 4870
rect 14932 4868 14988 4870
rect 15012 4868 15068 4870
rect 15092 4868 15148 4870
rect 10220 4378 10276 4380
rect 10300 4378 10356 4380
rect 10380 4378 10436 4380
rect 10460 4378 10516 4380
rect 10220 4326 10266 4378
rect 10266 4326 10276 4378
rect 10300 4326 10330 4378
rect 10330 4326 10342 4378
rect 10342 4326 10356 4378
rect 10380 4326 10394 4378
rect 10394 4326 10406 4378
rect 10406 4326 10436 4378
rect 10460 4326 10470 4378
rect 10470 4326 10516 4378
rect 10220 4324 10276 4326
rect 10300 4324 10356 4326
rect 10380 4324 10436 4326
rect 10460 4324 10516 4326
rect 10220 3290 10276 3292
rect 10300 3290 10356 3292
rect 10380 3290 10436 3292
rect 10460 3290 10516 3292
rect 10220 3238 10266 3290
rect 10266 3238 10276 3290
rect 10300 3238 10330 3290
rect 10330 3238 10342 3290
rect 10342 3238 10356 3290
rect 10380 3238 10394 3290
rect 10394 3238 10406 3290
rect 10406 3238 10436 3290
rect 10460 3238 10470 3290
rect 10470 3238 10516 3290
rect 10220 3236 10276 3238
rect 10300 3236 10356 3238
rect 10380 3236 10436 3238
rect 10460 3236 10516 3238
rect 10220 2202 10276 2204
rect 10300 2202 10356 2204
rect 10380 2202 10436 2204
rect 10460 2202 10516 2204
rect 10220 2150 10266 2202
rect 10266 2150 10276 2202
rect 10300 2150 10330 2202
rect 10330 2150 10342 2202
rect 10342 2150 10356 2202
rect 10380 2150 10394 2202
rect 10394 2150 10406 2202
rect 10406 2150 10436 2202
rect 10460 2150 10470 2202
rect 10470 2150 10516 2202
rect 10220 2148 10276 2150
rect 10300 2148 10356 2150
rect 10380 2148 10436 2150
rect 10460 2148 10516 2150
rect 14852 3834 14908 3836
rect 14932 3834 14988 3836
rect 15012 3834 15068 3836
rect 15092 3834 15148 3836
rect 14852 3782 14898 3834
rect 14898 3782 14908 3834
rect 14932 3782 14962 3834
rect 14962 3782 14974 3834
rect 14974 3782 14988 3834
rect 15012 3782 15026 3834
rect 15026 3782 15038 3834
rect 15038 3782 15068 3834
rect 15092 3782 15102 3834
rect 15102 3782 15148 3834
rect 14852 3780 14908 3782
rect 14932 3780 14988 3782
rect 15012 3780 15068 3782
rect 15092 3780 15148 3782
rect 14646 3576 14702 3632
rect 14852 2746 14908 2748
rect 14932 2746 14988 2748
rect 15012 2746 15068 2748
rect 15092 2746 15148 2748
rect 14852 2694 14898 2746
rect 14898 2694 14908 2746
rect 14932 2694 14962 2746
rect 14962 2694 14974 2746
rect 14974 2694 14988 2746
rect 15012 2694 15026 2746
rect 15026 2694 15038 2746
rect 15038 2694 15068 2746
rect 15092 2694 15102 2746
rect 15102 2694 15148 2746
rect 14852 2692 14908 2694
rect 14932 2692 14988 2694
rect 15012 2692 15068 2694
rect 15092 2692 15148 2694
rect 18326 35148 18382 35184
rect 18326 35128 18328 35148
rect 18328 35128 18380 35148
rect 18380 35128 18382 35148
rect 19484 38106 19540 38108
rect 19564 38106 19620 38108
rect 19644 38106 19700 38108
rect 19724 38106 19780 38108
rect 19484 38054 19530 38106
rect 19530 38054 19540 38106
rect 19564 38054 19594 38106
rect 19594 38054 19606 38106
rect 19606 38054 19620 38106
rect 19644 38054 19658 38106
rect 19658 38054 19670 38106
rect 19670 38054 19700 38106
rect 19724 38054 19734 38106
rect 19734 38054 19780 38106
rect 19484 38052 19540 38054
rect 19564 38052 19620 38054
rect 19644 38052 19700 38054
rect 19724 38052 19780 38054
rect 19484 37018 19540 37020
rect 19564 37018 19620 37020
rect 19644 37018 19700 37020
rect 19724 37018 19780 37020
rect 19484 36966 19530 37018
rect 19530 36966 19540 37018
rect 19564 36966 19594 37018
rect 19594 36966 19606 37018
rect 19606 36966 19620 37018
rect 19644 36966 19658 37018
rect 19658 36966 19670 37018
rect 19670 36966 19700 37018
rect 19724 36966 19734 37018
rect 19734 36966 19780 37018
rect 19484 36964 19540 36966
rect 19564 36964 19620 36966
rect 19644 36964 19700 36966
rect 19724 36964 19780 36966
rect 19484 35930 19540 35932
rect 19564 35930 19620 35932
rect 19644 35930 19700 35932
rect 19724 35930 19780 35932
rect 19484 35878 19530 35930
rect 19530 35878 19540 35930
rect 19564 35878 19594 35930
rect 19594 35878 19606 35930
rect 19606 35878 19620 35930
rect 19644 35878 19658 35930
rect 19658 35878 19670 35930
rect 19670 35878 19700 35930
rect 19724 35878 19734 35930
rect 19734 35878 19780 35930
rect 19484 35876 19540 35878
rect 19564 35876 19620 35878
rect 19644 35876 19700 35878
rect 19724 35876 19780 35878
rect 19484 34842 19540 34844
rect 19564 34842 19620 34844
rect 19644 34842 19700 34844
rect 19724 34842 19780 34844
rect 19484 34790 19530 34842
rect 19530 34790 19540 34842
rect 19564 34790 19594 34842
rect 19594 34790 19606 34842
rect 19606 34790 19620 34842
rect 19644 34790 19658 34842
rect 19658 34790 19670 34842
rect 19670 34790 19700 34842
rect 19724 34790 19734 34842
rect 19734 34790 19780 34842
rect 19484 34788 19540 34790
rect 19564 34788 19620 34790
rect 19644 34788 19700 34790
rect 19724 34788 19780 34790
rect 19484 33754 19540 33756
rect 19564 33754 19620 33756
rect 19644 33754 19700 33756
rect 19724 33754 19780 33756
rect 19484 33702 19530 33754
rect 19530 33702 19540 33754
rect 19564 33702 19594 33754
rect 19594 33702 19606 33754
rect 19606 33702 19620 33754
rect 19644 33702 19658 33754
rect 19658 33702 19670 33754
rect 19670 33702 19700 33754
rect 19724 33702 19734 33754
rect 19734 33702 19780 33754
rect 19484 33700 19540 33702
rect 19564 33700 19620 33702
rect 19644 33700 19700 33702
rect 19724 33700 19780 33702
rect 19484 32666 19540 32668
rect 19564 32666 19620 32668
rect 19644 32666 19700 32668
rect 19724 32666 19780 32668
rect 19484 32614 19530 32666
rect 19530 32614 19540 32666
rect 19564 32614 19594 32666
rect 19594 32614 19606 32666
rect 19606 32614 19620 32666
rect 19644 32614 19658 32666
rect 19658 32614 19670 32666
rect 19670 32614 19700 32666
rect 19724 32614 19734 32666
rect 19734 32614 19780 32666
rect 19484 32612 19540 32614
rect 19564 32612 19620 32614
rect 19644 32612 19700 32614
rect 19724 32612 19780 32614
rect 19484 31578 19540 31580
rect 19564 31578 19620 31580
rect 19644 31578 19700 31580
rect 19724 31578 19780 31580
rect 19484 31526 19530 31578
rect 19530 31526 19540 31578
rect 19564 31526 19594 31578
rect 19594 31526 19606 31578
rect 19606 31526 19620 31578
rect 19644 31526 19658 31578
rect 19658 31526 19670 31578
rect 19670 31526 19700 31578
rect 19724 31526 19734 31578
rect 19734 31526 19780 31578
rect 19484 31524 19540 31526
rect 19564 31524 19620 31526
rect 19644 31524 19700 31526
rect 19724 31524 19780 31526
rect 19484 30490 19540 30492
rect 19564 30490 19620 30492
rect 19644 30490 19700 30492
rect 19724 30490 19780 30492
rect 19484 30438 19530 30490
rect 19530 30438 19540 30490
rect 19564 30438 19594 30490
rect 19594 30438 19606 30490
rect 19606 30438 19620 30490
rect 19644 30438 19658 30490
rect 19658 30438 19670 30490
rect 19670 30438 19700 30490
rect 19724 30438 19734 30490
rect 19734 30438 19780 30490
rect 19484 30436 19540 30438
rect 19564 30436 19620 30438
rect 19644 30436 19700 30438
rect 19724 30436 19780 30438
rect 19484 29402 19540 29404
rect 19564 29402 19620 29404
rect 19644 29402 19700 29404
rect 19724 29402 19780 29404
rect 19484 29350 19530 29402
rect 19530 29350 19540 29402
rect 19564 29350 19594 29402
rect 19594 29350 19606 29402
rect 19606 29350 19620 29402
rect 19644 29350 19658 29402
rect 19658 29350 19670 29402
rect 19670 29350 19700 29402
rect 19724 29350 19734 29402
rect 19734 29350 19780 29402
rect 19484 29348 19540 29350
rect 19564 29348 19620 29350
rect 19644 29348 19700 29350
rect 19724 29348 19780 29350
rect 19484 28314 19540 28316
rect 19564 28314 19620 28316
rect 19644 28314 19700 28316
rect 19724 28314 19780 28316
rect 19484 28262 19530 28314
rect 19530 28262 19540 28314
rect 19564 28262 19594 28314
rect 19594 28262 19606 28314
rect 19606 28262 19620 28314
rect 19644 28262 19658 28314
rect 19658 28262 19670 28314
rect 19670 28262 19700 28314
rect 19724 28262 19734 28314
rect 19734 28262 19780 28314
rect 19484 28260 19540 28262
rect 19564 28260 19620 28262
rect 19644 28260 19700 28262
rect 19724 28260 19780 28262
rect 19484 27226 19540 27228
rect 19564 27226 19620 27228
rect 19644 27226 19700 27228
rect 19724 27226 19780 27228
rect 19484 27174 19530 27226
rect 19530 27174 19540 27226
rect 19564 27174 19594 27226
rect 19594 27174 19606 27226
rect 19606 27174 19620 27226
rect 19644 27174 19658 27226
rect 19658 27174 19670 27226
rect 19670 27174 19700 27226
rect 19724 27174 19734 27226
rect 19734 27174 19780 27226
rect 19484 27172 19540 27174
rect 19564 27172 19620 27174
rect 19644 27172 19700 27174
rect 19724 27172 19780 27174
rect 19484 26138 19540 26140
rect 19564 26138 19620 26140
rect 19644 26138 19700 26140
rect 19724 26138 19780 26140
rect 19484 26086 19530 26138
rect 19530 26086 19540 26138
rect 19564 26086 19594 26138
rect 19594 26086 19606 26138
rect 19606 26086 19620 26138
rect 19644 26086 19658 26138
rect 19658 26086 19670 26138
rect 19670 26086 19700 26138
rect 19724 26086 19734 26138
rect 19734 26086 19780 26138
rect 19484 26084 19540 26086
rect 19564 26084 19620 26086
rect 19644 26084 19700 26086
rect 19724 26084 19780 26086
rect 19484 25050 19540 25052
rect 19564 25050 19620 25052
rect 19644 25050 19700 25052
rect 19724 25050 19780 25052
rect 19484 24998 19530 25050
rect 19530 24998 19540 25050
rect 19564 24998 19594 25050
rect 19594 24998 19606 25050
rect 19606 24998 19620 25050
rect 19644 24998 19658 25050
rect 19658 24998 19670 25050
rect 19670 24998 19700 25050
rect 19724 24998 19734 25050
rect 19734 24998 19780 25050
rect 19484 24996 19540 24998
rect 19564 24996 19620 24998
rect 19644 24996 19700 24998
rect 19724 24996 19780 24998
rect 26146 49000 26202 49056
rect 25594 47640 25650 47696
rect 24116 47354 24172 47356
rect 24196 47354 24252 47356
rect 24276 47354 24332 47356
rect 24356 47354 24412 47356
rect 24116 47302 24162 47354
rect 24162 47302 24172 47354
rect 24196 47302 24226 47354
rect 24226 47302 24238 47354
rect 24238 47302 24252 47354
rect 24276 47302 24290 47354
rect 24290 47302 24302 47354
rect 24302 47302 24332 47354
rect 24356 47302 24366 47354
rect 24366 47302 24412 47354
rect 24116 47300 24172 47302
rect 24196 47300 24252 47302
rect 24276 47300 24332 47302
rect 24356 47300 24412 47302
rect 25962 46280 26018 46336
rect 24116 46266 24172 46268
rect 24196 46266 24252 46268
rect 24276 46266 24332 46268
rect 24356 46266 24412 46268
rect 24116 46214 24162 46266
rect 24162 46214 24172 46266
rect 24196 46214 24226 46266
rect 24226 46214 24238 46266
rect 24238 46214 24252 46266
rect 24276 46214 24290 46266
rect 24290 46214 24302 46266
rect 24302 46214 24332 46266
rect 24356 46214 24366 46266
rect 24366 46214 24412 46266
rect 24116 46212 24172 46214
rect 24196 46212 24252 46214
rect 24276 46212 24332 46214
rect 24356 46212 24412 46214
rect 22006 44240 22062 44296
rect 19484 23962 19540 23964
rect 19564 23962 19620 23964
rect 19644 23962 19700 23964
rect 19724 23962 19780 23964
rect 19484 23910 19530 23962
rect 19530 23910 19540 23962
rect 19564 23910 19594 23962
rect 19594 23910 19606 23962
rect 19606 23910 19620 23962
rect 19644 23910 19658 23962
rect 19658 23910 19670 23962
rect 19670 23910 19700 23962
rect 19724 23910 19734 23962
rect 19734 23910 19780 23962
rect 19484 23908 19540 23910
rect 19564 23908 19620 23910
rect 19644 23908 19700 23910
rect 19724 23908 19780 23910
rect 19484 22874 19540 22876
rect 19564 22874 19620 22876
rect 19644 22874 19700 22876
rect 19724 22874 19780 22876
rect 19484 22822 19530 22874
rect 19530 22822 19540 22874
rect 19564 22822 19594 22874
rect 19594 22822 19606 22874
rect 19606 22822 19620 22874
rect 19644 22822 19658 22874
rect 19658 22822 19670 22874
rect 19670 22822 19700 22874
rect 19724 22822 19734 22874
rect 19734 22822 19780 22874
rect 19484 22820 19540 22822
rect 19564 22820 19620 22822
rect 19644 22820 19700 22822
rect 19724 22820 19780 22822
rect 19484 21786 19540 21788
rect 19564 21786 19620 21788
rect 19644 21786 19700 21788
rect 19724 21786 19780 21788
rect 19484 21734 19530 21786
rect 19530 21734 19540 21786
rect 19564 21734 19594 21786
rect 19594 21734 19606 21786
rect 19606 21734 19620 21786
rect 19644 21734 19658 21786
rect 19658 21734 19670 21786
rect 19670 21734 19700 21786
rect 19724 21734 19734 21786
rect 19734 21734 19780 21786
rect 19484 21732 19540 21734
rect 19564 21732 19620 21734
rect 19644 21732 19700 21734
rect 19724 21732 19780 21734
rect 19484 20698 19540 20700
rect 19564 20698 19620 20700
rect 19644 20698 19700 20700
rect 19724 20698 19780 20700
rect 19484 20646 19530 20698
rect 19530 20646 19540 20698
rect 19564 20646 19594 20698
rect 19594 20646 19606 20698
rect 19606 20646 19620 20698
rect 19644 20646 19658 20698
rect 19658 20646 19670 20698
rect 19670 20646 19700 20698
rect 19724 20646 19734 20698
rect 19734 20646 19780 20698
rect 19484 20644 19540 20646
rect 19564 20644 19620 20646
rect 19644 20644 19700 20646
rect 19724 20644 19780 20646
rect 19484 19610 19540 19612
rect 19564 19610 19620 19612
rect 19644 19610 19700 19612
rect 19724 19610 19780 19612
rect 19484 19558 19530 19610
rect 19530 19558 19540 19610
rect 19564 19558 19594 19610
rect 19594 19558 19606 19610
rect 19606 19558 19620 19610
rect 19644 19558 19658 19610
rect 19658 19558 19670 19610
rect 19670 19558 19700 19610
rect 19724 19558 19734 19610
rect 19734 19558 19780 19610
rect 19484 19556 19540 19558
rect 19564 19556 19620 19558
rect 19644 19556 19700 19558
rect 19724 19556 19780 19558
rect 21822 33940 21824 33960
rect 21824 33940 21876 33960
rect 21876 33940 21878 33960
rect 21822 33904 21878 33940
rect 24116 45178 24172 45180
rect 24196 45178 24252 45180
rect 24276 45178 24332 45180
rect 24356 45178 24412 45180
rect 24116 45126 24162 45178
rect 24162 45126 24172 45178
rect 24196 45126 24226 45178
rect 24226 45126 24238 45178
rect 24238 45126 24252 45178
rect 24276 45126 24290 45178
rect 24290 45126 24302 45178
rect 24302 45126 24332 45178
rect 24356 45126 24366 45178
rect 24366 45126 24412 45178
rect 24116 45124 24172 45126
rect 24196 45124 24252 45126
rect 24276 45124 24332 45126
rect 24356 45124 24412 45126
rect 24116 44090 24172 44092
rect 24196 44090 24252 44092
rect 24276 44090 24332 44092
rect 24356 44090 24412 44092
rect 24116 44038 24162 44090
rect 24162 44038 24172 44090
rect 24196 44038 24226 44090
rect 24226 44038 24238 44090
rect 24238 44038 24252 44090
rect 24276 44038 24290 44090
rect 24290 44038 24302 44090
rect 24302 44038 24332 44090
rect 24356 44038 24366 44090
rect 24366 44038 24412 44090
rect 24116 44036 24172 44038
rect 24196 44036 24252 44038
rect 24276 44036 24332 44038
rect 24356 44036 24412 44038
rect 24116 43002 24172 43004
rect 24196 43002 24252 43004
rect 24276 43002 24332 43004
rect 24356 43002 24412 43004
rect 24116 42950 24162 43002
rect 24162 42950 24172 43002
rect 24196 42950 24226 43002
rect 24226 42950 24238 43002
rect 24238 42950 24252 43002
rect 24276 42950 24290 43002
rect 24290 42950 24302 43002
rect 24302 42950 24332 43002
rect 24356 42950 24366 43002
rect 24366 42950 24412 43002
rect 24116 42948 24172 42950
rect 24196 42948 24252 42950
rect 24276 42948 24332 42950
rect 24356 42948 24412 42950
rect 26054 42200 26110 42256
rect 24116 41914 24172 41916
rect 24196 41914 24252 41916
rect 24276 41914 24332 41916
rect 24356 41914 24412 41916
rect 24116 41862 24162 41914
rect 24162 41862 24172 41914
rect 24196 41862 24226 41914
rect 24226 41862 24238 41914
rect 24238 41862 24252 41914
rect 24276 41862 24290 41914
rect 24290 41862 24302 41914
rect 24302 41862 24332 41914
rect 24356 41862 24366 41914
rect 24366 41862 24412 41914
rect 24116 41860 24172 41862
rect 24196 41860 24252 41862
rect 24276 41860 24332 41862
rect 24356 41860 24412 41862
rect 25962 41520 26018 41576
rect 24116 40826 24172 40828
rect 24196 40826 24252 40828
rect 24276 40826 24332 40828
rect 24356 40826 24412 40828
rect 24116 40774 24162 40826
rect 24162 40774 24172 40826
rect 24196 40774 24226 40826
rect 24226 40774 24238 40826
rect 24238 40774 24252 40826
rect 24276 40774 24290 40826
rect 24290 40774 24302 40826
rect 24302 40774 24332 40826
rect 24356 40774 24366 40826
rect 24366 40774 24412 40826
rect 24116 40772 24172 40774
rect 24196 40772 24252 40774
rect 24276 40772 24332 40774
rect 24356 40772 24412 40774
rect 24116 39738 24172 39740
rect 24196 39738 24252 39740
rect 24276 39738 24332 39740
rect 24356 39738 24412 39740
rect 24116 39686 24162 39738
rect 24162 39686 24172 39738
rect 24196 39686 24226 39738
rect 24226 39686 24238 39738
rect 24238 39686 24252 39738
rect 24276 39686 24290 39738
rect 24290 39686 24302 39738
rect 24302 39686 24332 39738
rect 24356 39686 24366 39738
rect 24366 39686 24412 39738
rect 24116 39684 24172 39686
rect 24196 39684 24252 39686
rect 24276 39684 24332 39686
rect 24356 39684 24412 39686
rect 24116 38650 24172 38652
rect 24196 38650 24252 38652
rect 24276 38650 24332 38652
rect 24356 38650 24412 38652
rect 24116 38598 24162 38650
rect 24162 38598 24172 38650
rect 24196 38598 24226 38650
rect 24226 38598 24238 38650
rect 24238 38598 24252 38650
rect 24276 38598 24290 38650
rect 24290 38598 24302 38650
rect 24302 38598 24332 38650
rect 24356 38598 24366 38650
rect 24366 38598 24412 38650
rect 24116 38596 24172 38598
rect 24196 38596 24252 38598
rect 24276 38596 24332 38598
rect 24356 38596 24412 38598
rect 24116 37562 24172 37564
rect 24196 37562 24252 37564
rect 24276 37562 24332 37564
rect 24356 37562 24412 37564
rect 24116 37510 24162 37562
rect 24162 37510 24172 37562
rect 24196 37510 24226 37562
rect 24226 37510 24238 37562
rect 24238 37510 24252 37562
rect 24276 37510 24290 37562
rect 24290 37510 24302 37562
rect 24302 37510 24332 37562
rect 24356 37510 24366 37562
rect 24366 37510 24412 37562
rect 24116 37508 24172 37510
rect 24196 37508 24252 37510
rect 24276 37508 24332 37510
rect 24356 37508 24412 37510
rect 24116 36474 24172 36476
rect 24196 36474 24252 36476
rect 24276 36474 24332 36476
rect 24356 36474 24412 36476
rect 24116 36422 24162 36474
rect 24162 36422 24172 36474
rect 24196 36422 24226 36474
rect 24226 36422 24238 36474
rect 24238 36422 24252 36474
rect 24276 36422 24290 36474
rect 24290 36422 24302 36474
rect 24302 36422 24332 36474
rect 24356 36422 24366 36474
rect 24366 36422 24412 36474
rect 24116 36420 24172 36422
rect 24196 36420 24252 36422
rect 24276 36420 24332 36422
rect 24356 36420 24412 36422
rect 22374 32272 22430 32328
rect 24116 35386 24172 35388
rect 24196 35386 24252 35388
rect 24276 35386 24332 35388
rect 24356 35386 24412 35388
rect 24116 35334 24162 35386
rect 24162 35334 24172 35386
rect 24196 35334 24226 35386
rect 24226 35334 24238 35386
rect 24238 35334 24252 35386
rect 24276 35334 24290 35386
rect 24290 35334 24302 35386
rect 24302 35334 24332 35386
rect 24356 35334 24366 35386
rect 24366 35334 24412 35386
rect 24116 35332 24172 35334
rect 24196 35332 24252 35334
rect 24276 35332 24332 35334
rect 24356 35332 24412 35334
rect 19484 18522 19540 18524
rect 19564 18522 19620 18524
rect 19644 18522 19700 18524
rect 19724 18522 19780 18524
rect 19484 18470 19530 18522
rect 19530 18470 19540 18522
rect 19564 18470 19594 18522
rect 19594 18470 19606 18522
rect 19606 18470 19620 18522
rect 19644 18470 19658 18522
rect 19658 18470 19670 18522
rect 19670 18470 19700 18522
rect 19724 18470 19734 18522
rect 19734 18470 19780 18522
rect 19484 18468 19540 18470
rect 19564 18468 19620 18470
rect 19644 18468 19700 18470
rect 19724 18468 19780 18470
rect 19484 17434 19540 17436
rect 19564 17434 19620 17436
rect 19644 17434 19700 17436
rect 19724 17434 19780 17436
rect 19484 17382 19530 17434
rect 19530 17382 19540 17434
rect 19564 17382 19594 17434
rect 19594 17382 19606 17434
rect 19606 17382 19620 17434
rect 19644 17382 19658 17434
rect 19658 17382 19670 17434
rect 19670 17382 19700 17434
rect 19724 17382 19734 17434
rect 19734 17382 19780 17434
rect 19484 17380 19540 17382
rect 19564 17380 19620 17382
rect 19644 17380 19700 17382
rect 19724 17380 19780 17382
rect 19484 16346 19540 16348
rect 19564 16346 19620 16348
rect 19644 16346 19700 16348
rect 19724 16346 19780 16348
rect 19484 16294 19530 16346
rect 19530 16294 19540 16346
rect 19564 16294 19594 16346
rect 19594 16294 19606 16346
rect 19606 16294 19620 16346
rect 19644 16294 19658 16346
rect 19658 16294 19670 16346
rect 19670 16294 19700 16346
rect 19724 16294 19734 16346
rect 19734 16294 19780 16346
rect 19484 16292 19540 16294
rect 19564 16292 19620 16294
rect 19644 16292 19700 16294
rect 19724 16292 19780 16294
rect 19484 15258 19540 15260
rect 19564 15258 19620 15260
rect 19644 15258 19700 15260
rect 19724 15258 19780 15260
rect 19484 15206 19530 15258
rect 19530 15206 19540 15258
rect 19564 15206 19594 15258
rect 19594 15206 19606 15258
rect 19606 15206 19620 15258
rect 19644 15206 19658 15258
rect 19658 15206 19670 15258
rect 19670 15206 19700 15258
rect 19724 15206 19734 15258
rect 19734 15206 19780 15258
rect 19484 15204 19540 15206
rect 19564 15204 19620 15206
rect 19644 15204 19700 15206
rect 19724 15204 19780 15206
rect 19484 14170 19540 14172
rect 19564 14170 19620 14172
rect 19644 14170 19700 14172
rect 19724 14170 19780 14172
rect 19484 14118 19530 14170
rect 19530 14118 19540 14170
rect 19564 14118 19594 14170
rect 19594 14118 19606 14170
rect 19606 14118 19620 14170
rect 19644 14118 19658 14170
rect 19658 14118 19670 14170
rect 19670 14118 19700 14170
rect 19724 14118 19734 14170
rect 19734 14118 19780 14170
rect 19484 14116 19540 14118
rect 19564 14116 19620 14118
rect 19644 14116 19700 14118
rect 19724 14116 19780 14118
rect 19484 13082 19540 13084
rect 19564 13082 19620 13084
rect 19644 13082 19700 13084
rect 19724 13082 19780 13084
rect 19484 13030 19530 13082
rect 19530 13030 19540 13082
rect 19564 13030 19594 13082
rect 19594 13030 19606 13082
rect 19606 13030 19620 13082
rect 19644 13030 19658 13082
rect 19658 13030 19670 13082
rect 19670 13030 19700 13082
rect 19724 13030 19734 13082
rect 19734 13030 19780 13082
rect 19484 13028 19540 13030
rect 19564 13028 19620 13030
rect 19644 13028 19700 13030
rect 19724 13028 19780 13030
rect 19484 11994 19540 11996
rect 19564 11994 19620 11996
rect 19644 11994 19700 11996
rect 19724 11994 19780 11996
rect 19484 11942 19530 11994
rect 19530 11942 19540 11994
rect 19564 11942 19594 11994
rect 19594 11942 19606 11994
rect 19606 11942 19620 11994
rect 19644 11942 19658 11994
rect 19658 11942 19670 11994
rect 19670 11942 19700 11994
rect 19724 11942 19734 11994
rect 19734 11942 19780 11994
rect 19484 11940 19540 11942
rect 19564 11940 19620 11942
rect 19644 11940 19700 11942
rect 19724 11940 19780 11942
rect 22006 23432 22062 23488
rect 22006 21548 22062 21584
rect 22006 21528 22008 21548
rect 22008 21528 22060 21548
rect 22060 21528 22062 21548
rect 24116 34298 24172 34300
rect 24196 34298 24252 34300
rect 24276 34298 24332 34300
rect 24356 34298 24412 34300
rect 24116 34246 24162 34298
rect 24162 34246 24172 34298
rect 24196 34246 24226 34298
rect 24226 34246 24238 34298
rect 24238 34246 24252 34298
rect 24276 34246 24290 34298
rect 24290 34246 24302 34298
rect 24302 34246 24332 34298
rect 24356 34246 24366 34298
rect 24366 34246 24412 34298
rect 24116 34244 24172 34246
rect 24196 34244 24252 34246
rect 24276 34244 24332 34246
rect 24356 34244 24412 34246
rect 24116 33210 24172 33212
rect 24196 33210 24252 33212
rect 24276 33210 24332 33212
rect 24356 33210 24412 33212
rect 24116 33158 24162 33210
rect 24162 33158 24172 33210
rect 24196 33158 24226 33210
rect 24226 33158 24238 33210
rect 24238 33158 24252 33210
rect 24276 33158 24290 33210
rect 24290 33158 24302 33210
rect 24302 33158 24332 33210
rect 24356 33158 24366 33210
rect 24366 33158 24412 33210
rect 24116 33156 24172 33158
rect 24196 33156 24252 33158
rect 24276 33156 24332 33158
rect 24356 33156 24412 33158
rect 24116 32122 24172 32124
rect 24196 32122 24252 32124
rect 24276 32122 24332 32124
rect 24356 32122 24412 32124
rect 24116 32070 24162 32122
rect 24162 32070 24172 32122
rect 24196 32070 24226 32122
rect 24226 32070 24238 32122
rect 24238 32070 24252 32122
rect 24276 32070 24290 32122
rect 24290 32070 24302 32122
rect 24302 32070 24332 32122
rect 24356 32070 24366 32122
rect 24366 32070 24412 32122
rect 24116 32068 24172 32070
rect 24196 32068 24252 32070
rect 24276 32068 24332 32070
rect 24356 32068 24412 32070
rect 24116 31034 24172 31036
rect 24196 31034 24252 31036
rect 24276 31034 24332 31036
rect 24356 31034 24412 31036
rect 24116 30982 24162 31034
rect 24162 30982 24172 31034
rect 24196 30982 24226 31034
rect 24226 30982 24238 31034
rect 24238 30982 24252 31034
rect 24276 30982 24290 31034
rect 24290 30982 24302 31034
rect 24302 30982 24332 31034
rect 24356 30982 24366 31034
rect 24366 30982 24412 31034
rect 24116 30980 24172 30982
rect 24196 30980 24252 30982
rect 24276 30980 24332 30982
rect 24356 30980 24412 30982
rect 24116 29946 24172 29948
rect 24196 29946 24252 29948
rect 24276 29946 24332 29948
rect 24356 29946 24412 29948
rect 24116 29894 24162 29946
rect 24162 29894 24172 29946
rect 24196 29894 24226 29946
rect 24226 29894 24238 29946
rect 24238 29894 24252 29946
rect 24276 29894 24290 29946
rect 24290 29894 24302 29946
rect 24302 29894 24332 29946
rect 24356 29894 24366 29946
rect 24366 29894 24412 29946
rect 24116 29892 24172 29894
rect 24196 29892 24252 29894
rect 24276 29892 24332 29894
rect 24356 29892 24412 29894
rect 24116 28858 24172 28860
rect 24196 28858 24252 28860
rect 24276 28858 24332 28860
rect 24356 28858 24412 28860
rect 24116 28806 24162 28858
rect 24162 28806 24172 28858
rect 24196 28806 24226 28858
rect 24226 28806 24238 28858
rect 24238 28806 24252 28858
rect 24276 28806 24290 28858
rect 24290 28806 24302 28858
rect 24302 28806 24332 28858
rect 24356 28806 24366 28858
rect 24366 28806 24412 28858
rect 24116 28804 24172 28806
rect 24196 28804 24252 28806
rect 24276 28804 24332 28806
rect 24356 28804 24412 28806
rect 24116 27770 24172 27772
rect 24196 27770 24252 27772
rect 24276 27770 24332 27772
rect 24356 27770 24412 27772
rect 24116 27718 24162 27770
rect 24162 27718 24172 27770
rect 24196 27718 24226 27770
rect 24226 27718 24238 27770
rect 24238 27718 24252 27770
rect 24276 27718 24290 27770
rect 24290 27718 24302 27770
rect 24302 27718 24332 27770
rect 24356 27718 24366 27770
rect 24366 27718 24412 27770
rect 24116 27716 24172 27718
rect 24196 27716 24252 27718
rect 24276 27716 24332 27718
rect 24356 27716 24412 27718
rect 24116 26682 24172 26684
rect 24196 26682 24252 26684
rect 24276 26682 24332 26684
rect 24356 26682 24412 26684
rect 24116 26630 24162 26682
rect 24162 26630 24172 26682
rect 24196 26630 24226 26682
rect 24226 26630 24238 26682
rect 24238 26630 24252 26682
rect 24276 26630 24290 26682
rect 24290 26630 24302 26682
rect 24302 26630 24332 26682
rect 24356 26630 24366 26682
rect 24366 26630 24412 26682
rect 24116 26628 24172 26630
rect 24196 26628 24252 26630
rect 24276 26628 24332 26630
rect 24356 26628 24412 26630
rect 24116 25594 24172 25596
rect 24196 25594 24252 25596
rect 24276 25594 24332 25596
rect 24356 25594 24412 25596
rect 24116 25542 24162 25594
rect 24162 25542 24172 25594
rect 24196 25542 24226 25594
rect 24226 25542 24238 25594
rect 24238 25542 24252 25594
rect 24276 25542 24290 25594
rect 24290 25542 24302 25594
rect 24302 25542 24332 25594
rect 24356 25542 24366 25594
rect 24366 25542 24412 25594
rect 24116 25540 24172 25542
rect 24196 25540 24252 25542
rect 24276 25540 24332 25542
rect 24356 25540 24412 25542
rect 19484 10906 19540 10908
rect 19564 10906 19620 10908
rect 19644 10906 19700 10908
rect 19724 10906 19780 10908
rect 19484 10854 19530 10906
rect 19530 10854 19540 10906
rect 19564 10854 19594 10906
rect 19594 10854 19606 10906
rect 19606 10854 19620 10906
rect 19644 10854 19658 10906
rect 19658 10854 19670 10906
rect 19670 10854 19700 10906
rect 19724 10854 19734 10906
rect 19734 10854 19780 10906
rect 19484 10852 19540 10854
rect 19564 10852 19620 10854
rect 19644 10852 19700 10854
rect 19724 10852 19780 10854
rect 24116 24506 24172 24508
rect 24196 24506 24252 24508
rect 24276 24506 24332 24508
rect 24356 24506 24412 24508
rect 24116 24454 24162 24506
rect 24162 24454 24172 24506
rect 24196 24454 24226 24506
rect 24226 24454 24238 24506
rect 24238 24454 24252 24506
rect 24276 24454 24290 24506
rect 24290 24454 24302 24506
rect 24302 24454 24332 24506
rect 24356 24454 24366 24506
rect 24366 24454 24412 24506
rect 24116 24452 24172 24454
rect 24196 24452 24252 24454
rect 24276 24452 24332 24454
rect 24356 24452 24412 24454
rect 24116 23418 24172 23420
rect 24196 23418 24252 23420
rect 24276 23418 24332 23420
rect 24356 23418 24412 23420
rect 24116 23366 24162 23418
rect 24162 23366 24172 23418
rect 24196 23366 24226 23418
rect 24226 23366 24238 23418
rect 24238 23366 24252 23418
rect 24276 23366 24290 23418
rect 24290 23366 24302 23418
rect 24302 23366 24332 23418
rect 24356 23366 24366 23418
rect 24366 23366 24412 23418
rect 24116 23364 24172 23366
rect 24196 23364 24252 23366
rect 24276 23364 24332 23366
rect 24356 23364 24412 23366
rect 25042 29280 25098 29336
rect 25042 24132 25098 24168
rect 25042 24112 25044 24132
rect 25044 24112 25096 24132
rect 25096 24112 25098 24132
rect 24116 22330 24172 22332
rect 24196 22330 24252 22332
rect 24276 22330 24332 22332
rect 24356 22330 24412 22332
rect 24116 22278 24162 22330
rect 24162 22278 24172 22330
rect 24196 22278 24226 22330
rect 24226 22278 24238 22330
rect 24238 22278 24252 22330
rect 24276 22278 24290 22330
rect 24290 22278 24302 22330
rect 24302 22278 24332 22330
rect 24356 22278 24366 22330
rect 24366 22278 24412 22330
rect 24116 22276 24172 22278
rect 24196 22276 24252 22278
rect 24276 22276 24332 22278
rect 24356 22276 24412 22278
rect 24116 21242 24172 21244
rect 24196 21242 24252 21244
rect 24276 21242 24332 21244
rect 24356 21242 24412 21244
rect 24116 21190 24162 21242
rect 24162 21190 24172 21242
rect 24196 21190 24226 21242
rect 24226 21190 24238 21242
rect 24238 21190 24252 21242
rect 24276 21190 24290 21242
rect 24290 21190 24302 21242
rect 24302 21190 24332 21242
rect 24356 21190 24366 21242
rect 24366 21190 24412 21242
rect 24116 21188 24172 21190
rect 24196 21188 24252 21190
rect 24276 21188 24332 21190
rect 24356 21188 24412 21190
rect 24116 20154 24172 20156
rect 24196 20154 24252 20156
rect 24276 20154 24332 20156
rect 24356 20154 24412 20156
rect 24116 20102 24162 20154
rect 24162 20102 24172 20154
rect 24196 20102 24226 20154
rect 24226 20102 24238 20154
rect 24238 20102 24252 20154
rect 24276 20102 24290 20154
rect 24290 20102 24302 20154
rect 24302 20102 24332 20154
rect 24356 20102 24366 20154
rect 24366 20102 24412 20154
rect 24116 20100 24172 20102
rect 24196 20100 24252 20102
rect 24276 20100 24332 20102
rect 24356 20100 24412 20102
rect 24116 19066 24172 19068
rect 24196 19066 24252 19068
rect 24276 19066 24332 19068
rect 24356 19066 24412 19068
rect 24116 19014 24162 19066
rect 24162 19014 24172 19066
rect 24196 19014 24226 19066
rect 24226 19014 24238 19066
rect 24238 19014 24252 19066
rect 24276 19014 24290 19066
rect 24290 19014 24302 19066
rect 24302 19014 24332 19066
rect 24356 19014 24366 19066
rect 24366 19014 24412 19066
rect 24116 19012 24172 19014
rect 24196 19012 24252 19014
rect 24276 19012 24332 19014
rect 24356 19012 24412 19014
rect 24116 17978 24172 17980
rect 24196 17978 24252 17980
rect 24276 17978 24332 17980
rect 24356 17978 24412 17980
rect 24116 17926 24162 17978
rect 24162 17926 24172 17978
rect 24196 17926 24226 17978
rect 24226 17926 24238 17978
rect 24238 17926 24252 17978
rect 24276 17926 24290 17978
rect 24290 17926 24302 17978
rect 24302 17926 24332 17978
rect 24356 17926 24366 17978
rect 24366 17926 24412 17978
rect 24116 17924 24172 17926
rect 24196 17924 24252 17926
rect 24276 17924 24332 17926
rect 24356 17924 24412 17926
rect 24116 16890 24172 16892
rect 24196 16890 24252 16892
rect 24276 16890 24332 16892
rect 24356 16890 24412 16892
rect 24116 16838 24162 16890
rect 24162 16838 24172 16890
rect 24196 16838 24226 16890
rect 24226 16838 24238 16890
rect 24238 16838 24252 16890
rect 24276 16838 24290 16890
rect 24290 16838 24302 16890
rect 24302 16838 24332 16890
rect 24356 16838 24366 16890
rect 24366 16838 24412 16890
rect 24116 16836 24172 16838
rect 24196 16836 24252 16838
rect 24276 16836 24332 16838
rect 24356 16836 24412 16838
rect 24116 15802 24172 15804
rect 24196 15802 24252 15804
rect 24276 15802 24332 15804
rect 24356 15802 24412 15804
rect 24116 15750 24162 15802
rect 24162 15750 24172 15802
rect 24196 15750 24226 15802
rect 24226 15750 24238 15802
rect 24238 15750 24252 15802
rect 24276 15750 24290 15802
rect 24290 15750 24302 15802
rect 24302 15750 24332 15802
rect 24356 15750 24366 15802
rect 24366 15750 24412 15802
rect 24116 15748 24172 15750
rect 24196 15748 24252 15750
rect 24276 15748 24332 15750
rect 24356 15748 24412 15750
rect 24116 14714 24172 14716
rect 24196 14714 24252 14716
rect 24276 14714 24332 14716
rect 24356 14714 24412 14716
rect 24116 14662 24162 14714
rect 24162 14662 24172 14714
rect 24196 14662 24226 14714
rect 24226 14662 24238 14714
rect 24238 14662 24252 14714
rect 24276 14662 24290 14714
rect 24290 14662 24302 14714
rect 24302 14662 24332 14714
rect 24356 14662 24366 14714
rect 24366 14662 24412 14714
rect 24116 14660 24172 14662
rect 24196 14660 24252 14662
rect 24276 14660 24332 14662
rect 24356 14660 24412 14662
rect 24116 13626 24172 13628
rect 24196 13626 24252 13628
rect 24276 13626 24332 13628
rect 24356 13626 24412 13628
rect 24116 13574 24162 13626
rect 24162 13574 24172 13626
rect 24196 13574 24226 13626
rect 24226 13574 24238 13626
rect 24238 13574 24252 13626
rect 24276 13574 24290 13626
rect 24290 13574 24302 13626
rect 24302 13574 24332 13626
rect 24356 13574 24366 13626
rect 24366 13574 24412 13626
rect 24116 13572 24172 13574
rect 24196 13572 24252 13574
rect 24276 13572 24332 13574
rect 24356 13572 24412 13574
rect 24858 15000 24914 15056
rect 24116 12538 24172 12540
rect 24196 12538 24252 12540
rect 24276 12538 24332 12540
rect 24356 12538 24412 12540
rect 24116 12486 24162 12538
rect 24162 12486 24172 12538
rect 24196 12486 24226 12538
rect 24226 12486 24238 12538
rect 24238 12486 24252 12538
rect 24276 12486 24290 12538
rect 24290 12486 24302 12538
rect 24302 12486 24332 12538
rect 24356 12486 24366 12538
rect 24366 12486 24412 12538
rect 24116 12484 24172 12486
rect 24196 12484 24252 12486
rect 24276 12484 24332 12486
rect 24356 12484 24412 12486
rect 25778 26560 25834 26616
rect 25226 15544 25282 15600
rect 25962 32680 26018 32736
rect 25962 24520 26018 24576
rect 26790 36760 26846 36816
rect 27526 44940 27582 44976
rect 27526 44920 27528 44940
rect 27528 44920 27580 44940
rect 27580 44920 27582 44940
rect 26146 21120 26202 21176
rect 27526 40840 27582 40896
rect 27526 36080 27582 36136
rect 27434 34620 27436 34640
rect 27436 34620 27488 34640
rect 27488 34620 27490 34640
rect 27434 34584 27490 34620
rect 27526 34060 27582 34096
rect 27526 34040 27528 34060
rect 27528 34040 27580 34060
rect 27580 34040 27582 34060
rect 27342 29960 27398 30016
rect 28814 46960 28870 47016
rect 28170 42880 28226 42936
rect 28170 40160 28226 40216
rect 28722 39480 28778 39536
rect 27526 30640 27582 30696
rect 27526 28620 27582 28656
rect 27526 28600 27528 28620
rect 27528 28600 27580 28620
rect 27580 28600 27582 28620
rect 27526 27240 27582 27296
rect 24116 11450 24172 11452
rect 24196 11450 24252 11452
rect 24276 11450 24332 11452
rect 24356 11450 24412 11452
rect 24116 11398 24162 11450
rect 24162 11398 24172 11450
rect 24196 11398 24226 11450
rect 24226 11398 24238 11450
rect 24238 11398 24252 11450
rect 24276 11398 24290 11450
rect 24290 11398 24302 11450
rect 24302 11398 24332 11450
rect 24356 11398 24366 11450
rect 24366 11398 24412 11450
rect 24116 11396 24172 11398
rect 24196 11396 24252 11398
rect 24276 11396 24332 11398
rect 24356 11396 24412 11398
rect 19484 9818 19540 9820
rect 19564 9818 19620 9820
rect 19644 9818 19700 9820
rect 19724 9818 19780 9820
rect 19484 9766 19530 9818
rect 19530 9766 19540 9818
rect 19564 9766 19594 9818
rect 19594 9766 19606 9818
rect 19606 9766 19620 9818
rect 19644 9766 19658 9818
rect 19658 9766 19670 9818
rect 19670 9766 19700 9818
rect 19724 9766 19734 9818
rect 19734 9766 19780 9818
rect 19484 9764 19540 9766
rect 19564 9764 19620 9766
rect 19644 9764 19700 9766
rect 19724 9764 19780 9766
rect 19484 8730 19540 8732
rect 19564 8730 19620 8732
rect 19644 8730 19700 8732
rect 19724 8730 19780 8732
rect 19484 8678 19530 8730
rect 19530 8678 19540 8730
rect 19564 8678 19594 8730
rect 19594 8678 19606 8730
rect 19606 8678 19620 8730
rect 19644 8678 19658 8730
rect 19658 8678 19670 8730
rect 19670 8678 19700 8730
rect 19724 8678 19734 8730
rect 19734 8678 19780 8730
rect 19484 8676 19540 8678
rect 19564 8676 19620 8678
rect 19644 8676 19700 8678
rect 19724 8676 19780 8678
rect 18694 7928 18750 7984
rect 19484 7642 19540 7644
rect 19564 7642 19620 7644
rect 19644 7642 19700 7644
rect 19724 7642 19780 7644
rect 19484 7590 19530 7642
rect 19530 7590 19540 7642
rect 19564 7590 19594 7642
rect 19594 7590 19606 7642
rect 19606 7590 19620 7642
rect 19644 7590 19658 7642
rect 19658 7590 19670 7642
rect 19670 7590 19700 7642
rect 19724 7590 19734 7642
rect 19734 7590 19780 7642
rect 19484 7588 19540 7590
rect 19564 7588 19620 7590
rect 19644 7588 19700 7590
rect 19724 7588 19780 7590
rect 19484 6554 19540 6556
rect 19564 6554 19620 6556
rect 19644 6554 19700 6556
rect 19724 6554 19780 6556
rect 19484 6502 19530 6554
rect 19530 6502 19540 6554
rect 19564 6502 19594 6554
rect 19594 6502 19606 6554
rect 19606 6502 19620 6554
rect 19644 6502 19658 6554
rect 19658 6502 19670 6554
rect 19670 6502 19700 6554
rect 19724 6502 19734 6554
rect 19734 6502 19780 6554
rect 19484 6500 19540 6502
rect 19564 6500 19620 6502
rect 19644 6500 19700 6502
rect 19724 6500 19780 6502
rect 19484 5466 19540 5468
rect 19564 5466 19620 5468
rect 19644 5466 19700 5468
rect 19724 5466 19780 5468
rect 19484 5414 19530 5466
rect 19530 5414 19540 5466
rect 19564 5414 19594 5466
rect 19594 5414 19606 5466
rect 19606 5414 19620 5466
rect 19644 5414 19658 5466
rect 19658 5414 19670 5466
rect 19670 5414 19700 5466
rect 19724 5414 19734 5466
rect 19734 5414 19780 5466
rect 19484 5412 19540 5414
rect 19564 5412 19620 5414
rect 19644 5412 19700 5414
rect 19724 5412 19780 5414
rect 19484 4378 19540 4380
rect 19564 4378 19620 4380
rect 19644 4378 19700 4380
rect 19724 4378 19780 4380
rect 19484 4326 19530 4378
rect 19530 4326 19540 4378
rect 19564 4326 19594 4378
rect 19594 4326 19606 4378
rect 19606 4326 19620 4378
rect 19644 4326 19658 4378
rect 19658 4326 19670 4378
rect 19670 4326 19700 4378
rect 19724 4326 19734 4378
rect 19734 4326 19780 4378
rect 19484 4324 19540 4326
rect 19564 4324 19620 4326
rect 19644 4324 19700 4326
rect 19724 4324 19780 4326
rect 19484 3290 19540 3292
rect 19564 3290 19620 3292
rect 19644 3290 19700 3292
rect 19724 3290 19780 3292
rect 19484 3238 19530 3290
rect 19530 3238 19540 3290
rect 19564 3238 19594 3290
rect 19594 3238 19606 3290
rect 19606 3238 19620 3290
rect 19644 3238 19658 3290
rect 19658 3238 19670 3290
rect 19670 3238 19700 3290
rect 19724 3238 19734 3290
rect 19734 3238 19780 3290
rect 19484 3236 19540 3238
rect 19564 3236 19620 3238
rect 19644 3236 19700 3238
rect 19724 3236 19780 3238
rect 19484 2202 19540 2204
rect 19564 2202 19620 2204
rect 19644 2202 19700 2204
rect 19724 2202 19780 2204
rect 19484 2150 19530 2202
rect 19530 2150 19540 2202
rect 19564 2150 19594 2202
rect 19594 2150 19606 2202
rect 19606 2150 19620 2202
rect 19644 2150 19658 2202
rect 19658 2150 19670 2202
rect 19670 2150 19700 2202
rect 19724 2150 19734 2202
rect 19734 2150 19780 2202
rect 19484 2148 19540 2150
rect 19564 2148 19620 2150
rect 19644 2148 19700 2150
rect 19724 2148 19780 2150
rect 24116 10362 24172 10364
rect 24196 10362 24252 10364
rect 24276 10362 24332 10364
rect 24356 10362 24412 10364
rect 24116 10310 24162 10362
rect 24162 10310 24172 10362
rect 24196 10310 24226 10362
rect 24226 10310 24238 10362
rect 24238 10310 24252 10362
rect 24276 10310 24290 10362
rect 24290 10310 24302 10362
rect 24302 10310 24332 10362
rect 24356 10310 24366 10362
rect 24366 10310 24412 10362
rect 24116 10308 24172 10310
rect 24196 10308 24252 10310
rect 24276 10308 24332 10310
rect 24356 10308 24412 10310
rect 24116 9274 24172 9276
rect 24196 9274 24252 9276
rect 24276 9274 24332 9276
rect 24356 9274 24412 9276
rect 24116 9222 24162 9274
rect 24162 9222 24172 9274
rect 24196 9222 24226 9274
rect 24226 9222 24238 9274
rect 24238 9222 24252 9274
rect 24276 9222 24290 9274
rect 24290 9222 24302 9274
rect 24302 9222 24332 9274
rect 24356 9222 24366 9274
rect 24366 9222 24412 9274
rect 24116 9220 24172 9222
rect 24196 9220 24252 9222
rect 24276 9220 24332 9222
rect 24356 9220 24412 9222
rect 24116 8186 24172 8188
rect 24196 8186 24252 8188
rect 24276 8186 24332 8188
rect 24356 8186 24412 8188
rect 24116 8134 24162 8186
rect 24162 8134 24172 8186
rect 24196 8134 24226 8186
rect 24226 8134 24238 8186
rect 24238 8134 24252 8186
rect 24276 8134 24290 8186
rect 24290 8134 24302 8186
rect 24302 8134 24332 8186
rect 24356 8134 24366 8186
rect 24366 8134 24412 8186
rect 24116 8132 24172 8134
rect 24196 8132 24252 8134
rect 24276 8132 24332 8134
rect 24356 8132 24412 8134
rect 24116 7098 24172 7100
rect 24196 7098 24252 7100
rect 24276 7098 24332 7100
rect 24356 7098 24412 7100
rect 24116 7046 24162 7098
rect 24162 7046 24172 7098
rect 24196 7046 24226 7098
rect 24226 7046 24238 7098
rect 24238 7046 24252 7098
rect 24276 7046 24290 7098
rect 24290 7046 24302 7098
rect 24302 7046 24332 7098
rect 24356 7046 24366 7098
rect 24366 7046 24412 7098
rect 24116 7044 24172 7046
rect 24196 7044 24252 7046
rect 24276 7044 24332 7046
rect 24356 7044 24412 7046
rect 25962 10240 26018 10296
rect 24116 6010 24172 6012
rect 24196 6010 24252 6012
rect 24276 6010 24332 6012
rect 24356 6010 24412 6012
rect 24116 5958 24162 6010
rect 24162 5958 24172 6010
rect 24196 5958 24226 6010
rect 24226 5958 24238 6010
rect 24238 5958 24252 6010
rect 24276 5958 24290 6010
rect 24290 5958 24302 6010
rect 24302 5958 24332 6010
rect 24356 5958 24366 6010
rect 24366 5958 24412 6010
rect 24116 5956 24172 5958
rect 24196 5956 24252 5958
rect 24276 5956 24332 5958
rect 24356 5956 24412 5958
rect 24116 4922 24172 4924
rect 24196 4922 24252 4924
rect 24276 4922 24332 4924
rect 24356 4922 24412 4924
rect 24116 4870 24162 4922
rect 24162 4870 24172 4922
rect 24196 4870 24226 4922
rect 24226 4870 24238 4922
rect 24238 4870 24252 4922
rect 24276 4870 24290 4922
rect 24290 4870 24302 4922
rect 24302 4870 24332 4922
rect 24356 4870 24366 4922
rect 24366 4870 24412 4922
rect 24116 4868 24172 4870
rect 24196 4868 24252 4870
rect 24276 4868 24332 4870
rect 24356 4868 24412 4870
rect 24116 3834 24172 3836
rect 24196 3834 24252 3836
rect 24276 3834 24332 3836
rect 24356 3834 24412 3836
rect 24116 3782 24162 3834
rect 24162 3782 24172 3834
rect 24196 3782 24226 3834
rect 24226 3782 24238 3834
rect 24238 3782 24252 3834
rect 24276 3782 24290 3834
rect 24290 3782 24302 3834
rect 24302 3782 24332 3834
rect 24356 3782 24366 3834
rect 24366 3782 24412 3834
rect 24116 3780 24172 3782
rect 24196 3780 24252 3782
rect 24276 3780 24332 3782
rect 24356 3780 24412 3782
rect 25042 3576 25098 3632
rect 24116 2746 24172 2748
rect 24196 2746 24252 2748
rect 24276 2746 24332 2748
rect 24356 2746 24412 2748
rect 24116 2694 24162 2746
rect 24162 2694 24172 2746
rect 24196 2694 24226 2746
rect 24226 2694 24238 2746
rect 24238 2694 24252 2746
rect 24276 2694 24290 2746
rect 24290 2694 24302 2746
rect 24302 2694 24332 2746
rect 24356 2694 24366 2746
rect 24366 2694 24412 2746
rect 24116 2692 24172 2694
rect 24196 2692 24252 2694
rect 24276 2692 24332 2694
rect 24356 2692 24412 2694
rect 26146 8880 26202 8936
rect 25962 8200 26018 8256
rect 27526 25200 27582 25256
rect 27526 23840 27582 23896
rect 27342 20304 27398 20360
rect 27342 19760 27398 19816
rect 27526 14320 27582 14376
rect 27526 12280 27582 12336
rect 27526 10920 27582 10976
rect 28170 21800 28226 21856
rect 28170 20440 28226 20496
rect 28078 16360 28134 16416
rect 28170 15680 28226 15736
rect 27802 13932 27858 13968
rect 27802 13912 27804 13932
rect 27804 13912 27856 13932
rect 27856 13912 27858 13932
rect 27526 7520 27582 7576
rect 27526 6860 27582 6896
rect 27526 6840 27528 6860
rect 27528 6840 27580 6860
rect 27580 6840 27582 6860
rect 25962 2760 26018 2816
rect 27434 3440 27490 3496
rect 28630 32000 28686 32056
rect 28170 5480 28226 5536
rect 28722 31320 28778 31376
rect 28998 2080 29054 2136
rect 27526 1400 27582 1456
<< metal3 >>
rect 0 49738 800 49828
rect 4061 49738 4127 49741
rect 0 49736 4127 49738
rect 0 49680 4066 49736
rect 4122 49680 4127 49736
rect 0 49678 4127 49680
rect 0 49588 800 49678
rect 4061 49675 4127 49678
rect 26141 49058 26207 49061
rect 29200 49058 30000 49148
rect 26141 49056 30000 49058
rect 26141 49000 26146 49056
rect 26202 49000 30000 49056
rect 26141 48998 30000 49000
rect 26141 48995 26207 48998
rect 29200 48908 30000 48998
rect 0 48228 800 48468
rect 29200 48228 30000 48468
rect 0 47548 800 47788
rect 25589 47698 25655 47701
rect 29200 47698 30000 47788
rect 25589 47696 30000 47698
rect 25589 47640 25594 47696
rect 25650 47640 30000 47696
rect 25589 47638 30000 47640
rect 25589 47635 25655 47638
rect 29200 47548 30000 47638
rect 5576 47360 5896 47361
rect 5576 47296 5584 47360
rect 5648 47296 5664 47360
rect 5728 47296 5744 47360
rect 5808 47296 5824 47360
rect 5888 47296 5896 47360
rect 5576 47295 5896 47296
rect 14840 47360 15160 47361
rect 14840 47296 14848 47360
rect 14912 47296 14928 47360
rect 14992 47296 15008 47360
rect 15072 47296 15088 47360
rect 15152 47296 15160 47360
rect 14840 47295 15160 47296
rect 24104 47360 24424 47361
rect 24104 47296 24112 47360
rect 24176 47296 24192 47360
rect 24256 47296 24272 47360
rect 24336 47296 24352 47360
rect 24416 47296 24424 47360
rect 24104 47295 24424 47296
rect 0 46868 800 47108
rect 28809 47018 28875 47021
rect 29200 47018 30000 47108
rect 28809 47016 30000 47018
rect 28809 46960 28814 47016
rect 28870 46960 30000 47016
rect 28809 46958 30000 46960
rect 28809 46955 28875 46958
rect 29200 46868 30000 46958
rect 10208 46816 10528 46817
rect 10208 46752 10216 46816
rect 10280 46752 10296 46816
rect 10360 46752 10376 46816
rect 10440 46752 10456 46816
rect 10520 46752 10528 46816
rect 10208 46751 10528 46752
rect 19472 46816 19792 46817
rect 19472 46752 19480 46816
rect 19544 46752 19560 46816
rect 19624 46752 19640 46816
rect 19704 46752 19720 46816
rect 19784 46752 19792 46816
rect 19472 46751 19792 46752
rect 0 46188 800 46428
rect 25957 46338 26023 46341
rect 29200 46338 30000 46428
rect 25957 46336 30000 46338
rect 25957 46280 25962 46336
rect 26018 46280 30000 46336
rect 25957 46278 30000 46280
rect 25957 46275 26023 46278
rect 5576 46272 5896 46273
rect 5576 46208 5584 46272
rect 5648 46208 5664 46272
rect 5728 46208 5744 46272
rect 5808 46208 5824 46272
rect 5888 46208 5896 46272
rect 5576 46207 5896 46208
rect 14840 46272 15160 46273
rect 14840 46208 14848 46272
rect 14912 46208 14928 46272
rect 14992 46208 15008 46272
rect 15072 46208 15088 46272
rect 15152 46208 15160 46272
rect 14840 46207 15160 46208
rect 24104 46272 24424 46273
rect 24104 46208 24112 46272
rect 24176 46208 24192 46272
rect 24256 46208 24272 46272
rect 24336 46208 24352 46272
rect 24416 46208 24424 46272
rect 24104 46207 24424 46208
rect 29200 46188 30000 46278
rect 0 45508 800 45748
rect 10208 45728 10528 45729
rect 10208 45664 10216 45728
rect 10280 45664 10296 45728
rect 10360 45664 10376 45728
rect 10440 45664 10456 45728
rect 10520 45664 10528 45728
rect 10208 45663 10528 45664
rect 19472 45728 19792 45729
rect 19472 45664 19480 45728
rect 19544 45664 19560 45728
rect 19624 45664 19640 45728
rect 19704 45664 19720 45728
rect 19784 45664 19792 45728
rect 19472 45663 19792 45664
rect 29200 45508 30000 45748
rect 5576 45184 5896 45185
rect 5576 45120 5584 45184
rect 5648 45120 5664 45184
rect 5728 45120 5744 45184
rect 5808 45120 5824 45184
rect 5888 45120 5896 45184
rect 5576 45119 5896 45120
rect 14840 45184 15160 45185
rect 14840 45120 14848 45184
rect 14912 45120 14928 45184
rect 14992 45120 15008 45184
rect 15072 45120 15088 45184
rect 15152 45120 15160 45184
rect 14840 45119 15160 45120
rect 24104 45184 24424 45185
rect 24104 45120 24112 45184
rect 24176 45120 24192 45184
rect 24256 45120 24272 45184
rect 24336 45120 24352 45184
rect 24416 45120 24424 45184
rect 24104 45119 24424 45120
rect 0 44978 800 45068
rect 3233 44978 3299 44981
rect 0 44976 3299 44978
rect 0 44920 3238 44976
rect 3294 44920 3299 44976
rect 0 44918 3299 44920
rect 0 44828 800 44918
rect 3233 44915 3299 44918
rect 27521 44978 27587 44981
rect 29200 44978 30000 45068
rect 27521 44976 30000 44978
rect 27521 44920 27526 44976
rect 27582 44920 30000 44976
rect 27521 44918 30000 44920
rect 27521 44915 27587 44918
rect 29200 44828 30000 44918
rect 10208 44640 10528 44641
rect 10208 44576 10216 44640
rect 10280 44576 10296 44640
rect 10360 44576 10376 44640
rect 10440 44576 10456 44640
rect 10520 44576 10528 44640
rect 10208 44575 10528 44576
rect 19472 44640 19792 44641
rect 19472 44576 19480 44640
rect 19544 44576 19560 44640
rect 19624 44576 19640 44640
rect 19704 44576 19720 44640
rect 19784 44576 19792 44640
rect 19472 44575 19792 44576
rect 0 44298 800 44388
rect 2865 44298 2931 44301
rect 22001 44300 22067 44301
rect 21950 44298 21956 44300
rect 0 44296 2931 44298
rect 0 44240 2870 44296
rect 2926 44240 2931 44296
rect 0 44238 2931 44240
rect 21910 44238 21956 44298
rect 22020 44296 22067 44300
rect 22062 44240 22067 44296
rect 0 44148 800 44238
rect 2865 44235 2931 44238
rect 21950 44236 21956 44238
rect 22020 44236 22067 44240
rect 22001 44235 22067 44236
rect 5576 44096 5896 44097
rect 5576 44032 5584 44096
rect 5648 44032 5664 44096
rect 5728 44032 5744 44096
rect 5808 44032 5824 44096
rect 5888 44032 5896 44096
rect 5576 44031 5896 44032
rect 14840 44096 15160 44097
rect 14840 44032 14848 44096
rect 14912 44032 14928 44096
rect 14992 44032 15008 44096
rect 15072 44032 15088 44096
rect 15152 44032 15160 44096
rect 14840 44031 15160 44032
rect 24104 44096 24424 44097
rect 24104 44032 24112 44096
rect 24176 44032 24192 44096
rect 24256 44032 24272 44096
rect 24336 44032 24352 44096
rect 24416 44032 24424 44096
rect 24104 44031 24424 44032
rect 10208 43552 10528 43553
rect 10208 43488 10216 43552
rect 10280 43488 10296 43552
rect 10360 43488 10376 43552
rect 10440 43488 10456 43552
rect 10520 43488 10528 43552
rect 10208 43487 10528 43488
rect 19472 43552 19792 43553
rect 19472 43488 19480 43552
rect 19544 43488 19560 43552
rect 19624 43488 19640 43552
rect 19704 43488 19720 43552
rect 19784 43488 19792 43552
rect 19472 43487 19792 43488
rect 29200 43468 30000 43708
rect 0 42788 800 43028
rect 5576 43008 5896 43009
rect 5576 42944 5584 43008
rect 5648 42944 5664 43008
rect 5728 42944 5744 43008
rect 5808 42944 5824 43008
rect 5888 42944 5896 43008
rect 5576 42943 5896 42944
rect 14840 43008 15160 43009
rect 14840 42944 14848 43008
rect 14912 42944 14928 43008
rect 14992 42944 15008 43008
rect 15072 42944 15088 43008
rect 15152 42944 15160 43008
rect 14840 42943 15160 42944
rect 24104 43008 24424 43009
rect 24104 42944 24112 43008
rect 24176 42944 24192 43008
rect 24256 42944 24272 43008
rect 24336 42944 24352 43008
rect 24416 42944 24424 43008
rect 24104 42943 24424 42944
rect 28165 42938 28231 42941
rect 29200 42938 30000 43028
rect 28165 42936 30000 42938
rect 28165 42880 28170 42936
rect 28226 42880 30000 42936
rect 28165 42878 30000 42880
rect 28165 42875 28231 42878
rect 29200 42788 30000 42878
rect 10208 42464 10528 42465
rect 10208 42400 10216 42464
rect 10280 42400 10296 42464
rect 10360 42400 10376 42464
rect 10440 42400 10456 42464
rect 10520 42400 10528 42464
rect 10208 42399 10528 42400
rect 19472 42464 19792 42465
rect 19472 42400 19480 42464
rect 19544 42400 19560 42464
rect 19624 42400 19640 42464
rect 19704 42400 19720 42464
rect 19784 42400 19792 42464
rect 19472 42399 19792 42400
rect 0 42258 800 42348
rect 1393 42258 1459 42261
rect 0 42256 1459 42258
rect 0 42200 1398 42256
rect 1454 42200 1459 42256
rect 0 42198 1459 42200
rect 0 42108 800 42198
rect 1393 42195 1459 42198
rect 26049 42258 26115 42261
rect 29200 42258 30000 42348
rect 26049 42256 30000 42258
rect 26049 42200 26054 42256
rect 26110 42200 30000 42256
rect 26049 42198 30000 42200
rect 26049 42195 26115 42198
rect 29200 42108 30000 42198
rect 5576 41920 5896 41921
rect 5576 41856 5584 41920
rect 5648 41856 5664 41920
rect 5728 41856 5744 41920
rect 5808 41856 5824 41920
rect 5888 41856 5896 41920
rect 5576 41855 5896 41856
rect 14840 41920 15160 41921
rect 14840 41856 14848 41920
rect 14912 41856 14928 41920
rect 14992 41856 15008 41920
rect 15072 41856 15088 41920
rect 15152 41856 15160 41920
rect 14840 41855 15160 41856
rect 24104 41920 24424 41921
rect 24104 41856 24112 41920
rect 24176 41856 24192 41920
rect 24256 41856 24272 41920
rect 24336 41856 24352 41920
rect 24416 41856 24424 41920
rect 24104 41855 24424 41856
rect 0 41578 800 41668
rect 2773 41578 2839 41581
rect 0 41576 2839 41578
rect 0 41520 2778 41576
rect 2834 41520 2839 41576
rect 0 41518 2839 41520
rect 0 41428 800 41518
rect 2773 41515 2839 41518
rect 25957 41578 26023 41581
rect 29200 41578 30000 41668
rect 25957 41576 30000 41578
rect 25957 41520 25962 41576
rect 26018 41520 30000 41576
rect 25957 41518 30000 41520
rect 25957 41515 26023 41518
rect 29200 41428 30000 41518
rect 10208 41376 10528 41377
rect 10208 41312 10216 41376
rect 10280 41312 10296 41376
rect 10360 41312 10376 41376
rect 10440 41312 10456 41376
rect 10520 41312 10528 41376
rect 10208 41311 10528 41312
rect 19472 41376 19792 41377
rect 19472 41312 19480 41376
rect 19544 41312 19560 41376
rect 19624 41312 19640 41376
rect 19704 41312 19720 41376
rect 19784 41312 19792 41376
rect 19472 41311 19792 41312
rect 0 40748 800 40988
rect 27521 40898 27587 40901
rect 29200 40898 30000 40988
rect 27521 40896 30000 40898
rect 27521 40840 27526 40896
rect 27582 40840 30000 40896
rect 27521 40838 30000 40840
rect 27521 40835 27587 40838
rect 5576 40832 5896 40833
rect 5576 40768 5584 40832
rect 5648 40768 5664 40832
rect 5728 40768 5744 40832
rect 5808 40768 5824 40832
rect 5888 40768 5896 40832
rect 5576 40767 5896 40768
rect 14840 40832 15160 40833
rect 14840 40768 14848 40832
rect 14912 40768 14928 40832
rect 14992 40768 15008 40832
rect 15072 40768 15088 40832
rect 15152 40768 15160 40832
rect 14840 40767 15160 40768
rect 24104 40832 24424 40833
rect 24104 40768 24112 40832
rect 24176 40768 24192 40832
rect 24256 40768 24272 40832
rect 24336 40768 24352 40832
rect 24416 40768 24424 40832
rect 24104 40767 24424 40768
rect 29200 40748 30000 40838
rect 0 40068 800 40308
rect 10208 40288 10528 40289
rect 10208 40224 10216 40288
rect 10280 40224 10296 40288
rect 10360 40224 10376 40288
rect 10440 40224 10456 40288
rect 10520 40224 10528 40288
rect 10208 40223 10528 40224
rect 19472 40288 19792 40289
rect 19472 40224 19480 40288
rect 19544 40224 19560 40288
rect 19624 40224 19640 40288
rect 19704 40224 19720 40288
rect 19784 40224 19792 40288
rect 19472 40223 19792 40224
rect 28165 40218 28231 40221
rect 29200 40218 30000 40308
rect 28165 40216 30000 40218
rect 28165 40160 28170 40216
rect 28226 40160 30000 40216
rect 28165 40158 30000 40160
rect 28165 40155 28231 40158
rect 29200 40068 30000 40158
rect 5576 39744 5896 39745
rect 5576 39680 5584 39744
rect 5648 39680 5664 39744
rect 5728 39680 5744 39744
rect 5808 39680 5824 39744
rect 5888 39680 5896 39744
rect 5576 39679 5896 39680
rect 14840 39744 15160 39745
rect 14840 39680 14848 39744
rect 14912 39680 14928 39744
rect 14992 39680 15008 39744
rect 15072 39680 15088 39744
rect 15152 39680 15160 39744
rect 14840 39679 15160 39680
rect 24104 39744 24424 39745
rect 24104 39680 24112 39744
rect 24176 39680 24192 39744
rect 24256 39680 24272 39744
rect 24336 39680 24352 39744
rect 24416 39680 24424 39744
rect 24104 39679 24424 39680
rect 0 39388 800 39628
rect 28717 39538 28783 39541
rect 29200 39538 30000 39628
rect 28717 39536 30000 39538
rect 28717 39480 28722 39536
rect 28778 39480 30000 39536
rect 28717 39478 30000 39480
rect 28717 39475 28783 39478
rect 29200 39388 30000 39478
rect 10208 39200 10528 39201
rect 10208 39136 10216 39200
rect 10280 39136 10296 39200
rect 10360 39136 10376 39200
rect 10440 39136 10456 39200
rect 10520 39136 10528 39200
rect 10208 39135 10528 39136
rect 19472 39200 19792 39201
rect 19472 39136 19480 39200
rect 19544 39136 19560 39200
rect 19624 39136 19640 39200
rect 19704 39136 19720 39200
rect 19784 39136 19792 39200
rect 19472 39135 19792 39136
rect 0 38858 800 38948
rect 2773 38858 2839 38861
rect 0 38856 2839 38858
rect 0 38800 2778 38856
rect 2834 38800 2839 38856
rect 0 38798 2839 38800
rect 0 38708 800 38798
rect 2773 38795 2839 38798
rect 5576 38656 5896 38657
rect 5576 38592 5584 38656
rect 5648 38592 5664 38656
rect 5728 38592 5744 38656
rect 5808 38592 5824 38656
rect 5888 38592 5896 38656
rect 5576 38591 5896 38592
rect 14840 38656 15160 38657
rect 14840 38592 14848 38656
rect 14912 38592 14928 38656
rect 14992 38592 15008 38656
rect 15072 38592 15088 38656
rect 15152 38592 15160 38656
rect 14840 38591 15160 38592
rect 24104 38656 24424 38657
rect 24104 38592 24112 38656
rect 24176 38592 24192 38656
rect 24256 38592 24272 38656
rect 24336 38592 24352 38656
rect 24416 38592 24424 38656
rect 24104 38591 24424 38592
rect 10208 38112 10528 38113
rect 10208 38048 10216 38112
rect 10280 38048 10296 38112
rect 10360 38048 10376 38112
rect 10440 38048 10456 38112
rect 10520 38048 10528 38112
rect 10208 38047 10528 38048
rect 19472 38112 19792 38113
rect 19472 38048 19480 38112
rect 19544 38048 19560 38112
rect 19624 38048 19640 38112
rect 19704 38048 19720 38112
rect 19784 38048 19792 38112
rect 19472 38047 19792 38048
rect 29200 38028 30000 38268
rect 0 37498 800 37588
rect 5576 37568 5896 37569
rect 5576 37504 5584 37568
rect 5648 37504 5664 37568
rect 5728 37504 5744 37568
rect 5808 37504 5824 37568
rect 5888 37504 5896 37568
rect 5576 37503 5896 37504
rect 14840 37568 15160 37569
rect 14840 37504 14848 37568
rect 14912 37504 14928 37568
rect 14992 37504 15008 37568
rect 15072 37504 15088 37568
rect 15152 37504 15160 37568
rect 14840 37503 15160 37504
rect 24104 37568 24424 37569
rect 24104 37504 24112 37568
rect 24176 37504 24192 37568
rect 24256 37504 24272 37568
rect 24336 37504 24352 37568
rect 24416 37504 24424 37568
rect 24104 37503 24424 37504
rect 1393 37498 1459 37501
rect 0 37496 1459 37498
rect 0 37440 1398 37496
rect 1454 37440 1459 37496
rect 0 37438 1459 37440
rect 0 37348 800 37438
rect 1393 37435 1459 37438
rect 29200 37348 30000 37588
rect 10208 37024 10528 37025
rect 10208 36960 10216 37024
rect 10280 36960 10296 37024
rect 10360 36960 10376 37024
rect 10440 36960 10456 37024
rect 10520 36960 10528 37024
rect 10208 36959 10528 36960
rect 19472 37024 19792 37025
rect 19472 36960 19480 37024
rect 19544 36960 19560 37024
rect 19624 36960 19640 37024
rect 19704 36960 19720 37024
rect 19784 36960 19792 37024
rect 19472 36959 19792 36960
rect 0 36818 800 36908
rect 1853 36818 1919 36821
rect 0 36816 1919 36818
rect 0 36760 1858 36816
rect 1914 36760 1919 36816
rect 0 36758 1919 36760
rect 0 36668 800 36758
rect 1853 36755 1919 36758
rect 26785 36818 26851 36821
rect 29200 36818 30000 36908
rect 26785 36816 30000 36818
rect 26785 36760 26790 36816
rect 26846 36760 30000 36816
rect 26785 36758 30000 36760
rect 26785 36755 26851 36758
rect 29200 36668 30000 36758
rect 5576 36480 5896 36481
rect 5576 36416 5584 36480
rect 5648 36416 5664 36480
rect 5728 36416 5744 36480
rect 5808 36416 5824 36480
rect 5888 36416 5896 36480
rect 5576 36415 5896 36416
rect 14840 36480 15160 36481
rect 14840 36416 14848 36480
rect 14912 36416 14928 36480
rect 14992 36416 15008 36480
rect 15072 36416 15088 36480
rect 15152 36416 15160 36480
rect 14840 36415 15160 36416
rect 24104 36480 24424 36481
rect 24104 36416 24112 36480
rect 24176 36416 24192 36480
rect 24256 36416 24272 36480
rect 24336 36416 24352 36480
rect 24416 36416 24424 36480
rect 24104 36415 24424 36416
rect 0 36138 800 36228
rect 2773 36138 2839 36141
rect 0 36136 2839 36138
rect 0 36080 2778 36136
rect 2834 36080 2839 36136
rect 0 36078 2839 36080
rect 0 35988 800 36078
rect 2773 36075 2839 36078
rect 27521 36138 27587 36141
rect 29200 36138 30000 36228
rect 27521 36136 30000 36138
rect 27521 36080 27526 36136
rect 27582 36080 30000 36136
rect 27521 36078 30000 36080
rect 27521 36075 27587 36078
rect 29200 35988 30000 36078
rect 10208 35936 10528 35937
rect 10208 35872 10216 35936
rect 10280 35872 10296 35936
rect 10360 35872 10376 35936
rect 10440 35872 10456 35936
rect 10520 35872 10528 35936
rect 10208 35871 10528 35872
rect 19472 35936 19792 35937
rect 19472 35872 19480 35936
rect 19544 35872 19560 35936
rect 19624 35872 19640 35936
rect 19704 35872 19720 35936
rect 19784 35872 19792 35936
rect 19472 35871 19792 35872
rect 0 35308 800 35548
rect 5576 35392 5896 35393
rect 5576 35328 5584 35392
rect 5648 35328 5664 35392
rect 5728 35328 5744 35392
rect 5808 35328 5824 35392
rect 5888 35328 5896 35392
rect 5576 35327 5896 35328
rect 14840 35392 15160 35393
rect 14840 35328 14848 35392
rect 14912 35328 14928 35392
rect 14992 35328 15008 35392
rect 15072 35328 15088 35392
rect 15152 35328 15160 35392
rect 14840 35327 15160 35328
rect 24104 35392 24424 35393
rect 24104 35328 24112 35392
rect 24176 35328 24192 35392
rect 24256 35328 24272 35392
rect 24336 35328 24352 35392
rect 24416 35328 24424 35392
rect 24104 35327 24424 35328
rect 29200 35308 30000 35548
rect 10593 35186 10659 35189
rect 18321 35186 18387 35189
rect 18638 35186 18644 35188
rect 10593 35184 18644 35186
rect 10593 35128 10598 35184
rect 10654 35128 18326 35184
rect 18382 35128 18644 35184
rect 10593 35126 18644 35128
rect 10593 35123 10659 35126
rect 18321 35123 18387 35126
rect 18638 35124 18644 35126
rect 18708 35124 18714 35188
rect 0 34778 800 34868
rect 10208 34848 10528 34849
rect 10208 34784 10216 34848
rect 10280 34784 10296 34848
rect 10360 34784 10376 34848
rect 10440 34784 10456 34848
rect 10520 34784 10528 34848
rect 10208 34783 10528 34784
rect 19472 34848 19792 34849
rect 19472 34784 19480 34848
rect 19544 34784 19560 34848
rect 19624 34784 19640 34848
rect 19704 34784 19720 34848
rect 19784 34784 19792 34848
rect 19472 34783 19792 34784
rect 1761 34778 1827 34781
rect 0 34776 1827 34778
rect 0 34720 1766 34776
rect 1822 34720 1827 34776
rect 0 34718 1827 34720
rect 0 34628 800 34718
rect 1761 34715 1827 34718
rect 27429 34644 27495 34645
rect 27429 34640 27476 34644
rect 27540 34642 27546 34644
rect 27429 34584 27434 34640
rect 27429 34580 27476 34584
rect 27540 34582 27586 34642
rect 29200 34628 30000 34868
rect 27540 34580 27546 34582
rect 27429 34579 27495 34580
rect 5576 34304 5896 34305
rect 5576 34240 5584 34304
rect 5648 34240 5664 34304
rect 5728 34240 5744 34304
rect 5808 34240 5824 34304
rect 5888 34240 5896 34304
rect 5576 34239 5896 34240
rect 14840 34304 15160 34305
rect 14840 34240 14848 34304
rect 14912 34240 14928 34304
rect 14992 34240 15008 34304
rect 15072 34240 15088 34304
rect 15152 34240 15160 34304
rect 14840 34239 15160 34240
rect 24104 34304 24424 34305
rect 24104 34240 24112 34304
rect 24176 34240 24192 34304
rect 24256 34240 24272 34304
rect 24336 34240 24352 34304
rect 24416 34240 24424 34304
rect 24104 34239 24424 34240
rect 0 33948 800 34188
rect 27521 34098 27587 34101
rect 29200 34098 30000 34188
rect 27521 34096 30000 34098
rect 27521 34040 27526 34096
rect 27582 34040 30000 34096
rect 27521 34038 30000 34040
rect 27521 34035 27587 34038
rect 21817 33964 21883 33965
rect 21766 33900 21772 33964
rect 21836 33962 21883 33964
rect 21836 33960 21928 33962
rect 21878 33904 21928 33960
rect 29200 33948 30000 34038
rect 21836 33902 21928 33904
rect 21836 33900 21883 33902
rect 21817 33899 21883 33900
rect 10208 33760 10528 33761
rect 10208 33696 10216 33760
rect 10280 33696 10296 33760
rect 10360 33696 10376 33760
rect 10440 33696 10456 33760
rect 10520 33696 10528 33760
rect 10208 33695 10528 33696
rect 19472 33760 19792 33761
rect 19472 33696 19480 33760
rect 19544 33696 19560 33760
rect 19624 33696 19640 33760
rect 19704 33696 19720 33760
rect 19784 33696 19792 33760
rect 19472 33695 19792 33696
rect 0 33418 800 33508
rect 3325 33418 3391 33421
rect 0 33416 3391 33418
rect 0 33360 3330 33416
rect 3386 33360 3391 33416
rect 0 33358 3391 33360
rect 0 33268 800 33358
rect 3325 33355 3391 33358
rect 5576 33216 5896 33217
rect 5576 33152 5584 33216
rect 5648 33152 5664 33216
rect 5728 33152 5744 33216
rect 5808 33152 5824 33216
rect 5888 33152 5896 33216
rect 5576 33151 5896 33152
rect 14840 33216 15160 33217
rect 14840 33152 14848 33216
rect 14912 33152 14928 33216
rect 14992 33152 15008 33216
rect 15072 33152 15088 33216
rect 15152 33152 15160 33216
rect 14840 33151 15160 33152
rect 24104 33216 24424 33217
rect 24104 33152 24112 33216
rect 24176 33152 24192 33216
rect 24256 33152 24272 33216
rect 24336 33152 24352 33216
rect 24416 33152 24424 33216
rect 24104 33151 24424 33152
rect 25957 32738 26023 32741
rect 29200 32738 30000 32828
rect 25957 32736 30000 32738
rect 25957 32680 25962 32736
rect 26018 32680 30000 32736
rect 25957 32678 30000 32680
rect 25957 32675 26023 32678
rect 10208 32672 10528 32673
rect 10208 32608 10216 32672
rect 10280 32608 10296 32672
rect 10360 32608 10376 32672
rect 10440 32608 10456 32672
rect 10520 32608 10528 32672
rect 10208 32607 10528 32608
rect 19472 32672 19792 32673
rect 19472 32608 19480 32672
rect 19544 32608 19560 32672
rect 19624 32608 19640 32672
rect 19704 32608 19720 32672
rect 19784 32608 19792 32672
rect 19472 32607 19792 32608
rect 29200 32588 30000 32678
rect 22369 32330 22435 32333
rect 22502 32330 22508 32332
rect 22369 32328 22508 32330
rect 22369 32272 22374 32328
rect 22430 32272 22508 32328
rect 22369 32270 22508 32272
rect 22369 32267 22435 32270
rect 22502 32268 22508 32270
rect 22572 32268 22578 32332
rect 0 32058 800 32148
rect 5576 32128 5896 32129
rect 5576 32064 5584 32128
rect 5648 32064 5664 32128
rect 5728 32064 5744 32128
rect 5808 32064 5824 32128
rect 5888 32064 5896 32128
rect 5576 32063 5896 32064
rect 14840 32128 15160 32129
rect 14840 32064 14848 32128
rect 14912 32064 14928 32128
rect 14992 32064 15008 32128
rect 15072 32064 15088 32128
rect 15152 32064 15160 32128
rect 14840 32063 15160 32064
rect 24104 32128 24424 32129
rect 24104 32064 24112 32128
rect 24176 32064 24192 32128
rect 24256 32064 24272 32128
rect 24336 32064 24352 32128
rect 24416 32064 24424 32128
rect 24104 32063 24424 32064
rect 1853 32058 1919 32061
rect 0 32056 1919 32058
rect 0 32000 1858 32056
rect 1914 32000 1919 32056
rect 0 31998 1919 32000
rect 0 31908 800 31998
rect 1853 31995 1919 31998
rect 28625 32058 28691 32061
rect 29200 32058 30000 32148
rect 28625 32056 30000 32058
rect 28625 32000 28630 32056
rect 28686 32000 30000 32056
rect 28625 31998 30000 32000
rect 28625 31995 28691 31998
rect 29200 31908 30000 31998
rect 10208 31584 10528 31585
rect 10208 31520 10216 31584
rect 10280 31520 10296 31584
rect 10360 31520 10376 31584
rect 10440 31520 10456 31584
rect 10520 31520 10528 31584
rect 10208 31519 10528 31520
rect 19472 31584 19792 31585
rect 19472 31520 19480 31584
rect 19544 31520 19560 31584
rect 19624 31520 19640 31584
rect 19704 31520 19720 31584
rect 19784 31520 19792 31584
rect 19472 31519 19792 31520
rect 0 31228 800 31468
rect 28717 31378 28783 31381
rect 29200 31378 30000 31468
rect 28717 31376 30000 31378
rect 28717 31320 28722 31376
rect 28778 31320 30000 31376
rect 28717 31318 30000 31320
rect 28717 31315 28783 31318
rect 29200 31228 30000 31318
rect 5576 31040 5896 31041
rect 5576 30976 5584 31040
rect 5648 30976 5664 31040
rect 5728 30976 5744 31040
rect 5808 30976 5824 31040
rect 5888 30976 5896 31040
rect 5576 30975 5896 30976
rect 14840 31040 15160 31041
rect 14840 30976 14848 31040
rect 14912 30976 14928 31040
rect 14992 30976 15008 31040
rect 15072 30976 15088 31040
rect 15152 30976 15160 31040
rect 14840 30975 15160 30976
rect 24104 31040 24424 31041
rect 24104 30976 24112 31040
rect 24176 30976 24192 31040
rect 24256 30976 24272 31040
rect 24336 30976 24352 31040
rect 24416 30976 24424 31040
rect 24104 30975 24424 30976
rect 0 30548 800 30788
rect 27521 30698 27587 30701
rect 29200 30698 30000 30788
rect 27521 30696 30000 30698
rect 27521 30640 27526 30696
rect 27582 30640 30000 30696
rect 27521 30638 30000 30640
rect 27521 30635 27587 30638
rect 29200 30548 30000 30638
rect 10208 30496 10528 30497
rect 10208 30432 10216 30496
rect 10280 30432 10296 30496
rect 10360 30432 10376 30496
rect 10440 30432 10456 30496
rect 10520 30432 10528 30496
rect 10208 30431 10528 30432
rect 19472 30496 19792 30497
rect 19472 30432 19480 30496
rect 19544 30432 19560 30496
rect 19624 30432 19640 30496
rect 19704 30432 19720 30496
rect 19784 30432 19792 30496
rect 19472 30431 19792 30432
rect 0 30018 800 30108
rect 1393 30018 1459 30021
rect 0 30016 1459 30018
rect 0 29960 1398 30016
rect 1454 29960 1459 30016
rect 0 29958 1459 29960
rect 0 29868 800 29958
rect 1393 29955 1459 29958
rect 27337 30018 27403 30021
rect 29200 30018 30000 30108
rect 27337 30016 30000 30018
rect 27337 29960 27342 30016
rect 27398 29960 30000 30016
rect 27337 29958 30000 29960
rect 27337 29955 27403 29958
rect 5576 29952 5896 29953
rect 5576 29888 5584 29952
rect 5648 29888 5664 29952
rect 5728 29888 5744 29952
rect 5808 29888 5824 29952
rect 5888 29888 5896 29952
rect 5576 29887 5896 29888
rect 14840 29952 15160 29953
rect 14840 29888 14848 29952
rect 14912 29888 14928 29952
rect 14992 29888 15008 29952
rect 15072 29888 15088 29952
rect 15152 29888 15160 29952
rect 14840 29887 15160 29888
rect 24104 29952 24424 29953
rect 24104 29888 24112 29952
rect 24176 29888 24192 29952
rect 24256 29888 24272 29952
rect 24336 29888 24352 29952
rect 24416 29888 24424 29952
rect 24104 29887 24424 29888
rect 29200 29868 30000 29958
rect 0 29188 800 29428
rect 10208 29408 10528 29409
rect 10208 29344 10216 29408
rect 10280 29344 10296 29408
rect 10360 29344 10376 29408
rect 10440 29344 10456 29408
rect 10520 29344 10528 29408
rect 10208 29343 10528 29344
rect 19472 29408 19792 29409
rect 19472 29344 19480 29408
rect 19544 29344 19560 29408
rect 19624 29344 19640 29408
rect 19704 29344 19720 29408
rect 19784 29344 19792 29408
rect 19472 29343 19792 29344
rect 25037 29338 25103 29341
rect 29200 29338 30000 29428
rect 25037 29336 30000 29338
rect 25037 29280 25042 29336
rect 25098 29280 30000 29336
rect 25037 29278 30000 29280
rect 25037 29275 25103 29278
rect 29200 29188 30000 29278
rect 5576 28864 5896 28865
rect 5576 28800 5584 28864
rect 5648 28800 5664 28864
rect 5728 28800 5744 28864
rect 5808 28800 5824 28864
rect 5888 28800 5896 28864
rect 5576 28799 5896 28800
rect 14840 28864 15160 28865
rect 14840 28800 14848 28864
rect 14912 28800 14928 28864
rect 14992 28800 15008 28864
rect 15072 28800 15088 28864
rect 15152 28800 15160 28864
rect 14840 28799 15160 28800
rect 24104 28864 24424 28865
rect 24104 28800 24112 28864
rect 24176 28800 24192 28864
rect 24256 28800 24272 28864
rect 24336 28800 24352 28864
rect 24416 28800 24424 28864
rect 24104 28799 24424 28800
rect 0 28508 800 28748
rect 27521 28658 27587 28661
rect 29200 28658 30000 28748
rect 27521 28656 30000 28658
rect 27521 28600 27526 28656
rect 27582 28600 30000 28656
rect 27521 28598 30000 28600
rect 27521 28595 27587 28598
rect 29200 28508 30000 28598
rect 10208 28320 10528 28321
rect 10208 28256 10216 28320
rect 10280 28256 10296 28320
rect 10360 28256 10376 28320
rect 10440 28256 10456 28320
rect 10520 28256 10528 28320
rect 10208 28255 10528 28256
rect 19472 28320 19792 28321
rect 19472 28256 19480 28320
rect 19544 28256 19560 28320
rect 19624 28256 19640 28320
rect 19704 28256 19720 28320
rect 19784 28256 19792 28320
rect 19472 28255 19792 28256
rect 0 27978 800 28068
rect 1393 27978 1459 27981
rect 0 27976 1459 27978
rect 0 27920 1398 27976
rect 1454 27920 1459 27976
rect 0 27918 1459 27920
rect 0 27828 800 27918
rect 1393 27915 1459 27918
rect 5576 27776 5896 27777
rect 5576 27712 5584 27776
rect 5648 27712 5664 27776
rect 5728 27712 5744 27776
rect 5808 27712 5824 27776
rect 5888 27712 5896 27776
rect 5576 27711 5896 27712
rect 14840 27776 15160 27777
rect 14840 27712 14848 27776
rect 14912 27712 14928 27776
rect 14992 27712 15008 27776
rect 15072 27712 15088 27776
rect 15152 27712 15160 27776
rect 14840 27711 15160 27712
rect 24104 27776 24424 27777
rect 24104 27712 24112 27776
rect 24176 27712 24192 27776
rect 24256 27712 24272 27776
rect 24336 27712 24352 27776
rect 24416 27712 24424 27776
rect 24104 27711 24424 27712
rect 27521 27298 27587 27301
rect 29200 27298 30000 27388
rect 27521 27296 30000 27298
rect 27521 27240 27526 27296
rect 27582 27240 30000 27296
rect 27521 27238 30000 27240
rect 27521 27235 27587 27238
rect 10208 27232 10528 27233
rect 10208 27168 10216 27232
rect 10280 27168 10296 27232
rect 10360 27168 10376 27232
rect 10440 27168 10456 27232
rect 10520 27168 10528 27232
rect 10208 27167 10528 27168
rect 19472 27232 19792 27233
rect 19472 27168 19480 27232
rect 19544 27168 19560 27232
rect 19624 27168 19640 27232
rect 19704 27168 19720 27232
rect 19784 27168 19792 27232
rect 19472 27167 19792 27168
rect 29200 27148 30000 27238
rect 0 26468 800 26708
rect 5576 26688 5896 26689
rect 5576 26624 5584 26688
rect 5648 26624 5664 26688
rect 5728 26624 5744 26688
rect 5808 26624 5824 26688
rect 5888 26624 5896 26688
rect 5576 26623 5896 26624
rect 14840 26688 15160 26689
rect 14840 26624 14848 26688
rect 14912 26624 14928 26688
rect 14992 26624 15008 26688
rect 15072 26624 15088 26688
rect 15152 26624 15160 26688
rect 14840 26623 15160 26624
rect 24104 26688 24424 26689
rect 24104 26624 24112 26688
rect 24176 26624 24192 26688
rect 24256 26624 24272 26688
rect 24336 26624 24352 26688
rect 24416 26624 24424 26688
rect 24104 26623 24424 26624
rect 25773 26618 25839 26621
rect 29200 26618 30000 26708
rect 25773 26616 30000 26618
rect 25773 26560 25778 26616
rect 25834 26560 30000 26616
rect 25773 26558 30000 26560
rect 25773 26555 25839 26558
rect 29200 26468 30000 26558
rect 10208 26144 10528 26145
rect 10208 26080 10216 26144
rect 10280 26080 10296 26144
rect 10360 26080 10376 26144
rect 10440 26080 10456 26144
rect 10520 26080 10528 26144
rect 10208 26079 10528 26080
rect 19472 26144 19792 26145
rect 19472 26080 19480 26144
rect 19544 26080 19560 26144
rect 19624 26080 19640 26144
rect 19704 26080 19720 26144
rect 19784 26080 19792 26144
rect 19472 26079 19792 26080
rect 0 25938 800 26028
rect 2773 25938 2839 25941
rect 0 25936 2839 25938
rect 0 25880 2778 25936
rect 2834 25880 2839 25936
rect 0 25878 2839 25880
rect 0 25788 800 25878
rect 2773 25875 2839 25878
rect 29200 25788 30000 26028
rect 5576 25600 5896 25601
rect 5576 25536 5584 25600
rect 5648 25536 5664 25600
rect 5728 25536 5744 25600
rect 5808 25536 5824 25600
rect 5888 25536 5896 25600
rect 5576 25535 5896 25536
rect 14840 25600 15160 25601
rect 14840 25536 14848 25600
rect 14912 25536 14928 25600
rect 14992 25536 15008 25600
rect 15072 25536 15088 25600
rect 15152 25536 15160 25600
rect 14840 25535 15160 25536
rect 24104 25600 24424 25601
rect 24104 25536 24112 25600
rect 24176 25536 24192 25600
rect 24256 25536 24272 25600
rect 24336 25536 24352 25600
rect 24416 25536 24424 25600
rect 24104 25535 24424 25536
rect 0 25258 800 25348
rect 1393 25258 1459 25261
rect 0 25256 1459 25258
rect 0 25200 1398 25256
rect 1454 25200 1459 25256
rect 0 25198 1459 25200
rect 0 25108 800 25198
rect 1393 25195 1459 25198
rect 27521 25258 27587 25261
rect 29200 25258 30000 25348
rect 27521 25256 30000 25258
rect 27521 25200 27526 25256
rect 27582 25200 30000 25256
rect 27521 25198 30000 25200
rect 27521 25195 27587 25198
rect 29200 25108 30000 25198
rect 10208 25056 10528 25057
rect 10208 24992 10216 25056
rect 10280 24992 10296 25056
rect 10360 24992 10376 25056
rect 10440 24992 10456 25056
rect 10520 24992 10528 25056
rect 10208 24991 10528 24992
rect 19472 25056 19792 25057
rect 19472 24992 19480 25056
rect 19544 24992 19560 25056
rect 19624 24992 19640 25056
rect 19704 24992 19720 25056
rect 19784 24992 19792 25056
rect 19472 24991 19792 24992
rect 0 24428 800 24668
rect 25957 24578 26023 24581
rect 29200 24578 30000 24668
rect 25957 24576 30000 24578
rect 25957 24520 25962 24576
rect 26018 24520 30000 24576
rect 25957 24518 30000 24520
rect 25957 24515 26023 24518
rect 5576 24512 5896 24513
rect 5576 24448 5584 24512
rect 5648 24448 5664 24512
rect 5728 24448 5744 24512
rect 5808 24448 5824 24512
rect 5888 24448 5896 24512
rect 5576 24447 5896 24448
rect 14840 24512 15160 24513
rect 14840 24448 14848 24512
rect 14912 24448 14928 24512
rect 14992 24448 15008 24512
rect 15072 24448 15088 24512
rect 15152 24448 15160 24512
rect 14840 24447 15160 24448
rect 24104 24512 24424 24513
rect 24104 24448 24112 24512
rect 24176 24448 24192 24512
rect 24256 24448 24272 24512
rect 24336 24448 24352 24512
rect 24416 24448 24424 24512
rect 24104 24447 24424 24448
rect 29200 24428 30000 24518
rect 21950 24108 21956 24172
rect 22020 24170 22026 24172
rect 25037 24170 25103 24173
rect 22020 24168 25103 24170
rect 22020 24112 25042 24168
rect 25098 24112 25103 24168
rect 22020 24110 25103 24112
rect 22020 24108 22026 24110
rect 25037 24107 25103 24110
rect 0 23748 800 23988
rect 10208 23968 10528 23969
rect 10208 23904 10216 23968
rect 10280 23904 10296 23968
rect 10360 23904 10376 23968
rect 10440 23904 10456 23968
rect 10520 23904 10528 23968
rect 10208 23903 10528 23904
rect 19472 23968 19792 23969
rect 19472 23904 19480 23968
rect 19544 23904 19560 23968
rect 19624 23904 19640 23968
rect 19704 23904 19720 23968
rect 19784 23904 19792 23968
rect 19472 23903 19792 23904
rect 27521 23898 27587 23901
rect 29200 23898 30000 23988
rect 27521 23896 30000 23898
rect 27521 23840 27526 23896
rect 27582 23840 30000 23896
rect 27521 23838 30000 23840
rect 27521 23835 27587 23838
rect 29200 23748 30000 23838
rect 21766 23428 21772 23492
rect 21836 23490 21842 23492
rect 22001 23490 22067 23493
rect 21836 23488 22067 23490
rect 21836 23432 22006 23488
rect 22062 23432 22067 23488
rect 21836 23430 22067 23432
rect 21836 23428 21842 23430
rect 22001 23427 22067 23430
rect 5576 23424 5896 23425
rect 5576 23360 5584 23424
rect 5648 23360 5664 23424
rect 5728 23360 5744 23424
rect 5808 23360 5824 23424
rect 5888 23360 5896 23424
rect 5576 23359 5896 23360
rect 14840 23424 15160 23425
rect 14840 23360 14848 23424
rect 14912 23360 14928 23424
rect 14992 23360 15008 23424
rect 15072 23360 15088 23424
rect 15152 23360 15160 23424
rect 14840 23359 15160 23360
rect 24104 23424 24424 23425
rect 24104 23360 24112 23424
rect 24176 23360 24192 23424
rect 24256 23360 24272 23424
rect 24336 23360 24352 23424
rect 24416 23360 24424 23424
rect 24104 23359 24424 23360
rect 0 23068 800 23308
rect 29200 23068 30000 23308
rect 10208 22880 10528 22881
rect 10208 22816 10216 22880
rect 10280 22816 10296 22880
rect 10360 22816 10376 22880
rect 10440 22816 10456 22880
rect 10520 22816 10528 22880
rect 10208 22815 10528 22816
rect 19472 22880 19792 22881
rect 19472 22816 19480 22880
rect 19544 22816 19560 22880
rect 19624 22816 19640 22880
rect 19704 22816 19720 22880
rect 19784 22816 19792 22880
rect 19472 22815 19792 22816
rect 0 22388 800 22628
rect 5576 22336 5896 22337
rect 5576 22272 5584 22336
rect 5648 22272 5664 22336
rect 5728 22272 5744 22336
rect 5808 22272 5824 22336
rect 5888 22272 5896 22336
rect 5576 22271 5896 22272
rect 14840 22336 15160 22337
rect 14840 22272 14848 22336
rect 14912 22272 14928 22336
rect 14992 22272 15008 22336
rect 15072 22272 15088 22336
rect 15152 22272 15160 22336
rect 14840 22271 15160 22272
rect 24104 22336 24424 22337
rect 24104 22272 24112 22336
rect 24176 22272 24192 22336
rect 24256 22272 24272 22336
rect 24336 22272 24352 22336
rect 24416 22272 24424 22336
rect 24104 22271 24424 22272
rect 28165 21858 28231 21861
rect 29200 21858 30000 21948
rect 28165 21856 30000 21858
rect 28165 21800 28170 21856
rect 28226 21800 30000 21856
rect 28165 21798 30000 21800
rect 28165 21795 28231 21798
rect 10208 21792 10528 21793
rect 10208 21728 10216 21792
rect 10280 21728 10296 21792
rect 10360 21728 10376 21792
rect 10440 21728 10456 21792
rect 10520 21728 10528 21792
rect 10208 21727 10528 21728
rect 19472 21792 19792 21793
rect 19472 21728 19480 21792
rect 19544 21728 19560 21792
rect 19624 21728 19640 21792
rect 19704 21728 19720 21792
rect 19784 21728 19792 21792
rect 19472 21727 19792 21728
rect 29200 21708 30000 21798
rect 22001 21586 22067 21589
rect 22502 21586 22508 21588
rect 22001 21584 22508 21586
rect 22001 21528 22006 21584
rect 22062 21528 22508 21584
rect 22001 21526 22508 21528
rect 22001 21523 22067 21526
rect 22502 21524 22508 21526
rect 22572 21524 22578 21588
rect 0 21028 800 21268
rect 5576 21248 5896 21249
rect 5576 21184 5584 21248
rect 5648 21184 5664 21248
rect 5728 21184 5744 21248
rect 5808 21184 5824 21248
rect 5888 21184 5896 21248
rect 5576 21183 5896 21184
rect 14840 21248 15160 21249
rect 14840 21184 14848 21248
rect 14912 21184 14928 21248
rect 14992 21184 15008 21248
rect 15072 21184 15088 21248
rect 15152 21184 15160 21248
rect 14840 21183 15160 21184
rect 24104 21248 24424 21249
rect 24104 21184 24112 21248
rect 24176 21184 24192 21248
rect 24256 21184 24272 21248
rect 24336 21184 24352 21248
rect 24416 21184 24424 21248
rect 24104 21183 24424 21184
rect 26141 21178 26207 21181
rect 29200 21178 30000 21268
rect 26141 21176 30000 21178
rect 26141 21120 26146 21176
rect 26202 21120 30000 21176
rect 26141 21118 30000 21120
rect 26141 21115 26207 21118
rect 29200 21028 30000 21118
rect 10208 20704 10528 20705
rect 10208 20640 10216 20704
rect 10280 20640 10296 20704
rect 10360 20640 10376 20704
rect 10440 20640 10456 20704
rect 10520 20640 10528 20704
rect 10208 20639 10528 20640
rect 19472 20704 19792 20705
rect 19472 20640 19480 20704
rect 19544 20640 19560 20704
rect 19624 20640 19640 20704
rect 19704 20640 19720 20704
rect 19784 20640 19792 20704
rect 19472 20639 19792 20640
rect 0 20348 800 20588
rect 28165 20498 28231 20501
rect 29200 20498 30000 20588
rect 28165 20496 30000 20498
rect 28165 20440 28170 20496
rect 28226 20440 30000 20496
rect 28165 20438 30000 20440
rect 28165 20435 28231 20438
rect 27337 20364 27403 20365
rect 27286 20300 27292 20364
rect 27356 20362 27403 20364
rect 27356 20360 27448 20362
rect 27398 20304 27448 20360
rect 29200 20348 30000 20438
rect 27356 20302 27448 20304
rect 27356 20300 27403 20302
rect 27337 20299 27403 20300
rect 5576 20160 5896 20161
rect 5576 20096 5584 20160
rect 5648 20096 5664 20160
rect 5728 20096 5744 20160
rect 5808 20096 5824 20160
rect 5888 20096 5896 20160
rect 5576 20095 5896 20096
rect 14840 20160 15160 20161
rect 14840 20096 14848 20160
rect 14912 20096 14928 20160
rect 14992 20096 15008 20160
rect 15072 20096 15088 20160
rect 15152 20096 15160 20160
rect 14840 20095 15160 20096
rect 24104 20160 24424 20161
rect 24104 20096 24112 20160
rect 24176 20096 24192 20160
rect 24256 20096 24272 20160
rect 24336 20096 24352 20160
rect 24416 20096 24424 20160
rect 24104 20095 24424 20096
rect 0 19818 800 19908
rect 2957 19818 3023 19821
rect 0 19816 3023 19818
rect 0 19760 2962 19816
rect 3018 19760 3023 19816
rect 0 19758 3023 19760
rect 0 19668 800 19758
rect 2957 19755 3023 19758
rect 27337 19818 27403 19821
rect 29200 19818 30000 19908
rect 27337 19816 30000 19818
rect 27337 19760 27342 19816
rect 27398 19760 30000 19816
rect 27337 19758 30000 19760
rect 27337 19755 27403 19758
rect 29200 19668 30000 19758
rect 10208 19616 10528 19617
rect 10208 19552 10216 19616
rect 10280 19552 10296 19616
rect 10360 19552 10376 19616
rect 10440 19552 10456 19616
rect 10520 19552 10528 19616
rect 10208 19551 10528 19552
rect 19472 19616 19792 19617
rect 19472 19552 19480 19616
rect 19544 19552 19560 19616
rect 19624 19552 19640 19616
rect 19704 19552 19720 19616
rect 19784 19552 19792 19616
rect 19472 19551 19792 19552
rect 0 19138 800 19228
rect 1853 19138 1919 19141
rect 0 19136 1919 19138
rect 0 19080 1858 19136
rect 1914 19080 1919 19136
rect 0 19078 1919 19080
rect 0 18988 800 19078
rect 1853 19075 1919 19078
rect 5576 19072 5896 19073
rect 5576 19008 5584 19072
rect 5648 19008 5664 19072
rect 5728 19008 5744 19072
rect 5808 19008 5824 19072
rect 5888 19008 5896 19072
rect 5576 19007 5896 19008
rect 14840 19072 15160 19073
rect 14840 19008 14848 19072
rect 14912 19008 14928 19072
rect 14992 19008 15008 19072
rect 15072 19008 15088 19072
rect 15152 19008 15160 19072
rect 14840 19007 15160 19008
rect 24104 19072 24424 19073
rect 24104 19008 24112 19072
rect 24176 19008 24192 19072
rect 24256 19008 24272 19072
rect 24336 19008 24352 19072
rect 24416 19008 24424 19072
rect 24104 19007 24424 19008
rect 29200 18988 30000 19228
rect 0 18458 800 18548
rect 10208 18528 10528 18529
rect 10208 18464 10216 18528
rect 10280 18464 10296 18528
rect 10360 18464 10376 18528
rect 10440 18464 10456 18528
rect 10520 18464 10528 18528
rect 10208 18463 10528 18464
rect 19472 18528 19792 18529
rect 19472 18464 19480 18528
rect 19544 18464 19560 18528
rect 19624 18464 19640 18528
rect 19704 18464 19720 18528
rect 19784 18464 19792 18528
rect 19472 18463 19792 18464
rect 2405 18458 2471 18461
rect 0 18456 2471 18458
rect 0 18400 2410 18456
rect 2466 18400 2471 18456
rect 0 18398 2471 18400
rect 0 18308 800 18398
rect 2405 18395 2471 18398
rect 29200 18308 30000 18548
rect 5576 17984 5896 17985
rect 5576 17920 5584 17984
rect 5648 17920 5664 17984
rect 5728 17920 5744 17984
rect 5808 17920 5824 17984
rect 5888 17920 5896 17984
rect 5576 17919 5896 17920
rect 14840 17984 15160 17985
rect 14840 17920 14848 17984
rect 14912 17920 14928 17984
rect 14992 17920 15008 17984
rect 15072 17920 15088 17984
rect 15152 17920 15160 17984
rect 14840 17919 15160 17920
rect 24104 17984 24424 17985
rect 24104 17920 24112 17984
rect 24176 17920 24192 17984
rect 24256 17920 24272 17984
rect 24336 17920 24352 17984
rect 24416 17920 24424 17984
rect 24104 17919 24424 17920
rect 0 17778 800 17868
rect 2773 17778 2839 17781
rect 0 17776 2839 17778
rect 0 17720 2778 17776
rect 2834 17720 2839 17776
rect 0 17718 2839 17720
rect 0 17628 800 17718
rect 2773 17715 2839 17718
rect 29200 17628 30000 17868
rect 10208 17440 10528 17441
rect 10208 17376 10216 17440
rect 10280 17376 10296 17440
rect 10360 17376 10376 17440
rect 10440 17376 10456 17440
rect 10520 17376 10528 17440
rect 10208 17375 10528 17376
rect 19472 17440 19792 17441
rect 19472 17376 19480 17440
rect 19544 17376 19560 17440
rect 19624 17376 19640 17440
rect 19704 17376 19720 17440
rect 19784 17376 19792 17440
rect 19472 17375 19792 17376
rect 0 16948 800 17188
rect 5576 16896 5896 16897
rect 5576 16832 5584 16896
rect 5648 16832 5664 16896
rect 5728 16832 5744 16896
rect 5808 16832 5824 16896
rect 5888 16832 5896 16896
rect 5576 16831 5896 16832
rect 14840 16896 15160 16897
rect 14840 16832 14848 16896
rect 14912 16832 14928 16896
rect 14992 16832 15008 16896
rect 15072 16832 15088 16896
rect 15152 16832 15160 16896
rect 14840 16831 15160 16832
rect 24104 16896 24424 16897
rect 24104 16832 24112 16896
rect 24176 16832 24192 16896
rect 24256 16832 24272 16896
rect 24336 16832 24352 16896
rect 24416 16832 24424 16896
rect 24104 16831 24424 16832
rect 28073 16418 28139 16421
rect 29200 16418 30000 16508
rect 28073 16416 30000 16418
rect 28073 16360 28078 16416
rect 28134 16360 30000 16416
rect 28073 16358 30000 16360
rect 28073 16355 28139 16358
rect 10208 16352 10528 16353
rect 10208 16288 10216 16352
rect 10280 16288 10296 16352
rect 10360 16288 10376 16352
rect 10440 16288 10456 16352
rect 10520 16288 10528 16352
rect 10208 16287 10528 16288
rect 19472 16352 19792 16353
rect 19472 16288 19480 16352
rect 19544 16288 19560 16352
rect 19624 16288 19640 16352
rect 19704 16288 19720 16352
rect 19784 16288 19792 16352
rect 19472 16287 19792 16288
rect 29200 16268 30000 16358
rect 0 15738 800 15828
rect 5576 15808 5896 15809
rect 5576 15744 5584 15808
rect 5648 15744 5664 15808
rect 5728 15744 5744 15808
rect 5808 15744 5824 15808
rect 5888 15744 5896 15808
rect 5576 15743 5896 15744
rect 14840 15808 15160 15809
rect 14840 15744 14848 15808
rect 14912 15744 14928 15808
rect 14992 15744 15008 15808
rect 15072 15744 15088 15808
rect 15152 15744 15160 15808
rect 14840 15743 15160 15744
rect 24104 15808 24424 15809
rect 24104 15744 24112 15808
rect 24176 15744 24192 15808
rect 24256 15744 24272 15808
rect 24336 15744 24352 15808
rect 24416 15744 24424 15808
rect 24104 15743 24424 15744
rect 2773 15738 2839 15741
rect 0 15736 2839 15738
rect 0 15680 2778 15736
rect 2834 15680 2839 15736
rect 0 15678 2839 15680
rect 0 15588 800 15678
rect 2773 15675 2839 15678
rect 28165 15738 28231 15741
rect 29200 15738 30000 15828
rect 28165 15736 30000 15738
rect 28165 15680 28170 15736
rect 28226 15680 30000 15736
rect 28165 15678 30000 15680
rect 28165 15675 28231 15678
rect 3969 15602 4035 15605
rect 25221 15602 25287 15605
rect 3969 15600 25287 15602
rect 3969 15544 3974 15600
rect 4030 15544 25226 15600
rect 25282 15544 25287 15600
rect 29200 15588 30000 15678
rect 3969 15542 25287 15544
rect 3969 15539 4035 15542
rect 25221 15539 25287 15542
rect 10208 15264 10528 15265
rect 10208 15200 10216 15264
rect 10280 15200 10296 15264
rect 10360 15200 10376 15264
rect 10440 15200 10456 15264
rect 10520 15200 10528 15264
rect 10208 15199 10528 15200
rect 19472 15264 19792 15265
rect 19472 15200 19480 15264
rect 19544 15200 19560 15264
rect 19624 15200 19640 15264
rect 19704 15200 19720 15264
rect 19784 15200 19792 15264
rect 19472 15199 19792 15200
rect 0 14908 800 15148
rect 24853 15058 24919 15061
rect 29200 15058 30000 15148
rect 24853 15056 30000 15058
rect 24853 15000 24858 15056
rect 24914 15000 30000 15056
rect 24853 14998 30000 15000
rect 24853 14995 24919 14998
rect 29200 14908 30000 14998
rect 5576 14720 5896 14721
rect 5576 14656 5584 14720
rect 5648 14656 5664 14720
rect 5728 14656 5744 14720
rect 5808 14656 5824 14720
rect 5888 14656 5896 14720
rect 5576 14655 5896 14656
rect 14840 14720 15160 14721
rect 14840 14656 14848 14720
rect 14912 14656 14928 14720
rect 14992 14656 15008 14720
rect 15072 14656 15088 14720
rect 15152 14656 15160 14720
rect 14840 14655 15160 14656
rect 24104 14720 24424 14721
rect 24104 14656 24112 14720
rect 24176 14656 24192 14720
rect 24256 14656 24272 14720
rect 24336 14656 24352 14720
rect 24416 14656 24424 14720
rect 24104 14655 24424 14656
rect 0 14378 800 14468
rect 1853 14378 1919 14381
rect 0 14376 1919 14378
rect 0 14320 1858 14376
rect 1914 14320 1919 14376
rect 0 14318 1919 14320
rect 0 14228 800 14318
rect 1853 14315 1919 14318
rect 27521 14378 27587 14381
rect 29200 14378 30000 14468
rect 27521 14376 30000 14378
rect 27521 14320 27526 14376
rect 27582 14320 30000 14376
rect 27521 14318 30000 14320
rect 27521 14315 27587 14318
rect 29200 14228 30000 14318
rect 10208 14176 10528 14177
rect 10208 14112 10216 14176
rect 10280 14112 10296 14176
rect 10360 14112 10376 14176
rect 10440 14112 10456 14176
rect 10520 14112 10528 14176
rect 10208 14111 10528 14112
rect 19472 14176 19792 14177
rect 19472 14112 19480 14176
rect 19544 14112 19560 14176
rect 19624 14112 19640 14176
rect 19704 14112 19720 14176
rect 19784 14112 19792 14176
rect 19472 14111 19792 14112
rect 27470 13908 27476 13972
rect 27540 13970 27546 13972
rect 27797 13970 27863 13973
rect 27540 13968 27863 13970
rect 27540 13912 27802 13968
rect 27858 13912 27863 13968
rect 27540 13910 27863 13912
rect 27540 13908 27546 13910
rect 27797 13907 27863 13910
rect 0 13698 800 13788
rect 1945 13698 2011 13701
rect 0 13696 2011 13698
rect 0 13640 1950 13696
rect 2006 13640 2011 13696
rect 0 13638 2011 13640
rect 0 13548 800 13638
rect 1945 13635 2011 13638
rect 5576 13632 5896 13633
rect 5576 13568 5584 13632
rect 5648 13568 5664 13632
rect 5728 13568 5744 13632
rect 5808 13568 5824 13632
rect 5888 13568 5896 13632
rect 5576 13567 5896 13568
rect 14840 13632 15160 13633
rect 14840 13568 14848 13632
rect 14912 13568 14928 13632
rect 14992 13568 15008 13632
rect 15072 13568 15088 13632
rect 15152 13568 15160 13632
rect 14840 13567 15160 13568
rect 24104 13632 24424 13633
rect 24104 13568 24112 13632
rect 24176 13568 24192 13632
rect 24256 13568 24272 13632
rect 24336 13568 24352 13632
rect 24416 13568 24424 13632
rect 24104 13567 24424 13568
rect 29200 13548 30000 13788
rect 0 12868 800 13108
rect 10208 13088 10528 13089
rect 10208 13024 10216 13088
rect 10280 13024 10296 13088
rect 10360 13024 10376 13088
rect 10440 13024 10456 13088
rect 10520 13024 10528 13088
rect 10208 13023 10528 13024
rect 19472 13088 19792 13089
rect 19472 13024 19480 13088
rect 19544 13024 19560 13088
rect 19624 13024 19640 13088
rect 19704 13024 19720 13088
rect 19784 13024 19792 13088
rect 19472 13023 19792 13024
rect 29200 12868 30000 13108
rect 5576 12544 5896 12545
rect 5576 12480 5584 12544
rect 5648 12480 5664 12544
rect 5728 12480 5744 12544
rect 5808 12480 5824 12544
rect 5888 12480 5896 12544
rect 5576 12479 5896 12480
rect 14840 12544 15160 12545
rect 14840 12480 14848 12544
rect 14912 12480 14928 12544
rect 14992 12480 15008 12544
rect 15072 12480 15088 12544
rect 15152 12480 15160 12544
rect 14840 12479 15160 12480
rect 24104 12544 24424 12545
rect 24104 12480 24112 12544
rect 24176 12480 24192 12544
rect 24256 12480 24272 12544
rect 24336 12480 24352 12544
rect 24416 12480 24424 12544
rect 24104 12479 24424 12480
rect 0 12338 800 12428
rect 3325 12338 3391 12341
rect 0 12336 3391 12338
rect 0 12280 3330 12336
rect 3386 12280 3391 12336
rect 0 12278 3391 12280
rect 0 12188 800 12278
rect 3325 12275 3391 12278
rect 27521 12338 27587 12341
rect 29200 12338 30000 12428
rect 27521 12336 30000 12338
rect 27521 12280 27526 12336
rect 27582 12280 30000 12336
rect 27521 12278 30000 12280
rect 27521 12275 27587 12278
rect 29200 12188 30000 12278
rect 10208 12000 10528 12001
rect 10208 11936 10216 12000
rect 10280 11936 10296 12000
rect 10360 11936 10376 12000
rect 10440 11936 10456 12000
rect 10520 11936 10528 12000
rect 10208 11935 10528 11936
rect 19472 12000 19792 12001
rect 19472 11936 19480 12000
rect 19544 11936 19560 12000
rect 19624 11936 19640 12000
rect 19704 11936 19720 12000
rect 19784 11936 19792 12000
rect 19472 11935 19792 11936
rect 0 11658 800 11748
rect 1945 11658 2011 11661
rect 0 11656 2011 11658
rect 0 11600 1950 11656
rect 2006 11600 2011 11656
rect 0 11598 2011 11600
rect 0 11508 800 11598
rect 1945 11595 2011 11598
rect 5576 11456 5896 11457
rect 5576 11392 5584 11456
rect 5648 11392 5664 11456
rect 5728 11392 5744 11456
rect 5808 11392 5824 11456
rect 5888 11392 5896 11456
rect 5576 11391 5896 11392
rect 14840 11456 15160 11457
rect 14840 11392 14848 11456
rect 14912 11392 14928 11456
rect 14992 11392 15008 11456
rect 15072 11392 15088 11456
rect 15152 11392 15160 11456
rect 14840 11391 15160 11392
rect 24104 11456 24424 11457
rect 24104 11392 24112 11456
rect 24176 11392 24192 11456
rect 24256 11392 24272 11456
rect 24336 11392 24352 11456
rect 24416 11392 24424 11456
rect 24104 11391 24424 11392
rect 27521 10978 27587 10981
rect 29200 10978 30000 11068
rect 27521 10976 30000 10978
rect 27521 10920 27526 10976
rect 27582 10920 30000 10976
rect 27521 10918 30000 10920
rect 27521 10915 27587 10918
rect 10208 10912 10528 10913
rect 10208 10848 10216 10912
rect 10280 10848 10296 10912
rect 10360 10848 10376 10912
rect 10440 10848 10456 10912
rect 10520 10848 10528 10912
rect 10208 10847 10528 10848
rect 19472 10912 19792 10913
rect 19472 10848 19480 10912
rect 19544 10848 19560 10912
rect 19624 10848 19640 10912
rect 19704 10848 19720 10912
rect 19784 10848 19792 10912
rect 19472 10847 19792 10848
rect 29200 10828 30000 10918
rect 0 10148 800 10388
rect 5576 10368 5896 10369
rect 5576 10304 5584 10368
rect 5648 10304 5664 10368
rect 5728 10304 5744 10368
rect 5808 10304 5824 10368
rect 5888 10304 5896 10368
rect 5576 10303 5896 10304
rect 14840 10368 15160 10369
rect 14840 10304 14848 10368
rect 14912 10304 14928 10368
rect 14992 10304 15008 10368
rect 15072 10304 15088 10368
rect 15152 10304 15160 10368
rect 14840 10303 15160 10304
rect 24104 10368 24424 10369
rect 24104 10304 24112 10368
rect 24176 10304 24192 10368
rect 24256 10304 24272 10368
rect 24336 10304 24352 10368
rect 24416 10304 24424 10368
rect 24104 10303 24424 10304
rect 25957 10298 26023 10301
rect 29200 10298 30000 10388
rect 25957 10296 30000 10298
rect 25957 10240 25962 10296
rect 26018 10240 30000 10296
rect 25957 10238 30000 10240
rect 25957 10235 26023 10238
rect 29200 10148 30000 10238
rect 10208 9824 10528 9825
rect 10208 9760 10216 9824
rect 10280 9760 10296 9824
rect 10360 9760 10376 9824
rect 10440 9760 10456 9824
rect 10520 9760 10528 9824
rect 10208 9759 10528 9760
rect 19472 9824 19792 9825
rect 19472 9760 19480 9824
rect 19544 9760 19560 9824
rect 19624 9760 19640 9824
rect 19704 9760 19720 9824
rect 19784 9760 19792 9824
rect 19472 9759 19792 9760
rect 0 9468 800 9708
rect 29200 9468 30000 9708
rect 5576 9280 5896 9281
rect 5576 9216 5584 9280
rect 5648 9216 5664 9280
rect 5728 9216 5744 9280
rect 5808 9216 5824 9280
rect 5888 9216 5896 9280
rect 5576 9215 5896 9216
rect 14840 9280 15160 9281
rect 14840 9216 14848 9280
rect 14912 9216 14928 9280
rect 14992 9216 15008 9280
rect 15072 9216 15088 9280
rect 15152 9216 15160 9280
rect 14840 9215 15160 9216
rect 24104 9280 24424 9281
rect 24104 9216 24112 9280
rect 24176 9216 24192 9280
rect 24256 9216 24272 9280
rect 24336 9216 24352 9280
rect 24416 9216 24424 9280
rect 24104 9215 24424 9216
rect 0 8938 800 9028
rect 1853 8938 1919 8941
rect 0 8936 1919 8938
rect 0 8880 1858 8936
rect 1914 8880 1919 8936
rect 0 8878 1919 8880
rect 0 8788 800 8878
rect 1853 8875 1919 8878
rect 26141 8938 26207 8941
rect 29200 8938 30000 9028
rect 26141 8936 30000 8938
rect 26141 8880 26146 8936
rect 26202 8880 30000 8936
rect 26141 8878 30000 8880
rect 26141 8875 26207 8878
rect 29200 8788 30000 8878
rect 10208 8736 10528 8737
rect 10208 8672 10216 8736
rect 10280 8672 10296 8736
rect 10360 8672 10376 8736
rect 10440 8672 10456 8736
rect 10520 8672 10528 8736
rect 10208 8671 10528 8672
rect 19472 8736 19792 8737
rect 19472 8672 19480 8736
rect 19544 8672 19560 8736
rect 19624 8672 19640 8736
rect 19704 8672 19720 8736
rect 19784 8672 19792 8736
rect 19472 8671 19792 8672
rect 0 8258 800 8348
rect 3417 8258 3483 8261
rect 0 8256 3483 8258
rect 0 8200 3422 8256
rect 3478 8200 3483 8256
rect 0 8198 3483 8200
rect 0 8108 800 8198
rect 3417 8195 3483 8198
rect 25957 8258 26023 8261
rect 29200 8258 30000 8348
rect 25957 8256 30000 8258
rect 25957 8200 25962 8256
rect 26018 8200 30000 8256
rect 25957 8198 30000 8200
rect 25957 8195 26023 8198
rect 5576 8192 5896 8193
rect 5576 8128 5584 8192
rect 5648 8128 5664 8192
rect 5728 8128 5744 8192
rect 5808 8128 5824 8192
rect 5888 8128 5896 8192
rect 5576 8127 5896 8128
rect 14840 8192 15160 8193
rect 14840 8128 14848 8192
rect 14912 8128 14928 8192
rect 14992 8128 15008 8192
rect 15072 8128 15088 8192
rect 15152 8128 15160 8192
rect 14840 8127 15160 8128
rect 24104 8192 24424 8193
rect 24104 8128 24112 8192
rect 24176 8128 24192 8192
rect 24256 8128 24272 8192
rect 24336 8128 24352 8192
rect 24416 8128 24424 8192
rect 24104 8127 24424 8128
rect 29200 8108 30000 8198
rect 18689 7988 18755 7989
rect 18638 7986 18644 7988
rect 18598 7926 18644 7986
rect 18708 7984 18755 7988
rect 18750 7928 18755 7984
rect 18638 7924 18644 7926
rect 18708 7924 18755 7928
rect 18689 7923 18755 7924
rect 0 7578 800 7668
rect 10208 7648 10528 7649
rect 10208 7584 10216 7648
rect 10280 7584 10296 7648
rect 10360 7584 10376 7648
rect 10440 7584 10456 7648
rect 10520 7584 10528 7648
rect 10208 7583 10528 7584
rect 19472 7648 19792 7649
rect 19472 7584 19480 7648
rect 19544 7584 19560 7648
rect 19624 7584 19640 7648
rect 19704 7584 19720 7648
rect 19784 7584 19792 7648
rect 19472 7583 19792 7584
rect 2865 7578 2931 7581
rect 0 7576 2931 7578
rect 0 7520 2870 7576
rect 2926 7520 2931 7576
rect 0 7518 2931 7520
rect 0 7428 800 7518
rect 2865 7515 2931 7518
rect 27521 7578 27587 7581
rect 29200 7578 30000 7668
rect 27521 7576 30000 7578
rect 27521 7520 27526 7576
rect 27582 7520 30000 7576
rect 27521 7518 30000 7520
rect 27521 7515 27587 7518
rect 29200 7428 30000 7518
rect 5576 7104 5896 7105
rect 5576 7040 5584 7104
rect 5648 7040 5664 7104
rect 5728 7040 5744 7104
rect 5808 7040 5824 7104
rect 5888 7040 5896 7104
rect 5576 7039 5896 7040
rect 14840 7104 15160 7105
rect 14840 7040 14848 7104
rect 14912 7040 14928 7104
rect 14992 7040 15008 7104
rect 15072 7040 15088 7104
rect 15152 7040 15160 7104
rect 14840 7039 15160 7040
rect 24104 7104 24424 7105
rect 24104 7040 24112 7104
rect 24176 7040 24192 7104
rect 24256 7040 24272 7104
rect 24336 7040 24352 7104
rect 24416 7040 24424 7104
rect 24104 7039 24424 7040
rect 0 6748 800 6988
rect 27521 6898 27587 6901
rect 29200 6898 30000 6988
rect 27521 6896 30000 6898
rect 27521 6840 27526 6896
rect 27582 6840 30000 6896
rect 27521 6838 30000 6840
rect 27521 6835 27587 6838
rect 29200 6748 30000 6838
rect 10208 6560 10528 6561
rect 10208 6496 10216 6560
rect 10280 6496 10296 6560
rect 10360 6496 10376 6560
rect 10440 6496 10456 6560
rect 10520 6496 10528 6560
rect 10208 6495 10528 6496
rect 19472 6560 19792 6561
rect 19472 6496 19480 6560
rect 19544 6496 19560 6560
rect 19624 6496 19640 6560
rect 19704 6496 19720 6560
rect 19784 6496 19792 6560
rect 19472 6495 19792 6496
rect 0 6218 800 6308
rect 3417 6218 3483 6221
rect 0 6216 3483 6218
rect 0 6160 3422 6216
rect 3478 6160 3483 6216
rect 0 6158 3483 6160
rect 0 6068 800 6158
rect 3417 6155 3483 6158
rect 5576 6016 5896 6017
rect 5576 5952 5584 6016
rect 5648 5952 5664 6016
rect 5728 5952 5744 6016
rect 5808 5952 5824 6016
rect 5888 5952 5896 6016
rect 5576 5951 5896 5952
rect 14840 6016 15160 6017
rect 14840 5952 14848 6016
rect 14912 5952 14928 6016
rect 14992 5952 15008 6016
rect 15072 5952 15088 6016
rect 15152 5952 15160 6016
rect 14840 5951 15160 5952
rect 24104 6016 24424 6017
rect 24104 5952 24112 6016
rect 24176 5952 24192 6016
rect 24256 5952 24272 6016
rect 24336 5952 24352 6016
rect 24416 5952 24424 6016
rect 24104 5951 24424 5952
rect 28165 5538 28231 5541
rect 29200 5538 30000 5628
rect 28165 5536 30000 5538
rect 28165 5480 28170 5536
rect 28226 5480 30000 5536
rect 28165 5478 30000 5480
rect 28165 5475 28231 5478
rect 10208 5472 10528 5473
rect 10208 5408 10216 5472
rect 10280 5408 10296 5472
rect 10360 5408 10376 5472
rect 10440 5408 10456 5472
rect 10520 5408 10528 5472
rect 10208 5407 10528 5408
rect 19472 5472 19792 5473
rect 19472 5408 19480 5472
rect 19544 5408 19560 5472
rect 19624 5408 19640 5472
rect 19704 5408 19720 5472
rect 19784 5408 19792 5472
rect 19472 5407 19792 5408
rect 29200 5388 30000 5478
rect 0 4858 800 4948
rect 5576 4928 5896 4929
rect 5576 4864 5584 4928
rect 5648 4864 5664 4928
rect 5728 4864 5744 4928
rect 5808 4864 5824 4928
rect 5888 4864 5896 4928
rect 5576 4863 5896 4864
rect 14840 4928 15160 4929
rect 14840 4864 14848 4928
rect 14912 4864 14928 4928
rect 14992 4864 15008 4928
rect 15072 4864 15088 4928
rect 15152 4864 15160 4928
rect 14840 4863 15160 4864
rect 24104 4928 24424 4929
rect 24104 4864 24112 4928
rect 24176 4864 24192 4928
rect 24256 4864 24272 4928
rect 24336 4864 24352 4928
rect 24416 4864 24424 4928
rect 24104 4863 24424 4864
rect 3325 4858 3391 4861
rect 0 4856 3391 4858
rect 0 4800 3330 4856
rect 3386 4800 3391 4856
rect 0 4798 3391 4800
rect 0 4708 800 4798
rect 3325 4795 3391 4798
rect 29200 4708 30000 4948
rect 10208 4384 10528 4385
rect 10208 4320 10216 4384
rect 10280 4320 10296 4384
rect 10360 4320 10376 4384
rect 10440 4320 10456 4384
rect 10520 4320 10528 4384
rect 10208 4319 10528 4320
rect 19472 4384 19792 4385
rect 19472 4320 19480 4384
rect 19544 4320 19560 4384
rect 19624 4320 19640 4384
rect 19704 4320 19720 4384
rect 19784 4320 19792 4384
rect 19472 4319 19792 4320
rect 0 4178 800 4268
rect 1393 4178 1459 4181
rect 0 4176 1459 4178
rect 0 4120 1398 4176
rect 1454 4120 1459 4176
rect 0 4118 1459 4120
rect 0 4028 800 4118
rect 1393 4115 1459 4118
rect 5257 4042 5323 4045
rect 27286 4042 27292 4044
rect 5257 4040 27292 4042
rect 5257 3984 5262 4040
rect 5318 3984 27292 4040
rect 5257 3982 27292 3984
rect 5257 3979 5323 3982
rect 27286 3980 27292 3982
rect 27356 3980 27362 4044
rect 29200 4028 30000 4268
rect 5576 3840 5896 3841
rect 5576 3776 5584 3840
rect 5648 3776 5664 3840
rect 5728 3776 5744 3840
rect 5808 3776 5824 3840
rect 5888 3776 5896 3840
rect 5576 3775 5896 3776
rect 14840 3840 15160 3841
rect 14840 3776 14848 3840
rect 14912 3776 14928 3840
rect 14992 3776 15008 3840
rect 15072 3776 15088 3840
rect 15152 3776 15160 3840
rect 14840 3775 15160 3776
rect 24104 3840 24424 3841
rect 24104 3776 24112 3840
rect 24176 3776 24192 3840
rect 24256 3776 24272 3840
rect 24336 3776 24352 3840
rect 24416 3776 24424 3840
rect 24104 3775 24424 3776
rect 14641 3634 14707 3637
rect 25037 3634 25103 3637
rect 14641 3632 25103 3634
rect 0 3498 800 3588
rect 14641 3576 14646 3632
rect 14702 3576 25042 3632
rect 25098 3576 25103 3632
rect 14641 3574 25103 3576
rect 14641 3571 14707 3574
rect 25037 3571 25103 3574
rect 3693 3498 3759 3501
rect 0 3496 3759 3498
rect 0 3440 3698 3496
rect 3754 3440 3759 3496
rect 0 3438 3759 3440
rect 0 3348 800 3438
rect 3693 3435 3759 3438
rect 27429 3498 27495 3501
rect 29200 3498 30000 3588
rect 27429 3496 30000 3498
rect 27429 3440 27434 3496
rect 27490 3440 30000 3496
rect 27429 3438 30000 3440
rect 27429 3435 27495 3438
rect 29200 3348 30000 3438
rect 10208 3296 10528 3297
rect 10208 3232 10216 3296
rect 10280 3232 10296 3296
rect 10360 3232 10376 3296
rect 10440 3232 10456 3296
rect 10520 3232 10528 3296
rect 10208 3231 10528 3232
rect 19472 3296 19792 3297
rect 19472 3232 19480 3296
rect 19544 3232 19560 3296
rect 19624 3232 19640 3296
rect 19704 3232 19720 3296
rect 19784 3232 19792 3296
rect 19472 3231 19792 3232
rect 0 2818 800 2908
rect 2773 2818 2839 2821
rect 0 2816 2839 2818
rect 0 2760 2778 2816
rect 2834 2760 2839 2816
rect 0 2758 2839 2760
rect 0 2668 800 2758
rect 2773 2755 2839 2758
rect 25957 2818 26023 2821
rect 29200 2818 30000 2908
rect 25957 2816 30000 2818
rect 25957 2760 25962 2816
rect 26018 2760 30000 2816
rect 25957 2758 30000 2760
rect 25957 2755 26023 2758
rect 5576 2752 5896 2753
rect 5576 2688 5584 2752
rect 5648 2688 5664 2752
rect 5728 2688 5744 2752
rect 5808 2688 5824 2752
rect 5888 2688 5896 2752
rect 5576 2687 5896 2688
rect 14840 2752 15160 2753
rect 14840 2688 14848 2752
rect 14912 2688 14928 2752
rect 14992 2688 15008 2752
rect 15072 2688 15088 2752
rect 15152 2688 15160 2752
rect 14840 2687 15160 2688
rect 24104 2752 24424 2753
rect 24104 2688 24112 2752
rect 24176 2688 24192 2752
rect 24256 2688 24272 2752
rect 24336 2688 24352 2752
rect 24416 2688 24424 2752
rect 24104 2687 24424 2688
rect 29200 2668 30000 2758
rect 0 2138 800 2228
rect 10208 2208 10528 2209
rect 10208 2144 10216 2208
rect 10280 2144 10296 2208
rect 10360 2144 10376 2208
rect 10440 2144 10456 2208
rect 10520 2144 10528 2208
rect 10208 2143 10528 2144
rect 19472 2208 19792 2209
rect 19472 2144 19480 2208
rect 19544 2144 19560 2208
rect 19624 2144 19640 2208
rect 19704 2144 19720 2208
rect 19784 2144 19792 2208
rect 19472 2143 19792 2144
rect 3417 2138 3483 2141
rect 0 2136 3483 2138
rect 0 2080 3422 2136
rect 3478 2080 3483 2136
rect 0 2078 3483 2080
rect 0 1988 800 2078
rect 3417 2075 3483 2078
rect 28993 2138 29059 2141
rect 29200 2138 30000 2228
rect 28993 2136 30000 2138
rect 28993 2080 28998 2136
rect 29054 2080 30000 2136
rect 28993 2078 30000 2080
rect 28993 2075 29059 2078
rect 29200 1988 30000 2078
rect 0 1458 800 1548
rect 3325 1458 3391 1461
rect 0 1456 3391 1458
rect 0 1400 3330 1456
rect 3386 1400 3391 1456
rect 0 1398 3391 1400
rect 0 1308 800 1398
rect 3325 1395 3391 1398
rect 27521 1458 27587 1461
rect 29200 1458 30000 1548
rect 27521 1456 30000 1458
rect 27521 1400 27526 1456
rect 27582 1400 30000 1456
rect 27521 1398 30000 1400
rect 27521 1395 27587 1398
rect 29200 1308 30000 1398
rect 0 628 800 868
rect 29200 -52 30000 188
<< via3 >>
rect 5584 47356 5648 47360
rect 5584 47300 5588 47356
rect 5588 47300 5644 47356
rect 5644 47300 5648 47356
rect 5584 47296 5648 47300
rect 5664 47356 5728 47360
rect 5664 47300 5668 47356
rect 5668 47300 5724 47356
rect 5724 47300 5728 47356
rect 5664 47296 5728 47300
rect 5744 47356 5808 47360
rect 5744 47300 5748 47356
rect 5748 47300 5804 47356
rect 5804 47300 5808 47356
rect 5744 47296 5808 47300
rect 5824 47356 5888 47360
rect 5824 47300 5828 47356
rect 5828 47300 5884 47356
rect 5884 47300 5888 47356
rect 5824 47296 5888 47300
rect 14848 47356 14912 47360
rect 14848 47300 14852 47356
rect 14852 47300 14908 47356
rect 14908 47300 14912 47356
rect 14848 47296 14912 47300
rect 14928 47356 14992 47360
rect 14928 47300 14932 47356
rect 14932 47300 14988 47356
rect 14988 47300 14992 47356
rect 14928 47296 14992 47300
rect 15008 47356 15072 47360
rect 15008 47300 15012 47356
rect 15012 47300 15068 47356
rect 15068 47300 15072 47356
rect 15008 47296 15072 47300
rect 15088 47356 15152 47360
rect 15088 47300 15092 47356
rect 15092 47300 15148 47356
rect 15148 47300 15152 47356
rect 15088 47296 15152 47300
rect 24112 47356 24176 47360
rect 24112 47300 24116 47356
rect 24116 47300 24172 47356
rect 24172 47300 24176 47356
rect 24112 47296 24176 47300
rect 24192 47356 24256 47360
rect 24192 47300 24196 47356
rect 24196 47300 24252 47356
rect 24252 47300 24256 47356
rect 24192 47296 24256 47300
rect 24272 47356 24336 47360
rect 24272 47300 24276 47356
rect 24276 47300 24332 47356
rect 24332 47300 24336 47356
rect 24272 47296 24336 47300
rect 24352 47356 24416 47360
rect 24352 47300 24356 47356
rect 24356 47300 24412 47356
rect 24412 47300 24416 47356
rect 24352 47296 24416 47300
rect 10216 46812 10280 46816
rect 10216 46756 10220 46812
rect 10220 46756 10276 46812
rect 10276 46756 10280 46812
rect 10216 46752 10280 46756
rect 10296 46812 10360 46816
rect 10296 46756 10300 46812
rect 10300 46756 10356 46812
rect 10356 46756 10360 46812
rect 10296 46752 10360 46756
rect 10376 46812 10440 46816
rect 10376 46756 10380 46812
rect 10380 46756 10436 46812
rect 10436 46756 10440 46812
rect 10376 46752 10440 46756
rect 10456 46812 10520 46816
rect 10456 46756 10460 46812
rect 10460 46756 10516 46812
rect 10516 46756 10520 46812
rect 10456 46752 10520 46756
rect 19480 46812 19544 46816
rect 19480 46756 19484 46812
rect 19484 46756 19540 46812
rect 19540 46756 19544 46812
rect 19480 46752 19544 46756
rect 19560 46812 19624 46816
rect 19560 46756 19564 46812
rect 19564 46756 19620 46812
rect 19620 46756 19624 46812
rect 19560 46752 19624 46756
rect 19640 46812 19704 46816
rect 19640 46756 19644 46812
rect 19644 46756 19700 46812
rect 19700 46756 19704 46812
rect 19640 46752 19704 46756
rect 19720 46812 19784 46816
rect 19720 46756 19724 46812
rect 19724 46756 19780 46812
rect 19780 46756 19784 46812
rect 19720 46752 19784 46756
rect 5584 46268 5648 46272
rect 5584 46212 5588 46268
rect 5588 46212 5644 46268
rect 5644 46212 5648 46268
rect 5584 46208 5648 46212
rect 5664 46268 5728 46272
rect 5664 46212 5668 46268
rect 5668 46212 5724 46268
rect 5724 46212 5728 46268
rect 5664 46208 5728 46212
rect 5744 46268 5808 46272
rect 5744 46212 5748 46268
rect 5748 46212 5804 46268
rect 5804 46212 5808 46268
rect 5744 46208 5808 46212
rect 5824 46268 5888 46272
rect 5824 46212 5828 46268
rect 5828 46212 5884 46268
rect 5884 46212 5888 46268
rect 5824 46208 5888 46212
rect 14848 46268 14912 46272
rect 14848 46212 14852 46268
rect 14852 46212 14908 46268
rect 14908 46212 14912 46268
rect 14848 46208 14912 46212
rect 14928 46268 14992 46272
rect 14928 46212 14932 46268
rect 14932 46212 14988 46268
rect 14988 46212 14992 46268
rect 14928 46208 14992 46212
rect 15008 46268 15072 46272
rect 15008 46212 15012 46268
rect 15012 46212 15068 46268
rect 15068 46212 15072 46268
rect 15008 46208 15072 46212
rect 15088 46268 15152 46272
rect 15088 46212 15092 46268
rect 15092 46212 15148 46268
rect 15148 46212 15152 46268
rect 15088 46208 15152 46212
rect 24112 46268 24176 46272
rect 24112 46212 24116 46268
rect 24116 46212 24172 46268
rect 24172 46212 24176 46268
rect 24112 46208 24176 46212
rect 24192 46268 24256 46272
rect 24192 46212 24196 46268
rect 24196 46212 24252 46268
rect 24252 46212 24256 46268
rect 24192 46208 24256 46212
rect 24272 46268 24336 46272
rect 24272 46212 24276 46268
rect 24276 46212 24332 46268
rect 24332 46212 24336 46268
rect 24272 46208 24336 46212
rect 24352 46268 24416 46272
rect 24352 46212 24356 46268
rect 24356 46212 24412 46268
rect 24412 46212 24416 46268
rect 24352 46208 24416 46212
rect 10216 45724 10280 45728
rect 10216 45668 10220 45724
rect 10220 45668 10276 45724
rect 10276 45668 10280 45724
rect 10216 45664 10280 45668
rect 10296 45724 10360 45728
rect 10296 45668 10300 45724
rect 10300 45668 10356 45724
rect 10356 45668 10360 45724
rect 10296 45664 10360 45668
rect 10376 45724 10440 45728
rect 10376 45668 10380 45724
rect 10380 45668 10436 45724
rect 10436 45668 10440 45724
rect 10376 45664 10440 45668
rect 10456 45724 10520 45728
rect 10456 45668 10460 45724
rect 10460 45668 10516 45724
rect 10516 45668 10520 45724
rect 10456 45664 10520 45668
rect 19480 45724 19544 45728
rect 19480 45668 19484 45724
rect 19484 45668 19540 45724
rect 19540 45668 19544 45724
rect 19480 45664 19544 45668
rect 19560 45724 19624 45728
rect 19560 45668 19564 45724
rect 19564 45668 19620 45724
rect 19620 45668 19624 45724
rect 19560 45664 19624 45668
rect 19640 45724 19704 45728
rect 19640 45668 19644 45724
rect 19644 45668 19700 45724
rect 19700 45668 19704 45724
rect 19640 45664 19704 45668
rect 19720 45724 19784 45728
rect 19720 45668 19724 45724
rect 19724 45668 19780 45724
rect 19780 45668 19784 45724
rect 19720 45664 19784 45668
rect 5584 45180 5648 45184
rect 5584 45124 5588 45180
rect 5588 45124 5644 45180
rect 5644 45124 5648 45180
rect 5584 45120 5648 45124
rect 5664 45180 5728 45184
rect 5664 45124 5668 45180
rect 5668 45124 5724 45180
rect 5724 45124 5728 45180
rect 5664 45120 5728 45124
rect 5744 45180 5808 45184
rect 5744 45124 5748 45180
rect 5748 45124 5804 45180
rect 5804 45124 5808 45180
rect 5744 45120 5808 45124
rect 5824 45180 5888 45184
rect 5824 45124 5828 45180
rect 5828 45124 5884 45180
rect 5884 45124 5888 45180
rect 5824 45120 5888 45124
rect 14848 45180 14912 45184
rect 14848 45124 14852 45180
rect 14852 45124 14908 45180
rect 14908 45124 14912 45180
rect 14848 45120 14912 45124
rect 14928 45180 14992 45184
rect 14928 45124 14932 45180
rect 14932 45124 14988 45180
rect 14988 45124 14992 45180
rect 14928 45120 14992 45124
rect 15008 45180 15072 45184
rect 15008 45124 15012 45180
rect 15012 45124 15068 45180
rect 15068 45124 15072 45180
rect 15008 45120 15072 45124
rect 15088 45180 15152 45184
rect 15088 45124 15092 45180
rect 15092 45124 15148 45180
rect 15148 45124 15152 45180
rect 15088 45120 15152 45124
rect 24112 45180 24176 45184
rect 24112 45124 24116 45180
rect 24116 45124 24172 45180
rect 24172 45124 24176 45180
rect 24112 45120 24176 45124
rect 24192 45180 24256 45184
rect 24192 45124 24196 45180
rect 24196 45124 24252 45180
rect 24252 45124 24256 45180
rect 24192 45120 24256 45124
rect 24272 45180 24336 45184
rect 24272 45124 24276 45180
rect 24276 45124 24332 45180
rect 24332 45124 24336 45180
rect 24272 45120 24336 45124
rect 24352 45180 24416 45184
rect 24352 45124 24356 45180
rect 24356 45124 24412 45180
rect 24412 45124 24416 45180
rect 24352 45120 24416 45124
rect 10216 44636 10280 44640
rect 10216 44580 10220 44636
rect 10220 44580 10276 44636
rect 10276 44580 10280 44636
rect 10216 44576 10280 44580
rect 10296 44636 10360 44640
rect 10296 44580 10300 44636
rect 10300 44580 10356 44636
rect 10356 44580 10360 44636
rect 10296 44576 10360 44580
rect 10376 44636 10440 44640
rect 10376 44580 10380 44636
rect 10380 44580 10436 44636
rect 10436 44580 10440 44636
rect 10376 44576 10440 44580
rect 10456 44636 10520 44640
rect 10456 44580 10460 44636
rect 10460 44580 10516 44636
rect 10516 44580 10520 44636
rect 10456 44576 10520 44580
rect 19480 44636 19544 44640
rect 19480 44580 19484 44636
rect 19484 44580 19540 44636
rect 19540 44580 19544 44636
rect 19480 44576 19544 44580
rect 19560 44636 19624 44640
rect 19560 44580 19564 44636
rect 19564 44580 19620 44636
rect 19620 44580 19624 44636
rect 19560 44576 19624 44580
rect 19640 44636 19704 44640
rect 19640 44580 19644 44636
rect 19644 44580 19700 44636
rect 19700 44580 19704 44636
rect 19640 44576 19704 44580
rect 19720 44636 19784 44640
rect 19720 44580 19724 44636
rect 19724 44580 19780 44636
rect 19780 44580 19784 44636
rect 19720 44576 19784 44580
rect 21956 44296 22020 44300
rect 21956 44240 22006 44296
rect 22006 44240 22020 44296
rect 21956 44236 22020 44240
rect 5584 44092 5648 44096
rect 5584 44036 5588 44092
rect 5588 44036 5644 44092
rect 5644 44036 5648 44092
rect 5584 44032 5648 44036
rect 5664 44092 5728 44096
rect 5664 44036 5668 44092
rect 5668 44036 5724 44092
rect 5724 44036 5728 44092
rect 5664 44032 5728 44036
rect 5744 44092 5808 44096
rect 5744 44036 5748 44092
rect 5748 44036 5804 44092
rect 5804 44036 5808 44092
rect 5744 44032 5808 44036
rect 5824 44092 5888 44096
rect 5824 44036 5828 44092
rect 5828 44036 5884 44092
rect 5884 44036 5888 44092
rect 5824 44032 5888 44036
rect 14848 44092 14912 44096
rect 14848 44036 14852 44092
rect 14852 44036 14908 44092
rect 14908 44036 14912 44092
rect 14848 44032 14912 44036
rect 14928 44092 14992 44096
rect 14928 44036 14932 44092
rect 14932 44036 14988 44092
rect 14988 44036 14992 44092
rect 14928 44032 14992 44036
rect 15008 44092 15072 44096
rect 15008 44036 15012 44092
rect 15012 44036 15068 44092
rect 15068 44036 15072 44092
rect 15008 44032 15072 44036
rect 15088 44092 15152 44096
rect 15088 44036 15092 44092
rect 15092 44036 15148 44092
rect 15148 44036 15152 44092
rect 15088 44032 15152 44036
rect 24112 44092 24176 44096
rect 24112 44036 24116 44092
rect 24116 44036 24172 44092
rect 24172 44036 24176 44092
rect 24112 44032 24176 44036
rect 24192 44092 24256 44096
rect 24192 44036 24196 44092
rect 24196 44036 24252 44092
rect 24252 44036 24256 44092
rect 24192 44032 24256 44036
rect 24272 44092 24336 44096
rect 24272 44036 24276 44092
rect 24276 44036 24332 44092
rect 24332 44036 24336 44092
rect 24272 44032 24336 44036
rect 24352 44092 24416 44096
rect 24352 44036 24356 44092
rect 24356 44036 24412 44092
rect 24412 44036 24416 44092
rect 24352 44032 24416 44036
rect 10216 43548 10280 43552
rect 10216 43492 10220 43548
rect 10220 43492 10276 43548
rect 10276 43492 10280 43548
rect 10216 43488 10280 43492
rect 10296 43548 10360 43552
rect 10296 43492 10300 43548
rect 10300 43492 10356 43548
rect 10356 43492 10360 43548
rect 10296 43488 10360 43492
rect 10376 43548 10440 43552
rect 10376 43492 10380 43548
rect 10380 43492 10436 43548
rect 10436 43492 10440 43548
rect 10376 43488 10440 43492
rect 10456 43548 10520 43552
rect 10456 43492 10460 43548
rect 10460 43492 10516 43548
rect 10516 43492 10520 43548
rect 10456 43488 10520 43492
rect 19480 43548 19544 43552
rect 19480 43492 19484 43548
rect 19484 43492 19540 43548
rect 19540 43492 19544 43548
rect 19480 43488 19544 43492
rect 19560 43548 19624 43552
rect 19560 43492 19564 43548
rect 19564 43492 19620 43548
rect 19620 43492 19624 43548
rect 19560 43488 19624 43492
rect 19640 43548 19704 43552
rect 19640 43492 19644 43548
rect 19644 43492 19700 43548
rect 19700 43492 19704 43548
rect 19640 43488 19704 43492
rect 19720 43548 19784 43552
rect 19720 43492 19724 43548
rect 19724 43492 19780 43548
rect 19780 43492 19784 43548
rect 19720 43488 19784 43492
rect 5584 43004 5648 43008
rect 5584 42948 5588 43004
rect 5588 42948 5644 43004
rect 5644 42948 5648 43004
rect 5584 42944 5648 42948
rect 5664 43004 5728 43008
rect 5664 42948 5668 43004
rect 5668 42948 5724 43004
rect 5724 42948 5728 43004
rect 5664 42944 5728 42948
rect 5744 43004 5808 43008
rect 5744 42948 5748 43004
rect 5748 42948 5804 43004
rect 5804 42948 5808 43004
rect 5744 42944 5808 42948
rect 5824 43004 5888 43008
rect 5824 42948 5828 43004
rect 5828 42948 5884 43004
rect 5884 42948 5888 43004
rect 5824 42944 5888 42948
rect 14848 43004 14912 43008
rect 14848 42948 14852 43004
rect 14852 42948 14908 43004
rect 14908 42948 14912 43004
rect 14848 42944 14912 42948
rect 14928 43004 14992 43008
rect 14928 42948 14932 43004
rect 14932 42948 14988 43004
rect 14988 42948 14992 43004
rect 14928 42944 14992 42948
rect 15008 43004 15072 43008
rect 15008 42948 15012 43004
rect 15012 42948 15068 43004
rect 15068 42948 15072 43004
rect 15008 42944 15072 42948
rect 15088 43004 15152 43008
rect 15088 42948 15092 43004
rect 15092 42948 15148 43004
rect 15148 42948 15152 43004
rect 15088 42944 15152 42948
rect 24112 43004 24176 43008
rect 24112 42948 24116 43004
rect 24116 42948 24172 43004
rect 24172 42948 24176 43004
rect 24112 42944 24176 42948
rect 24192 43004 24256 43008
rect 24192 42948 24196 43004
rect 24196 42948 24252 43004
rect 24252 42948 24256 43004
rect 24192 42944 24256 42948
rect 24272 43004 24336 43008
rect 24272 42948 24276 43004
rect 24276 42948 24332 43004
rect 24332 42948 24336 43004
rect 24272 42944 24336 42948
rect 24352 43004 24416 43008
rect 24352 42948 24356 43004
rect 24356 42948 24412 43004
rect 24412 42948 24416 43004
rect 24352 42944 24416 42948
rect 10216 42460 10280 42464
rect 10216 42404 10220 42460
rect 10220 42404 10276 42460
rect 10276 42404 10280 42460
rect 10216 42400 10280 42404
rect 10296 42460 10360 42464
rect 10296 42404 10300 42460
rect 10300 42404 10356 42460
rect 10356 42404 10360 42460
rect 10296 42400 10360 42404
rect 10376 42460 10440 42464
rect 10376 42404 10380 42460
rect 10380 42404 10436 42460
rect 10436 42404 10440 42460
rect 10376 42400 10440 42404
rect 10456 42460 10520 42464
rect 10456 42404 10460 42460
rect 10460 42404 10516 42460
rect 10516 42404 10520 42460
rect 10456 42400 10520 42404
rect 19480 42460 19544 42464
rect 19480 42404 19484 42460
rect 19484 42404 19540 42460
rect 19540 42404 19544 42460
rect 19480 42400 19544 42404
rect 19560 42460 19624 42464
rect 19560 42404 19564 42460
rect 19564 42404 19620 42460
rect 19620 42404 19624 42460
rect 19560 42400 19624 42404
rect 19640 42460 19704 42464
rect 19640 42404 19644 42460
rect 19644 42404 19700 42460
rect 19700 42404 19704 42460
rect 19640 42400 19704 42404
rect 19720 42460 19784 42464
rect 19720 42404 19724 42460
rect 19724 42404 19780 42460
rect 19780 42404 19784 42460
rect 19720 42400 19784 42404
rect 5584 41916 5648 41920
rect 5584 41860 5588 41916
rect 5588 41860 5644 41916
rect 5644 41860 5648 41916
rect 5584 41856 5648 41860
rect 5664 41916 5728 41920
rect 5664 41860 5668 41916
rect 5668 41860 5724 41916
rect 5724 41860 5728 41916
rect 5664 41856 5728 41860
rect 5744 41916 5808 41920
rect 5744 41860 5748 41916
rect 5748 41860 5804 41916
rect 5804 41860 5808 41916
rect 5744 41856 5808 41860
rect 5824 41916 5888 41920
rect 5824 41860 5828 41916
rect 5828 41860 5884 41916
rect 5884 41860 5888 41916
rect 5824 41856 5888 41860
rect 14848 41916 14912 41920
rect 14848 41860 14852 41916
rect 14852 41860 14908 41916
rect 14908 41860 14912 41916
rect 14848 41856 14912 41860
rect 14928 41916 14992 41920
rect 14928 41860 14932 41916
rect 14932 41860 14988 41916
rect 14988 41860 14992 41916
rect 14928 41856 14992 41860
rect 15008 41916 15072 41920
rect 15008 41860 15012 41916
rect 15012 41860 15068 41916
rect 15068 41860 15072 41916
rect 15008 41856 15072 41860
rect 15088 41916 15152 41920
rect 15088 41860 15092 41916
rect 15092 41860 15148 41916
rect 15148 41860 15152 41916
rect 15088 41856 15152 41860
rect 24112 41916 24176 41920
rect 24112 41860 24116 41916
rect 24116 41860 24172 41916
rect 24172 41860 24176 41916
rect 24112 41856 24176 41860
rect 24192 41916 24256 41920
rect 24192 41860 24196 41916
rect 24196 41860 24252 41916
rect 24252 41860 24256 41916
rect 24192 41856 24256 41860
rect 24272 41916 24336 41920
rect 24272 41860 24276 41916
rect 24276 41860 24332 41916
rect 24332 41860 24336 41916
rect 24272 41856 24336 41860
rect 24352 41916 24416 41920
rect 24352 41860 24356 41916
rect 24356 41860 24412 41916
rect 24412 41860 24416 41916
rect 24352 41856 24416 41860
rect 10216 41372 10280 41376
rect 10216 41316 10220 41372
rect 10220 41316 10276 41372
rect 10276 41316 10280 41372
rect 10216 41312 10280 41316
rect 10296 41372 10360 41376
rect 10296 41316 10300 41372
rect 10300 41316 10356 41372
rect 10356 41316 10360 41372
rect 10296 41312 10360 41316
rect 10376 41372 10440 41376
rect 10376 41316 10380 41372
rect 10380 41316 10436 41372
rect 10436 41316 10440 41372
rect 10376 41312 10440 41316
rect 10456 41372 10520 41376
rect 10456 41316 10460 41372
rect 10460 41316 10516 41372
rect 10516 41316 10520 41372
rect 10456 41312 10520 41316
rect 19480 41372 19544 41376
rect 19480 41316 19484 41372
rect 19484 41316 19540 41372
rect 19540 41316 19544 41372
rect 19480 41312 19544 41316
rect 19560 41372 19624 41376
rect 19560 41316 19564 41372
rect 19564 41316 19620 41372
rect 19620 41316 19624 41372
rect 19560 41312 19624 41316
rect 19640 41372 19704 41376
rect 19640 41316 19644 41372
rect 19644 41316 19700 41372
rect 19700 41316 19704 41372
rect 19640 41312 19704 41316
rect 19720 41372 19784 41376
rect 19720 41316 19724 41372
rect 19724 41316 19780 41372
rect 19780 41316 19784 41372
rect 19720 41312 19784 41316
rect 5584 40828 5648 40832
rect 5584 40772 5588 40828
rect 5588 40772 5644 40828
rect 5644 40772 5648 40828
rect 5584 40768 5648 40772
rect 5664 40828 5728 40832
rect 5664 40772 5668 40828
rect 5668 40772 5724 40828
rect 5724 40772 5728 40828
rect 5664 40768 5728 40772
rect 5744 40828 5808 40832
rect 5744 40772 5748 40828
rect 5748 40772 5804 40828
rect 5804 40772 5808 40828
rect 5744 40768 5808 40772
rect 5824 40828 5888 40832
rect 5824 40772 5828 40828
rect 5828 40772 5884 40828
rect 5884 40772 5888 40828
rect 5824 40768 5888 40772
rect 14848 40828 14912 40832
rect 14848 40772 14852 40828
rect 14852 40772 14908 40828
rect 14908 40772 14912 40828
rect 14848 40768 14912 40772
rect 14928 40828 14992 40832
rect 14928 40772 14932 40828
rect 14932 40772 14988 40828
rect 14988 40772 14992 40828
rect 14928 40768 14992 40772
rect 15008 40828 15072 40832
rect 15008 40772 15012 40828
rect 15012 40772 15068 40828
rect 15068 40772 15072 40828
rect 15008 40768 15072 40772
rect 15088 40828 15152 40832
rect 15088 40772 15092 40828
rect 15092 40772 15148 40828
rect 15148 40772 15152 40828
rect 15088 40768 15152 40772
rect 24112 40828 24176 40832
rect 24112 40772 24116 40828
rect 24116 40772 24172 40828
rect 24172 40772 24176 40828
rect 24112 40768 24176 40772
rect 24192 40828 24256 40832
rect 24192 40772 24196 40828
rect 24196 40772 24252 40828
rect 24252 40772 24256 40828
rect 24192 40768 24256 40772
rect 24272 40828 24336 40832
rect 24272 40772 24276 40828
rect 24276 40772 24332 40828
rect 24332 40772 24336 40828
rect 24272 40768 24336 40772
rect 24352 40828 24416 40832
rect 24352 40772 24356 40828
rect 24356 40772 24412 40828
rect 24412 40772 24416 40828
rect 24352 40768 24416 40772
rect 10216 40284 10280 40288
rect 10216 40228 10220 40284
rect 10220 40228 10276 40284
rect 10276 40228 10280 40284
rect 10216 40224 10280 40228
rect 10296 40284 10360 40288
rect 10296 40228 10300 40284
rect 10300 40228 10356 40284
rect 10356 40228 10360 40284
rect 10296 40224 10360 40228
rect 10376 40284 10440 40288
rect 10376 40228 10380 40284
rect 10380 40228 10436 40284
rect 10436 40228 10440 40284
rect 10376 40224 10440 40228
rect 10456 40284 10520 40288
rect 10456 40228 10460 40284
rect 10460 40228 10516 40284
rect 10516 40228 10520 40284
rect 10456 40224 10520 40228
rect 19480 40284 19544 40288
rect 19480 40228 19484 40284
rect 19484 40228 19540 40284
rect 19540 40228 19544 40284
rect 19480 40224 19544 40228
rect 19560 40284 19624 40288
rect 19560 40228 19564 40284
rect 19564 40228 19620 40284
rect 19620 40228 19624 40284
rect 19560 40224 19624 40228
rect 19640 40284 19704 40288
rect 19640 40228 19644 40284
rect 19644 40228 19700 40284
rect 19700 40228 19704 40284
rect 19640 40224 19704 40228
rect 19720 40284 19784 40288
rect 19720 40228 19724 40284
rect 19724 40228 19780 40284
rect 19780 40228 19784 40284
rect 19720 40224 19784 40228
rect 5584 39740 5648 39744
rect 5584 39684 5588 39740
rect 5588 39684 5644 39740
rect 5644 39684 5648 39740
rect 5584 39680 5648 39684
rect 5664 39740 5728 39744
rect 5664 39684 5668 39740
rect 5668 39684 5724 39740
rect 5724 39684 5728 39740
rect 5664 39680 5728 39684
rect 5744 39740 5808 39744
rect 5744 39684 5748 39740
rect 5748 39684 5804 39740
rect 5804 39684 5808 39740
rect 5744 39680 5808 39684
rect 5824 39740 5888 39744
rect 5824 39684 5828 39740
rect 5828 39684 5884 39740
rect 5884 39684 5888 39740
rect 5824 39680 5888 39684
rect 14848 39740 14912 39744
rect 14848 39684 14852 39740
rect 14852 39684 14908 39740
rect 14908 39684 14912 39740
rect 14848 39680 14912 39684
rect 14928 39740 14992 39744
rect 14928 39684 14932 39740
rect 14932 39684 14988 39740
rect 14988 39684 14992 39740
rect 14928 39680 14992 39684
rect 15008 39740 15072 39744
rect 15008 39684 15012 39740
rect 15012 39684 15068 39740
rect 15068 39684 15072 39740
rect 15008 39680 15072 39684
rect 15088 39740 15152 39744
rect 15088 39684 15092 39740
rect 15092 39684 15148 39740
rect 15148 39684 15152 39740
rect 15088 39680 15152 39684
rect 24112 39740 24176 39744
rect 24112 39684 24116 39740
rect 24116 39684 24172 39740
rect 24172 39684 24176 39740
rect 24112 39680 24176 39684
rect 24192 39740 24256 39744
rect 24192 39684 24196 39740
rect 24196 39684 24252 39740
rect 24252 39684 24256 39740
rect 24192 39680 24256 39684
rect 24272 39740 24336 39744
rect 24272 39684 24276 39740
rect 24276 39684 24332 39740
rect 24332 39684 24336 39740
rect 24272 39680 24336 39684
rect 24352 39740 24416 39744
rect 24352 39684 24356 39740
rect 24356 39684 24412 39740
rect 24412 39684 24416 39740
rect 24352 39680 24416 39684
rect 10216 39196 10280 39200
rect 10216 39140 10220 39196
rect 10220 39140 10276 39196
rect 10276 39140 10280 39196
rect 10216 39136 10280 39140
rect 10296 39196 10360 39200
rect 10296 39140 10300 39196
rect 10300 39140 10356 39196
rect 10356 39140 10360 39196
rect 10296 39136 10360 39140
rect 10376 39196 10440 39200
rect 10376 39140 10380 39196
rect 10380 39140 10436 39196
rect 10436 39140 10440 39196
rect 10376 39136 10440 39140
rect 10456 39196 10520 39200
rect 10456 39140 10460 39196
rect 10460 39140 10516 39196
rect 10516 39140 10520 39196
rect 10456 39136 10520 39140
rect 19480 39196 19544 39200
rect 19480 39140 19484 39196
rect 19484 39140 19540 39196
rect 19540 39140 19544 39196
rect 19480 39136 19544 39140
rect 19560 39196 19624 39200
rect 19560 39140 19564 39196
rect 19564 39140 19620 39196
rect 19620 39140 19624 39196
rect 19560 39136 19624 39140
rect 19640 39196 19704 39200
rect 19640 39140 19644 39196
rect 19644 39140 19700 39196
rect 19700 39140 19704 39196
rect 19640 39136 19704 39140
rect 19720 39196 19784 39200
rect 19720 39140 19724 39196
rect 19724 39140 19780 39196
rect 19780 39140 19784 39196
rect 19720 39136 19784 39140
rect 5584 38652 5648 38656
rect 5584 38596 5588 38652
rect 5588 38596 5644 38652
rect 5644 38596 5648 38652
rect 5584 38592 5648 38596
rect 5664 38652 5728 38656
rect 5664 38596 5668 38652
rect 5668 38596 5724 38652
rect 5724 38596 5728 38652
rect 5664 38592 5728 38596
rect 5744 38652 5808 38656
rect 5744 38596 5748 38652
rect 5748 38596 5804 38652
rect 5804 38596 5808 38652
rect 5744 38592 5808 38596
rect 5824 38652 5888 38656
rect 5824 38596 5828 38652
rect 5828 38596 5884 38652
rect 5884 38596 5888 38652
rect 5824 38592 5888 38596
rect 14848 38652 14912 38656
rect 14848 38596 14852 38652
rect 14852 38596 14908 38652
rect 14908 38596 14912 38652
rect 14848 38592 14912 38596
rect 14928 38652 14992 38656
rect 14928 38596 14932 38652
rect 14932 38596 14988 38652
rect 14988 38596 14992 38652
rect 14928 38592 14992 38596
rect 15008 38652 15072 38656
rect 15008 38596 15012 38652
rect 15012 38596 15068 38652
rect 15068 38596 15072 38652
rect 15008 38592 15072 38596
rect 15088 38652 15152 38656
rect 15088 38596 15092 38652
rect 15092 38596 15148 38652
rect 15148 38596 15152 38652
rect 15088 38592 15152 38596
rect 24112 38652 24176 38656
rect 24112 38596 24116 38652
rect 24116 38596 24172 38652
rect 24172 38596 24176 38652
rect 24112 38592 24176 38596
rect 24192 38652 24256 38656
rect 24192 38596 24196 38652
rect 24196 38596 24252 38652
rect 24252 38596 24256 38652
rect 24192 38592 24256 38596
rect 24272 38652 24336 38656
rect 24272 38596 24276 38652
rect 24276 38596 24332 38652
rect 24332 38596 24336 38652
rect 24272 38592 24336 38596
rect 24352 38652 24416 38656
rect 24352 38596 24356 38652
rect 24356 38596 24412 38652
rect 24412 38596 24416 38652
rect 24352 38592 24416 38596
rect 10216 38108 10280 38112
rect 10216 38052 10220 38108
rect 10220 38052 10276 38108
rect 10276 38052 10280 38108
rect 10216 38048 10280 38052
rect 10296 38108 10360 38112
rect 10296 38052 10300 38108
rect 10300 38052 10356 38108
rect 10356 38052 10360 38108
rect 10296 38048 10360 38052
rect 10376 38108 10440 38112
rect 10376 38052 10380 38108
rect 10380 38052 10436 38108
rect 10436 38052 10440 38108
rect 10376 38048 10440 38052
rect 10456 38108 10520 38112
rect 10456 38052 10460 38108
rect 10460 38052 10516 38108
rect 10516 38052 10520 38108
rect 10456 38048 10520 38052
rect 19480 38108 19544 38112
rect 19480 38052 19484 38108
rect 19484 38052 19540 38108
rect 19540 38052 19544 38108
rect 19480 38048 19544 38052
rect 19560 38108 19624 38112
rect 19560 38052 19564 38108
rect 19564 38052 19620 38108
rect 19620 38052 19624 38108
rect 19560 38048 19624 38052
rect 19640 38108 19704 38112
rect 19640 38052 19644 38108
rect 19644 38052 19700 38108
rect 19700 38052 19704 38108
rect 19640 38048 19704 38052
rect 19720 38108 19784 38112
rect 19720 38052 19724 38108
rect 19724 38052 19780 38108
rect 19780 38052 19784 38108
rect 19720 38048 19784 38052
rect 5584 37564 5648 37568
rect 5584 37508 5588 37564
rect 5588 37508 5644 37564
rect 5644 37508 5648 37564
rect 5584 37504 5648 37508
rect 5664 37564 5728 37568
rect 5664 37508 5668 37564
rect 5668 37508 5724 37564
rect 5724 37508 5728 37564
rect 5664 37504 5728 37508
rect 5744 37564 5808 37568
rect 5744 37508 5748 37564
rect 5748 37508 5804 37564
rect 5804 37508 5808 37564
rect 5744 37504 5808 37508
rect 5824 37564 5888 37568
rect 5824 37508 5828 37564
rect 5828 37508 5884 37564
rect 5884 37508 5888 37564
rect 5824 37504 5888 37508
rect 14848 37564 14912 37568
rect 14848 37508 14852 37564
rect 14852 37508 14908 37564
rect 14908 37508 14912 37564
rect 14848 37504 14912 37508
rect 14928 37564 14992 37568
rect 14928 37508 14932 37564
rect 14932 37508 14988 37564
rect 14988 37508 14992 37564
rect 14928 37504 14992 37508
rect 15008 37564 15072 37568
rect 15008 37508 15012 37564
rect 15012 37508 15068 37564
rect 15068 37508 15072 37564
rect 15008 37504 15072 37508
rect 15088 37564 15152 37568
rect 15088 37508 15092 37564
rect 15092 37508 15148 37564
rect 15148 37508 15152 37564
rect 15088 37504 15152 37508
rect 24112 37564 24176 37568
rect 24112 37508 24116 37564
rect 24116 37508 24172 37564
rect 24172 37508 24176 37564
rect 24112 37504 24176 37508
rect 24192 37564 24256 37568
rect 24192 37508 24196 37564
rect 24196 37508 24252 37564
rect 24252 37508 24256 37564
rect 24192 37504 24256 37508
rect 24272 37564 24336 37568
rect 24272 37508 24276 37564
rect 24276 37508 24332 37564
rect 24332 37508 24336 37564
rect 24272 37504 24336 37508
rect 24352 37564 24416 37568
rect 24352 37508 24356 37564
rect 24356 37508 24412 37564
rect 24412 37508 24416 37564
rect 24352 37504 24416 37508
rect 10216 37020 10280 37024
rect 10216 36964 10220 37020
rect 10220 36964 10276 37020
rect 10276 36964 10280 37020
rect 10216 36960 10280 36964
rect 10296 37020 10360 37024
rect 10296 36964 10300 37020
rect 10300 36964 10356 37020
rect 10356 36964 10360 37020
rect 10296 36960 10360 36964
rect 10376 37020 10440 37024
rect 10376 36964 10380 37020
rect 10380 36964 10436 37020
rect 10436 36964 10440 37020
rect 10376 36960 10440 36964
rect 10456 37020 10520 37024
rect 10456 36964 10460 37020
rect 10460 36964 10516 37020
rect 10516 36964 10520 37020
rect 10456 36960 10520 36964
rect 19480 37020 19544 37024
rect 19480 36964 19484 37020
rect 19484 36964 19540 37020
rect 19540 36964 19544 37020
rect 19480 36960 19544 36964
rect 19560 37020 19624 37024
rect 19560 36964 19564 37020
rect 19564 36964 19620 37020
rect 19620 36964 19624 37020
rect 19560 36960 19624 36964
rect 19640 37020 19704 37024
rect 19640 36964 19644 37020
rect 19644 36964 19700 37020
rect 19700 36964 19704 37020
rect 19640 36960 19704 36964
rect 19720 37020 19784 37024
rect 19720 36964 19724 37020
rect 19724 36964 19780 37020
rect 19780 36964 19784 37020
rect 19720 36960 19784 36964
rect 5584 36476 5648 36480
rect 5584 36420 5588 36476
rect 5588 36420 5644 36476
rect 5644 36420 5648 36476
rect 5584 36416 5648 36420
rect 5664 36476 5728 36480
rect 5664 36420 5668 36476
rect 5668 36420 5724 36476
rect 5724 36420 5728 36476
rect 5664 36416 5728 36420
rect 5744 36476 5808 36480
rect 5744 36420 5748 36476
rect 5748 36420 5804 36476
rect 5804 36420 5808 36476
rect 5744 36416 5808 36420
rect 5824 36476 5888 36480
rect 5824 36420 5828 36476
rect 5828 36420 5884 36476
rect 5884 36420 5888 36476
rect 5824 36416 5888 36420
rect 14848 36476 14912 36480
rect 14848 36420 14852 36476
rect 14852 36420 14908 36476
rect 14908 36420 14912 36476
rect 14848 36416 14912 36420
rect 14928 36476 14992 36480
rect 14928 36420 14932 36476
rect 14932 36420 14988 36476
rect 14988 36420 14992 36476
rect 14928 36416 14992 36420
rect 15008 36476 15072 36480
rect 15008 36420 15012 36476
rect 15012 36420 15068 36476
rect 15068 36420 15072 36476
rect 15008 36416 15072 36420
rect 15088 36476 15152 36480
rect 15088 36420 15092 36476
rect 15092 36420 15148 36476
rect 15148 36420 15152 36476
rect 15088 36416 15152 36420
rect 24112 36476 24176 36480
rect 24112 36420 24116 36476
rect 24116 36420 24172 36476
rect 24172 36420 24176 36476
rect 24112 36416 24176 36420
rect 24192 36476 24256 36480
rect 24192 36420 24196 36476
rect 24196 36420 24252 36476
rect 24252 36420 24256 36476
rect 24192 36416 24256 36420
rect 24272 36476 24336 36480
rect 24272 36420 24276 36476
rect 24276 36420 24332 36476
rect 24332 36420 24336 36476
rect 24272 36416 24336 36420
rect 24352 36476 24416 36480
rect 24352 36420 24356 36476
rect 24356 36420 24412 36476
rect 24412 36420 24416 36476
rect 24352 36416 24416 36420
rect 10216 35932 10280 35936
rect 10216 35876 10220 35932
rect 10220 35876 10276 35932
rect 10276 35876 10280 35932
rect 10216 35872 10280 35876
rect 10296 35932 10360 35936
rect 10296 35876 10300 35932
rect 10300 35876 10356 35932
rect 10356 35876 10360 35932
rect 10296 35872 10360 35876
rect 10376 35932 10440 35936
rect 10376 35876 10380 35932
rect 10380 35876 10436 35932
rect 10436 35876 10440 35932
rect 10376 35872 10440 35876
rect 10456 35932 10520 35936
rect 10456 35876 10460 35932
rect 10460 35876 10516 35932
rect 10516 35876 10520 35932
rect 10456 35872 10520 35876
rect 19480 35932 19544 35936
rect 19480 35876 19484 35932
rect 19484 35876 19540 35932
rect 19540 35876 19544 35932
rect 19480 35872 19544 35876
rect 19560 35932 19624 35936
rect 19560 35876 19564 35932
rect 19564 35876 19620 35932
rect 19620 35876 19624 35932
rect 19560 35872 19624 35876
rect 19640 35932 19704 35936
rect 19640 35876 19644 35932
rect 19644 35876 19700 35932
rect 19700 35876 19704 35932
rect 19640 35872 19704 35876
rect 19720 35932 19784 35936
rect 19720 35876 19724 35932
rect 19724 35876 19780 35932
rect 19780 35876 19784 35932
rect 19720 35872 19784 35876
rect 5584 35388 5648 35392
rect 5584 35332 5588 35388
rect 5588 35332 5644 35388
rect 5644 35332 5648 35388
rect 5584 35328 5648 35332
rect 5664 35388 5728 35392
rect 5664 35332 5668 35388
rect 5668 35332 5724 35388
rect 5724 35332 5728 35388
rect 5664 35328 5728 35332
rect 5744 35388 5808 35392
rect 5744 35332 5748 35388
rect 5748 35332 5804 35388
rect 5804 35332 5808 35388
rect 5744 35328 5808 35332
rect 5824 35388 5888 35392
rect 5824 35332 5828 35388
rect 5828 35332 5884 35388
rect 5884 35332 5888 35388
rect 5824 35328 5888 35332
rect 14848 35388 14912 35392
rect 14848 35332 14852 35388
rect 14852 35332 14908 35388
rect 14908 35332 14912 35388
rect 14848 35328 14912 35332
rect 14928 35388 14992 35392
rect 14928 35332 14932 35388
rect 14932 35332 14988 35388
rect 14988 35332 14992 35388
rect 14928 35328 14992 35332
rect 15008 35388 15072 35392
rect 15008 35332 15012 35388
rect 15012 35332 15068 35388
rect 15068 35332 15072 35388
rect 15008 35328 15072 35332
rect 15088 35388 15152 35392
rect 15088 35332 15092 35388
rect 15092 35332 15148 35388
rect 15148 35332 15152 35388
rect 15088 35328 15152 35332
rect 24112 35388 24176 35392
rect 24112 35332 24116 35388
rect 24116 35332 24172 35388
rect 24172 35332 24176 35388
rect 24112 35328 24176 35332
rect 24192 35388 24256 35392
rect 24192 35332 24196 35388
rect 24196 35332 24252 35388
rect 24252 35332 24256 35388
rect 24192 35328 24256 35332
rect 24272 35388 24336 35392
rect 24272 35332 24276 35388
rect 24276 35332 24332 35388
rect 24332 35332 24336 35388
rect 24272 35328 24336 35332
rect 24352 35388 24416 35392
rect 24352 35332 24356 35388
rect 24356 35332 24412 35388
rect 24412 35332 24416 35388
rect 24352 35328 24416 35332
rect 18644 35124 18708 35188
rect 10216 34844 10280 34848
rect 10216 34788 10220 34844
rect 10220 34788 10276 34844
rect 10276 34788 10280 34844
rect 10216 34784 10280 34788
rect 10296 34844 10360 34848
rect 10296 34788 10300 34844
rect 10300 34788 10356 34844
rect 10356 34788 10360 34844
rect 10296 34784 10360 34788
rect 10376 34844 10440 34848
rect 10376 34788 10380 34844
rect 10380 34788 10436 34844
rect 10436 34788 10440 34844
rect 10376 34784 10440 34788
rect 10456 34844 10520 34848
rect 10456 34788 10460 34844
rect 10460 34788 10516 34844
rect 10516 34788 10520 34844
rect 10456 34784 10520 34788
rect 19480 34844 19544 34848
rect 19480 34788 19484 34844
rect 19484 34788 19540 34844
rect 19540 34788 19544 34844
rect 19480 34784 19544 34788
rect 19560 34844 19624 34848
rect 19560 34788 19564 34844
rect 19564 34788 19620 34844
rect 19620 34788 19624 34844
rect 19560 34784 19624 34788
rect 19640 34844 19704 34848
rect 19640 34788 19644 34844
rect 19644 34788 19700 34844
rect 19700 34788 19704 34844
rect 19640 34784 19704 34788
rect 19720 34844 19784 34848
rect 19720 34788 19724 34844
rect 19724 34788 19780 34844
rect 19780 34788 19784 34844
rect 19720 34784 19784 34788
rect 27476 34640 27540 34644
rect 27476 34584 27490 34640
rect 27490 34584 27540 34640
rect 27476 34580 27540 34584
rect 5584 34300 5648 34304
rect 5584 34244 5588 34300
rect 5588 34244 5644 34300
rect 5644 34244 5648 34300
rect 5584 34240 5648 34244
rect 5664 34300 5728 34304
rect 5664 34244 5668 34300
rect 5668 34244 5724 34300
rect 5724 34244 5728 34300
rect 5664 34240 5728 34244
rect 5744 34300 5808 34304
rect 5744 34244 5748 34300
rect 5748 34244 5804 34300
rect 5804 34244 5808 34300
rect 5744 34240 5808 34244
rect 5824 34300 5888 34304
rect 5824 34244 5828 34300
rect 5828 34244 5884 34300
rect 5884 34244 5888 34300
rect 5824 34240 5888 34244
rect 14848 34300 14912 34304
rect 14848 34244 14852 34300
rect 14852 34244 14908 34300
rect 14908 34244 14912 34300
rect 14848 34240 14912 34244
rect 14928 34300 14992 34304
rect 14928 34244 14932 34300
rect 14932 34244 14988 34300
rect 14988 34244 14992 34300
rect 14928 34240 14992 34244
rect 15008 34300 15072 34304
rect 15008 34244 15012 34300
rect 15012 34244 15068 34300
rect 15068 34244 15072 34300
rect 15008 34240 15072 34244
rect 15088 34300 15152 34304
rect 15088 34244 15092 34300
rect 15092 34244 15148 34300
rect 15148 34244 15152 34300
rect 15088 34240 15152 34244
rect 24112 34300 24176 34304
rect 24112 34244 24116 34300
rect 24116 34244 24172 34300
rect 24172 34244 24176 34300
rect 24112 34240 24176 34244
rect 24192 34300 24256 34304
rect 24192 34244 24196 34300
rect 24196 34244 24252 34300
rect 24252 34244 24256 34300
rect 24192 34240 24256 34244
rect 24272 34300 24336 34304
rect 24272 34244 24276 34300
rect 24276 34244 24332 34300
rect 24332 34244 24336 34300
rect 24272 34240 24336 34244
rect 24352 34300 24416 34304
rect 24352 34244 24356 34300
rect 24356 34244 24412 34300
rect 24412 34244 24416 34300
rect 24352 34240 24416 34244
rect 21772 33960 21836 33964
rect 21772 33904 21822 33960
rect 21822 33904 21836 33960
rect 21772 33900 21836 33904
rect 10216 33756 10280 33760
rect 10216 33700 10220 33756
rect 10220 33700 10276 33756
rect 10276 33700 10280 33756
rect 10216 33696 10280 33700
rect 10296 33756 10360 33760
rect 10296 33700 10300 33756
rect 10300 33700 10356 33756
rect 10356 33700 10360 33756
rect 10296 33696 10360 33700
rect 10376 33756 10440 33760
rect 10376 33700 10380 33756
rect 10380 33700 10436 33756
rect 10436 33700 10440 33756
rect 10376 33696 10440 33700
rect 10456 33756 10520 33760
rect 10456 33700 10460 33756
rect 10460 33700 10516 33756
rect 10516 33700 10520 33756
rect 10456 33696 10520 33700
rect 19480 33756 19544 33760
rect 19480 33700 19484 33756
rect 19484 33700 19540 33756
rect 19540 33700 19544 33756
rect 19480 33696 19544 33700
rect 19560 33756 19624 33760
rect 19560 33700 19564 33756
rect 19564 33700 19620 33756
rect 19620 33700 19624 33756
rect 19560 33696 19624 33700
rect 19640 33756 19704 33760
rect 19640 33700 19644 33756
rect 19644 33700 19700 33756
rect 19700 33700 19704 33756
rect 19640 33696 19704 33700
rect 19720 33756 19784 33760
rect 19720 33700 19724 33756
rect 19724 33700 19780 33756
rect 19780 33700 19784 33756
rect 19720 33696 19784 33700
rect 5584 33212 5648 33216
rect 5584 33156 5588 33212
rect 5588 33156 5644 33212
rect 5644 33156 5648 33212
rect 5584 33152 5648 33156
rect 5664 33212 5728 33216
rect 5664 33156 5668 33212
rect 5668 33156 5724 33212
rect 5724 33156 5728 33212
rect 5664 33152 5728 33156
rect 5744 33212 5808 33216
rect 5744 33156 5748 33212
rect 5748 33156 5804 33212
rect 5804 33156 5808 33212
rect 5744 33152 5808 33156
rect 5824 33212 5888 33216
rect 5824 33156 5828 33212
rect 5828 33156 5884 33212
rect 5884 33156 5888 33212
rect 5824 33152 5888 33156
rect 14848 33212 14912 33216
rect 14848 33156 14852 33212
rect 14852 33156 14908 33212
rect 14908 33156 14912 33212
rect 14848 33152 14912 33156
rect 14928 33212 14992 33216
rect 14928 33156 14932 33212
rect 14932 33156 14988 33212
rect 14988 33156 14992 33212
rect 14928 33152 14992 33156
rect 15008 33212 15072 33216
rect 15008 33156 15012 33212
rect 15012 33156 15068 33212
rect 15068 33156 15072 33212
rect 15008 33152 15072 33156
rect 15088 33212 15152 33216
rect 15088 33156 15092 33212
rect 15092 33156 15148 33212
rect 15148 33156 15152 33212
rect 15088 33152 15152 33156
rect 24112 33212 24176 33216
rect 24112 33156 24116 33212
rect 24116 33156 24172 33212
rect 24172 33156 24176 33212
rect 24112 33152 24176 33156
rect 24192 33212 24256 33216
rect 24192 33156 24196 33212
rect 24196 33156 24252 33212
rect 24252 33156 24256 33212
rect 24192 33152 24256 33156
rect 24272 33212 24336 33216
rect 24272 33156 24276 33212
rect 24276 33156 24332 33212
rect 24332 33156 24336 33212
rect 24272 33152 24336 33156
rect 24352 33212 24416 33216
rect 24352 33156 24356 33212
rect 24356 33156 24412 33212
rect 24412 33156 24416 33212
rect 24352 33152 24416 33156
rect 10216 32668 10280 32672
rect 10216 32612 10220 32668
rect 10220 32612 10276 32668
rect 10276 32612 10280 32668
rect 10216 32608 10280 32612
rect 10296 32668 10360 32672
rect 10296 32612 10300 32668
rect 10300 32612 10356 32668
rect 10356 32612 10360 32668
rect 10296 32608 10360 32612
rect 10376 32668 10440 32672
rect 10376 32612 10380 32668
rect 10380 32612 10436 32668
rect 10436 32612 10440 32668
rect 10376 32608 10440 32612
rect 10456 32668 10520 32672
rect 10456 32612 10460 32668
rect 10460 32612 10516 32668
rect 10516 32612 10520 32668
rect 10456 32608 10520 32612
rect 19480 32668 19544 32672
rect 19480 32612 19484 32668
rect 19484 32612 19540 32668
rect 19540 32612 19544 32668
rect 19480 32608 19544 32612
rect 19560 32668 19624 32672
rect 19560 32612 19564 32668
rect 19564 32612 19620 32668
rect 19620 32612 19624 32668
rect 19560 32608 19624 32612
rect 19640 32668 19704 32672
rect 19640 32612 19644 32668
rect 19644 32612 19700 32668
rect 19700 32612 19704 32668
rect 19640 32608 19704 32612
rect 19720 32668 19784 32672
rect 19720 32612 19724 32668
rect 19724 32612 19780 32668
rect 19780 32612 19784 32668
rect 19720 32608 19784 32612
rect 22508 32268 22572 32332
rect 5584 32124 5648 32128
rect 5584 32068 5588 32124
rect 5588 32068 5644 32124
rect 5644 32068 5648 32124
rect 5584 32064 5648 32068
rect 5664 32124 5728 32128
rect 5664 32068 5668 32124
rect 5668 32068 5724 32124
rect 5724 32068 5728 32124
rect 5664 32064 5728 32068
rect 5744 32124 5808 32128
rect 5744 32068 5748 32124
rect 5748 32068 5804 32124
rect 5804 32068 5808 32124
rect 5744 32064 5808 32068
rect 5824 32124 5888 32128
rect 5824 32068 5828 32124
rect 5828 32068 5884 32124
rect 5884 32068 5888 32124
rect 5824 32064 5888 32068
rect 14848 32124 14912 32128
rect 14848 32068 14852 32124
rect 14852 32068 14908 32124
rect 14908 32068 14912 32124
rect 14848 32064 14912 32068
rect 14928 32124 14992 32128
rect 14928 32068 14932 32124
rect 14932 32068 14988 32124
rect 14988 32068 14992 32124
rect 14928 32064 14992 32068
rect 15008 32124 15072 32128
rect 15008 32068 15012 32124
rect 15012 32068 15068 32124
rect 15068 32068 15072 32124
rect 15008 32064 15072 32068
rect 15088 32124 15152 32128
rect 15088 32068 15092 32124
rect 15092 32068 15148 32124
rect 15148 32068 15152 32124
rect 15088 32064 15152 32068
rect 24112 32124 24176 32128
rect 24112 32068 24116 32124
rect 24116 32068 24172 32124
rect 24172 32068 24176 32124
rect 24112 32064 24176 32068
rect 24192 32124 24256 32128
rect 24192 32068 24196 32124
rect 24196 32068 24252 32124
rect 24252 32068 24256 32124
rect 24192 32064 24256 32068
rect 24272 32124 24336 32128
rect 24272 32068 24276 32124
rect 24276 32068 24332 32124
rect 24332 32068 24336 32124
rect 24272 32064 24336 32068
rect 24352 32124 24416 32128
rect 24352 32068 24356 32124
rect 24356 32068 24412 32124
rect 24412 32068 24416 32124
rect 24352 32064 24416 32068
rect 10216 31580 10280 31584
rect 10216 31524 10220 31580
rect 10220 31524 10276 31580
rect 10276 31524 10280 31580
rect 10216 31520 10280 31524
rect 10296 31580 10360 31584
rect 10296 31524 10300 31580
rect 10300 31524 10356 31580
rect 10356 31524 10360 31580
rect 10296 31520 10360 31524
rect 10376 31580 10440 31584
rect 10376 31524 10380 31580
rect 10380 31524 10436 31580
rect 10436 31524 10440 31580
rect 10376 31520 10440 31524
rect 10456 31580 10520 31584
rect 10456 31524 10460 31580
rect 10460 31524 10516 31580
rect 10516 31524 10520 31580
rect 10456 31520 10520 31524
rect 19480 31580 19544 31584
rect 19480 31524 19484 31580
rect 19484 31524 19540 31580
rect 19540 31524 19544 31580
rect 19480 31520 19544 31524
rect 19560 31580 19624 31584
rect 19560 31524 19564 31580
rect 19564 31524 19620 31580
rect 19620 31524 19624 31580
rect 19560 31520 19624 31524
rect 19640 31580 19704 31584
rect 19640 31524 19644 31580
rect 19644 31524 19700 31580
rect 19700 31524 19704 31580
rect 19640 31520 19704 31524
rect 19720 31580 19784 31584
rect 19720 31524 19724 31580
rect 19724 31524 19780 31580
rect 19780 31524 19784 31580
rect 19720 31520 19784 31524
rect 5584 31036 5648 31040
rect 5584 30980 5588 31036
rect 5588 30980 5644 31036
rect 5644 30980 5648 31036
rect 5584 30976 5648 30980
rect 5664 31036 5728 31040
rect 5664 30980 5668 31036
rect 5668 30980 5724 31036
rect 5724 30980 5728 31036
rect 5664 30976 5728 30980
rect 5744 31036 5808 31040
rect 5744 30980 5748 31036
rect 5748 30980 5804 31036
rect 5804 30980 5808 31036
rect 5744 30976 5808 30980
rect 5824 31036 5888 31040
rect 5824 30980 5828 31036
rect 5828 30980 5884 31036
rect 5884 30980 5888 31036
rect 5824 30976 5888 30980
rect 14848 31036 14912 31040
rect 14848 30980 14852 31036
rect 14852 30980 14908 31036
rect 14908 30980 14912 31036
rect 14848 30976 14912 30980
rect 14928 31036 14992 31040
rect 14928 30980 14932 31036
rect 14932 30980 14988 31036
rect 14988 30980 14992 31036
rect 14928 30976 14992 30980
rect 15008 31036 15072 31040
rect 15008 30980 15012 31036
rect 15012 30980 15068 31036
rect 15068 30980 15072 31036
rect 15008 30976 15072 30980
rect 15088 31036 15152 31040
rect 15088 30980 15092 31036
rect 15092 30980 15148 31036
rect 15148 30980 15152 31036
rect 15088 30976 15152 30980
rect 24112 31036 24176 31040
rect 24112 30980 24116 31036
rect 24116 30980 24172 31036
rect 24172 30980 24176 31036
rect 24112 30976 24176 30980
rect 24192 31036 24256 31040
rect 24192 30980 24196 31036
rect 24196 30980 24252 31036
rect 24252 30980 24256 31036
rect 24192 30976 24256 30980
rect 24272 31036 24336 31040
rect 24272 30980 24276 31036
rect 24276 30980 24332 31036
rect 24332 30980 24336 31036
rect 24272 30976 24336 30980
rect 24352 31036 24416 31040
rect 24352 30980 24356 31036
rect 24356 30980 24412 31036
rect 24412 30980 24416 31036
rect 24352 30976 24416 30980
rect 10216 30492 10280 30496
rect 10216 30436 10220 30492
rect 10220 30436 10276 30492
rect 10276 30436 10280 30492
rect 10216 30432 10280 30436
rect 10296 30492 10360 30496
rect 10296 30436 10300 30492
rect 10300 30436 10356 30492
rect 10356 30436 10360 30492
rect 10296 30432 10360 30436
rect 10376 30492 10440 30496
rect 10376 30436 10380 30492
rect 10380 30436 10436 30492
rect 10436 30436 10440 30492
rect 10376 30432 10440 30436
rect 10456 30492 10520 30496
rect 10456 30436 10460 30492
rect 10460 30436 10516 30492
rect 10516 30436 10520 30492
rect 10456 30432 10520 30436
rect 19480 30492 19544 30496
rect 19480 30436 19484 30492
rect 19484 30436 19540 30492
rect 19540 30436 19544 30492
rect 19480 30432 19544 30436
rect 19560 30492 19624 30496
rect 19560 30436 19564 30492
rect 19564 30436 19620 30492
rect 19620 30436 19624 30492
rect 19560 30432 19624 30436
rect 19640 30492 19704 30496
rect 19640 30436 19644 30492
rect 19644 30436 19700 30492
rect 19700 30436 19704 30492
rect 19640 30432 19704 30436
rect 19720 30492 19784 30496
rect 19720 30436 19724 30492
rect 19724 30436 19780 30492
rect 19780 30436 19784 30492
rect 19720 30432 19784 30436
rect 5584 29948 5648 29952
rect 5584 29892 5588 29948
rect 5588 29892 5644 29948
rect 5644 29892 5648 29948
rect 5584 29888 5648 29892
rect 5664 29948 5728 29952
rect 5664 29892 5668 29948
rect 5668 29892 5724 29948
rect 5724 29892 5728 29948
rect 5664 29888 5728 29892
rect 5744 29948 5808 29952
rect 5744 29892 5748 29948
rect 5748 29892 5804 29948
rect 5804 29892 5808 29948
rect 5744 29888 5808 29892
rect 5824 29948 5888 29952
rect 5824 29892 5828 29948
rect 5828 29892 5884 29948
rect 5884 29892 5888 29948
rect 5824 29888 5888 29892
rect 14848 29948 14912 29952
rect 14848 29892 14852 29948
rect 14852 29892 14908 29948
rect 14908 29892 14912 29948
rect 14848 29888 14912 29892
rect 14928 29948 14992 29952
rect 14928 29892 14932 29948
rect 14932 29892 14988 29948
rect 14988 29892 14992 29948
rect 14928 29888 14992 29892
rect 15008 29948 15072 29952
rect 15008 29892 15012 29948
rect 15012 29892 15068 29948
rect 15068 29892 15072 29948
rect 15008 29888 15072 29892
rect 15088 29948 15152 29952
rect 15088 29892 15092 29948
rect 15092 29892 15148 29948
rect 15148 29892 15152 29948
rect 15088 29888 15152 29892
rect 24112 29948 24176 29952
rect 24112 29892 24116 29948
rect 24116 29892 24172 29948
rect 24172 29892 24176 29948
rect 24112 29888 24176 29892
rect 24192 29948 24256 29952
rect 24192 29892 24196 29948
rect 24196 29892 24252 29948
rect 24252 29892 24256 29948
rect 24192 29888 24256 29892
rect 24272 29948 24336 29952
rect 24272 29892 24276 29948
rect 24276 29892 24332 29948
rect 24332 29892 24336 29948
rect 24272 29888 24336 29892
rect 24352 29948 24416 29952
rect 24352 29892 24356 29948
rect 24356 29892 24412 29948
rect 24412 29892 24416 29948
rect 24352 29888 24416 29892
rect 10216 29404 10280 29408
rect 10216 29348 10220 29404
rect 10220 29348 10276 29404
rect 10276 29348 10280 29404
rect 10216 29344 10280 29348
rect 10296 29404 10360 29408
rect 10296 29348 10300 29404
rect 10300 29348 10356 29404
rect 10356 29348 10360 29404
rect 10296 29344 10360 29348
rect 10376 29404 10440 29408
rect 10376 29348 10380 29404
rect 10380 29348 10436 29404
rect 10436 29348 10440 29404
rect 10376 29344 10440 29348
rect 10456 29404 10520 29408
rect 10456 29348 10460 29404
rect 10460 29348 10516 29404
rect 10516 29348 10520 29404
rect 10456 29344 10520 29348
rect 19480 29404 19544 29408
rect 19480 29348 19484 29404
rect 19484 29348 19540 29404
rect 19540 29348 19544 29404
rect 19480 29344 19544 29348
rect 19560 29404 19624 29408
rect 19560 29348 19564 29404
rect 19564 29348 19620 29404
rect 19620 29348 19624 29404
rect 19560 29344 19624 29348
rect 19640 29404 19704 29408
rect 19640 29348 19644 29404
rect 19644 29348 19700 29404
rect 19700 29348 19704 29404
rect 19640 29344 19704 29348
rect 19720 29404 19784 29408
rect 19720 29348 19724 29404
rect 19724 29348 19780 29404
rect 19780 29348 19784 29404
rect 19720 29344 19784 29348
rect 5584 28860 5648 28864
rect 5584 28804 5588 28860
rect 5588 28804 5644 28860
rect 5644 28804 5648 28860
rect 5584 28800 5648 28804
rect 5664 28860 5728 28864
rect 5664 28804 5668 28860
rect 5668 28804 5724 28860
rect 5724 28804 5728 28860
rect 5664 28800 5728 28804
rect 5744 28860 5808 28864
rect 5744 28804 5748 28860
rect 5748 28804 5804 28860
rect 5804 28804 5808 28860
rect 5744 28800 5808 28804
rect 5824 28860 5888 28864
rect 5824 28804 5828 28860
rect 5828 28804 5884 28860
rect 5884 28804 5888 28860
rect 5824 28800 5888 28804
rect 14848 28860 14912 28864
rect 14848 28804 14852 28860
rect 14852 28804 14908 28860
rect 14908 28804 14912 28860
rect 14848 28800 14912 28804
rect 14928 28860 14992 28864
rect 14928 28804 14932 28860
rect 14932 28804 14988 28860
rect 14988 28804 14992 28860
rect 14928 28800 14992 28804
rect 15008 28860 15072 28864
rect 15008 28804 15012 28860
rect 15012 28804 15068 28860
rect 15068 28804 15072 28860
rect 15008 28800 15072 28804
rect 15088 28860 15152 28864
rect 15088 28804 15092 28860
rect 15092 28804 15148 28860
rect 15148 28804 15152 28860
rect 15088 28800 15152 28804
rect 24112 28860 24176 28864
rect 24112 28804 24116 28860
rect 24116 28804 24172 28860
rect 24172 28804 24176 28860
rect 24112 28800 24176 28804
rect 24192 28860 24256 28864
rect 24192 28804 24196 28860
rect 24196 28804 24252 28860
rect 24252 28804 24256 28860
rect 24192 28800 24256 28804
rect 24272 28860 24336 28864
rect 24272 28804 24276 28860
rect 24276 28804 24332 28860
rect 24332 28804 24336 28860
rect 24272 28800 24336 28804
rect 24352 28860 24416 28864
rect 24352 28804 24356 28860
rect 24356 28804 24412 28860
rect 24412 28804 24416 28860
rect 24352 28800 24416 28804
rect 10216 28316 10280 28320
rect 10216 28260 10220 28316
rect 10220 28260 10276 28316
rect 10276 28260 10280 28316
rect 10216 28256 10280 28260
rect 10296 28316 10360 28320
rect 10296 28260 10300 28316
rect 10300 28260 10356 28316
rect 10356 28260 10360 28316
rect 10296 28256 10360 28260
rect 10376 28316 10440 28320
rect 10376 28260 10380 28316
rect 10380 28260 10436 28316
rect 10436 28260 10440 28316
rect 10376 28256 10440 28260
rect 10456 28316 10520 28320
rect 10456 28260 10460 28316
rect 10460 28260 10516 28316
rect 10516 28260 10520 28316
rect 10456 28256 10520 28260
rect 19480 28316 19544 28320
rect 19480 28260 19484 28316
rect 19484 28260 19540 28316
rect 19540 28260 19544 28316
rect 19480 28256 19544 28260
rect 19560 28316 19624 28320
rect 19560 28260 19564 28316
rect 19564 28260 19620 28316
rect 19620 28260 19624 28316
rect 19560 28256 19624 28260
rect 19640 28316 19704 28320
rect 19640 28260 19644 28316
rect 19644 28260 19700 28316
rect 19700 28260 19704 28316
rect 19640 28256 19704 28260
rect 19720 28316 19784 28320
rect 19720 28260 19724 28316
rect 19724 28260 19780 28316
rect 19780 28260 19784 28316
rect 19720 28256 19784 28260
rect 5584 27772 5648 27776
rect 5584 27716 5588 27772
rect 5588 27716 5644 27772
rect 5644 27716 5648 27772
rect 5584 27712 5648 27716
rect 5664 27772 5728 27776
rect 5664 27716 5668 27772
rect 5668 27716 5724 27772
rect 5724 27716 5728 27772
rect 5664 27712 5728 27716
rect 5744 27772 5808 27776
rect 5744 27716 5748 27772
rect 5748 27716 5804 27772
rect 5804 27716 5808 27772
rect 5744 27712 5808 27716
rect 5824 27772 5888 27776
rect 5824 27716 5828 27772
rect 5828 27716 5884 27772
rect 5884 27716 5888 27772
rect 5824 27712 5888 27716
rect 14848 27772 14912 27776
rect 14848 27716 14852 27772
rect 14852 27716 14908 27772
rect 14908 27716 14912 27772
rect 14848 27712 14912 27716
rect 14928 27772 14992 27776
rect 14928 27716 14932 27772
rect 14932 27716 14988 27772
rect 14988 27716 14992 27772
rect 14928 27712 14992 27716
rect 15008 27772 15072 27776
rect 15008 27716 15012 27772
rect 15012 27716 15068 27772
rect 15068 27716 15072 27772
rect 15008 27712 15072 27716
rect 15088 27772 15152 27776
rect 15088 27716 15092 27772
rect 15092 27716 15148 27772
rect 15148 27716 15152 27772
rect 15088 27712 15152 27716
rect 24112 27772 24176 27776
rect 24112 27716 24116 27772
rect 24116 27716 24172 27772
rect 24172 27716 24176 27772
rect 24112 27712 24176 27716
rect 24192 27772 24256 27776
rect 24192 27716 24196 27772
rect 24196 27716 24252 27772
rect 24252 27716 24256 27772
rect 24192 27712 24256 27716
rect 24272 27772 24336 27776
rect 24272 27716 24276 27772
rect 24276 27716 24332 27772
rect 24332 27716 24336 27772
rect 24272 27712 24336 27716
rect 24352 27772 24416 27776
rect 24352 27716 24356 27772
rect 24356 27716 24412 27772
rect 24412 27716 24416 27772
rect 24352 27712 24416 27716
rect 10216 27228 10280 27232
rect 10216 27172 10220 27228
rect 10220 27172 10276 27228
rect 10276 27172 10280 27228
rect 10216 27168 10280 27172
rect 10296 27228 10360 27232
rect 10296 27172 10300 27228
rect 10300 27172 10356 27228
rect 10356 27172 10360 27228
rect 10296 27168 10360 27172
rect 10376 27228 10440 27232
rect 10376 27172 10380 27228
rect 10380 27172 10436 27228
rect 10436 27172 10440 27228
rect 10376 27168 10440 27172
rect 10456 27228 10520 27232
rect 10456 27172 10460 27228
rect 10460 27172 10516 27228
rect 10516 27172 10520 27228
rect 10456 27168 10520 27172
rect 19480 27228 19544 27232
rect 19480 27172 19484 27228
rect 19484 27172 19540 27228
rect 19540 27172 19544 27228
rect 19480 27168 19544 27172
rect 19560 27228 19624 27232
rect 19560 27172 19564 27228
rect 19564 27172 19620 27228
rect 19620 27172 19624 27228
rect 19560 27168 19624 27172
rect 19640 27228 19704 27232
rect 19640 27172 19644 27228
rect 19644 27172 19700 27228
rect 19700 27172 19704 27228
rect 19640 27168 19704 27172
rect 19720 27228 19784 27232
rect 19720 27172 19724 27228
rect 19724 27172 19780 27228
rect 19780 27172 19784 27228
rect 19720 27168 19784 27172
rect 5584 26684 5648 26688
rect 5584 26628 5588 26684
rect 5588 26628 5644 26684
rect 5644 26628 5648 26684
rect 5584 26624 5648 26628
rect 5664 26684 5728 26688
rect 5664 26628 5668 26684
rect 5668 26628 5724 26684
rect 5724 26628 5728 26684
rect 5664 26624 5728 26628
rect 5744 26684 5808 26688
rect 5744 26628 5748 26684
rect 5748 26628 5804 26684
rect 5804 26628 5808 26684
rect 5744 26624 5808 26628
rect 5824 26684 5888 26688
rect 5824 26628 5828 26684
rect 5828 26628 5884 26684
rect 5884 26628 5888 26684
rect 5824 26624 5888 26628
rect 14848 26684 14912 26688
rect 14848 26628 14852 26684
rect 14852 26628 14908 26684
rect 14908 26628 14912 26684
rect 14848 26624 14912 26628
rect 14928 26684 14992 26688
rect 14928 26628 14932 26684
rect 14932 26628 14988 26684
rect 14988 26628 14992 26684
rect 14928 26624 14992 26628
rect 15008 26684 15072 26688
rect 15008 26628 15012 26684
rect 15012 26628 15068 26684
rect 15068 26628 15072 26684
rect 15008 26624 15072 26628
rect 15088 26684 15152 26688
rect 15088 26628 15092 26684
rect 15092 26628 15148 26684
rect 15148 26628 15152 26684
rect 15088 26624 15152 26628
rect 24112 26684 24176 26688
rect 24112 26628 24116 26684
rect 24116 26628 24172 26684
rect 24172 26628 24176 26684
rect 24112 26624 24176 26628
rect 24192 26684 24256 26688
rect 24192 26628 24196 26684
rect 24196 26628 24252 26684
rect 24252 26628 24256 26684
rect 24192 26624 24256 26628
rect 24272 26684 24336 26688
rect 24272 26628 24276 26684
rect 24276 26628 24332 26684
rect 24332 26628 24336 26684
rect 24272 26624 24336 26628
rect 24352 26684 24416 26688
rect 24352 26628 24356 26684
rect 24356 26628 24412 26684
rect 24412 26628 24416 26684
rect 24352 26624 24416 26628
rect 10216 26140 10280 26144
rect 10216 26084 10220 26140
rect 10220 26084 10276 26140
rect 10276 26084 10280 26140
rect 10216 26080 10280 26084
rect 10296 26140 10360 26144
rect 10296 26084 10300 26140
rect 10300 26084 10356 26140
rect 10356 26084 10360 26140
rect 10296 26080 10360 26084
rect 10376 26140 10440 26144
rect 10376 26084 10380 26140
rect 10380 26084 10436 26140
rect 10436 26084 10440 26140
rect 10376 26080 10440 26084
rect 10456 26140 10520 26144
rect 10456 26084 10460 26140
rect 10460 26084 10516 26140
rect 10516 26084 10520 26140
rect 10456 26080 10520 26084
rect 19480 26140 19544 26144
rect 19480 26084 19484 26140
rect 19484 26084 19540 26140
rect 19540 26084 19544 26140
rect 19480 26080 19544 26084
rect 19560 26140 19624 26144
rect 19560 26084 19564 26140
rect 19564 26084 19620 26140
rect 19620 26084 19624 26140
rect 19560 26080 19624 26084
rect 19640 26140 19704 26144
rect 19640 26084 19644 26140
rect 19644 26084 19700 26140
rect 19700 26084 19704 26140
rect 19640 26080 19704 26084
rect 19720 26140 19784 26144
rect 19720 26084 19724 26140
rect 19724 26084 19780 26140
rect 19780 26084 19784 26140
rect 19720 26080 19784 26084
rect 5584 25596 5648 25600
rect 5584 25540 5588 25596
rect 5588 25540 5644 25596
rect 5644 25540 5648 25596
rect 5584 25536 5648 25540
rect 5664 25596 5728 25600
rect 5664 25540 5668 25596
rect 5668 25540 5724 25596
rect 5724 25540 5728 25596
rect 5664 25536 5728 25540
rect 5744 25596 5808 25600
rect 5744 25540 5748 25596
rect 5748 25540 5804 25596
rect 5804 25540 5808 25596
rect 5744 25536 5808 25540
rect 5824 25596 5888 25600
rect 5824 25540 5828 25596
rect 5828 25540 5884 25596
rect 5884 25540 5888 25596
rect 5824 25536 5888 25540
rect 14848 25596 14912 25600
rect 14848 25540 14852 25596
rect 14852 25540 14908 25596
rect 14908 25540 14912 25596
rect 14848 25536 14912 25540
rect 14928 25596 14992 25600
rect 14928 25540 14932 25596
rect 14932 25540 14988 25596
rect 14988 25540 14992 25596
rect 14928 25536 14992 25540
rect 15008 25596 15072 25600
rect 15008 25540 15012 25596
rect 15012 25540 15068 25596
rect 15068 25540 15072 25596
rect 15008 25536 15072 25540
rect 15088 25596 15152 25600
rect 15088 25540 15092 25596
rect 15092 25540 15148 25596
rect 15148 25540 15152 25596
rect 15088 25536 15152 25540
rect 24112 25596 24176 25600
rect 24112 25540 24116 25596
rect 24116 25540 24172 25596
rect 24172 25540 24176 25596
rect 24112 25536 24176 25540
rect 24192 25596 24256 25600
rect 24192 25540 24196 25596
rect 24196 25540 24252 25596
rect 24252 25540 24256 25596
rect 24192 25536 24256 25540
rect 24272 25596 24336 25600
rect 24272 25540 24276 25596
rect 24276 25540 24332 25596
rect 24332 25540 24336 25596
rect 24272 25536 24336 25540
rect 24352 25596 24416 25600
rect 24352 25540 24356 25596
rect 24356 25540 24412 25596
rect 24412 25540 24416 25596
rect 24352 25536 24416 25540
rect 10216 25052 10280 25056
rect 10216 24996 10220 25052
rect 10220 24996 10276 25052
rect 10276 24996 10280 25052
rect 10216 24992 10280 24996
rect 10296 25052 10360 25056
rect 10296 24996 10300 25052
rect 10300 24996 10356 25052
rect 10356 24996 10360 25052
rect 10296 24992 10360 24996
rect 10376 25052 10440 25056
rect 10376 24996 10380 25052
rect 10380 24996 10436 25052
rect 10436 24996 10440 25052
rect 10376 24992 10440 24996
rect 10456 25052 10520 25056
rect 10456 24996 10460 25052
rect 10460 24996 10516 25052
rect 10516 24996 10520 25052
rect 10456 24992 10520 24996
rect 19480 25052 19544 25056
rect 19480 24996 19484 25052
rect 19484 24996 19540 25052
rect 19540 24996 19544 25052
rect 19480 24992 19544 24996
rect 19560 25052 19624 25056
rect 19560 24996 19564 25052
rect 19564 24996 19620 25052
rect 19620 24996 19624 25052
rect 19560 24992 19624 24996
rect 19640 25052 19704 25056
rect 19640 24996 19644 25052
rect 19644 24996 19700 25052
rect 19700 24996 19704 25052
rect 19640 24992 19704 24996
rect 19720 25052 19784 25056
rect 19720 24996 19724 25052
rect 19724 24996 19780 25052
rect 19780 24996 19784 25052
rect 19720 24992 19784 24996
rect 5584 24508 5648 24512
rect 5584 24452 5588 24508
rect 5588 24452 5644 24508
rect 5644 24452 5648 24508
rect 5584 24448 5648 24452
rect 5664 24508 5728 24512
rect 5664 24452 5668 24508
rect 5668 24452 5724 24508
rect 5724 24452 5728 24508
rect 5664 24448 5728 24452
rect 5744 24508 5808 24512
rect 5744 24452 5748 24508
rect 5748 24452 5804 24508
rect 5804 24452 5808 24508
rect 5744 24448 5808 24452
rect 5824 24508 5888 24512
rect 5824 24452 5828 24508
rect 5828 24452 5884 24508
rect 5884 24452 5888 24508
rect 5824 24448 5888 24452
rect 14848 24508 14912 24512
rect 14848 24452 14852 24508
rect 14852 24452 14908 24508
rect 14908 24452 14912 24508
rect 14848 24448 14912 24452
rect 14928 24508 14992 24512
rect 14928 24452 14932 24508
rect 14932 24452 14988 24508
rect 14988 24452 14992 24508
rect 14928 24448 14992 24452
rect 15008 24508 15072 24512
rect 15008 24452 15012 24508
rect 15012 24452 15068 24508
rect 15068 24452 15072 24508
rect 15008 24448 15072 24452
rect 15088 24508 15152 24512
rect 15088 24452 15092 24508
rect 15092 24452 15148 24508
rect 15148 24452 15152 24508
rect 15088 24448 15152 24452
rect 24112 24508 24176 24512
rect 24112 24452 24116 24508
rect 24116 24452 24172 24508
rect 24172 24452 24176 24508
rect 24112 24448 24176 24452
rect 24192 24508 24256 24512
rect 24192 24452 24196 24508
rect 24196 24452 24252 24508
rect 24252 24452 24256 24508
rect 24192 24448 24256 24452
rect 24272 24508 24336 24512
rect 24272 24452 24276 24508
rect 24276 24452 24332 24508
rect 24332 24452 24336 24508
rect 24272 24448 24336 24452
rect 24352 24508 24416 24512
rect 24352 24452 24356 24508
rect 24356 24452 24412 24508
rect 24412 24452 24416 24508
rect 24352 24448 24416 24452
rect 21956 24108 22020 24172
rect 10216 23964 10280 23968
rect 10216 23908 10220 23964
rect 10220 23908 10276 23964
rect 10276 23908 10280 23964
rect 10216 23904 10280 23908
rect 10296 23964 10360 23968
rect 10296 23908 10300 23964
rect 10300 23908 10356 23964
rect 10356 23908 10360 23964
rect 10296 23904 10360 23908
rect 10376 23964 10440 23968
rect 10376 23908 10380 23964
rect 10380 23908 10436 23964
rect 10436 23908 10440 23964
rect 10376 23904 10440 23908
rect 10456 23964 10520 23968
rect 10456 23908 10460 23964
rect 10460 23908 10516 23964
rect 10516 23908 10520 23964
rect 10456 23904 10520 23908
rect 19480 23964 19544 23968
rect 19480 23908 19484 23964
rect 19484 23908 19540 23964
rect 19540 23908 19544 23964
rect 19480 23904 19544 23908
rect 19560 23964 19624 23968
rect 19560 23908 19564 23964
rect 19564 23908 19620 23964
rect 19620 23908 19624 23964
rect 19560 23904 19624 23908
rect 19640 23964 19704 23968
rect 19640 23908 19644 23964
rect 19644 23908 19700 23964
rect 19700 23908 19704 23964
rect 19640 23904 19704 23908
rect 19720 23964 19784 23968
rect 19720 23908 19724 23964
rect 19724 23908 19780 23964
rect 19780 23908 19784 23964
rect 19720 23904 19784 23908
rect 21772 23428 21836 23492
rect 5584 23420 5648 23424
rect 5584 23364 5588 23420
rect 5588 23364 5644 23420
rect 5644 23364 5648 23420
rect 5584 23360 5648 23364
rect 5664 23420 5728 23424
rect 5664 23364 5668 23420
rect 5668 23364 5724 23420
rect 5724 23364 5728 23420
rect 5664 23360 5728 23364
rect 5744 23420 5808 23424
rect 5744 23364 5748 23420
rect 5748 23364 5804 23420
rect 5804 23364 5808 23420
rect 5744 23360 5808 23364
rect 5824 23420 5888 23424
rect 5824 23364 5828 23420
rect 5828 23364 5884 23420
rect 5884 23364 5888 23420
rect 5824 23360 5888 23364
rect 14848 23420 14912 23424
rect 14848 23364 14852 23420
rect 14852 23364 14908 23420
rect 14908 23364 14912 23420
rect 14848 23360 14912 23364
rect 14928 23420 14992 23424
rect 14928 23364 14932 23420
rect 14932 23364 14988 23420
rect 14988 23364 14992 23420
rect 14928 23360 14992 23364
rect 15008 23420 15072 23424
rect 15008 23364 15012 23420
rect 15012 23364 15068 23420
rect 15068 23364 15072 23420
rect 15008 23360 15072 23364
rect 15088 23420 15152 23424
rect 15088 23364 15092 23420
rect 15092 23364 15148 23420
rect 15148 23364 15152 23420
rect 15088 23360 15152 23364
rect 24112 23420 24176 23424
rect 24112 23364 24116 23420
rect 24116 23364 24172 23420
rect 24172 23364 24176 23420
rect 24112 23360 24176 23364
rect 24192 23420 24256 23424
rect 24192 23364 24196 23420
rect 24196 23364 24252 23420
rect 24252 23364 24256 23420
rect 24192 23360 24256 23364
rect 24272 23420 24336 23424
rect 24272 23364 24276 23420
rect 24276 23364 24332 23420
rect 24332 23364 24336 23420
rect 24272 23360 24336 23364
rect 24352 23420 24416 23424
rect 24352 23364 24356 23420
rect 24356 23364 24412 23420
rect 24412 23364 24416 23420
rect 24352 23360 24416 23364
rect 10216 22876 10280 22880
rect 10216 22820 10220 22876
rect 10220 22820 10276 22876
rect 10276 22820 10280 22876
rect 10216 22816 10280 22820
rect 10296 22876 10360 22880
rect 10296 22820 10300 22876
rect 10300 22820 10356 22876
rect 10356 22820 10360 22876
rect 10296 22816 10360 22820
rect 10376 22876 10440 22880
rect 10376 22820 10380 22876
rect 10380 22820 10436 22876
rect 10436 22820 10440 22876
rect 10376 22816 10440 22820
rect 10456 22876 10520 22880
rect 10456 22820 10460 22876
rect 10460 22820 10516 22876
rect 10516 22820 10520 22876
rect 10456 22816 10520 22820
rect 19480 22876 19544 22880
rect 19480 22820 19484 22876
rect 19484 22820 19540 22876
rect 19540 22820 19544 22876
rect 19480 22816 19544 22820
rect 19560 22876 19624 22880
rect 19560 22820 19564 22876
rect 19564 22820 19620 22876
rect 19620 22820 19624 22876
rect 19560 22816 19624 22820
rect 19640 22876 19704 22880
rect 19640 22820 19644 22876
rect 19644 22820 19700 22876
rect 19700 22820 19704 22876
rect 19640 22816 19704 22820
rect 19720 22876 19784 22880
rect 19720 22820 19724 22876
rect 19724 22820 19780 22876
rect 19780 22820 19784 22876
rect 19720 22816 19784 22820
rect 5584 22332 5648 22336
rect 5584 22276 5588 22332
rect 5588 22276 5644 22332
rect 5644 22276 5648 22332
rect 5584 22272 5648 22276
rect 5664 22332 5728 22336
rect 5664 22276 5668 22332
rect 5668 22276 5724 22332
rect 5724 22276 5728 22332
rect 5664 22272 5728 22276
rect 5744 22332 5808 22336
rect 5744 22276 5748 22332
rect 5748 22276 5804 22332
rect 5804 22276 5808 22332
rect 5744 22272 5808 22276
rect 5824 22332 5888 22336
rect 5824 22276 5828 22332
rect 5828 22276 5884 22332
rect 5884 22276 5888 22332
rect 5824 22272 5888 22276
rect 14848 22332 14912 22336
rect 14848 22276 14852 22332
rect 14852 22276 14908 22332
rect 14908 22276 14912 22332
rect 14848 22272 14912 22276
rect 14928 22332 14992 22336
rect 14928 22276 14932 22332
rect 14932 22276 14988 22332
rect 14988 22276 14992 22332
rect 14928 22272 14992 22276
rect 15008 22332 15072 22336
rect 15008 22276 15012 22332
rect 15012 22276 15068 22332
rect 15068 22276 15072 22332
rect 15008 22272 15072 22276
rect 15088 22332 15152 22336
rect 15088 22276 15092 22332
rect 15092 22276 15148 22332
rect 15148 22276 15152 22332
rect 15088 22272 15152 22276
rect 24112 22332 24176 22336
rect 24112 22276 24116 22332
rect 24116 22276 24172 22332
rect 24172 22276 24176 22332
rect 24112 22272 24176 22276
rect 24192 22332 24256 22336
rect 24192 22276 24196 22332
rect 24196 22276 24252 22332
rect 24252 22276 24256 22332
rect 24192 22272 24256 22276
rect 24272 22332 24336 22336
rect 24272 22276 24276 22332
rect 24276 22276 24332 22332
rect 24332 22276 24336 22332
rect 24272 22272 24336 22276
rect 24352 22332 24416 22336
rect 24352 22276 24356 22332
rect 24356 22276 24412 22332
rect 24412 22276 24416 22332
rect 24352 22272 24416 22276
rect 10216 21788 10280 21792
rect 10216 21732 10220 21788
rect 10220 21732 10276 21788
rect 10276 21732 10280 21788
rect 10216 21728 10280 21732
rect 10296 21788 10360 21792
rect 10296 21732 10300 21788
rect 10300 21732 10356 21788
rect 10356 21732 10360 21788
rect 10296 21728 10360 21732
rect 10376 21788 10440 21792
rect 10376 21732 10380 21788
rect 10380 21732 10436 21788
rect 10436 21732 10440 21788
rect 10376 21728 10440 21732
rect 10456 21788 10520 21792
rect 10456 21732 10460 21788
rect 10460 21732 10516 21788
rect 10516 21732 10520 21788
rect 10456 21728 10520 21732
rect 19480 21788 19544 21792
rect 19480 21732 19484 21788
rect 19484 21732 19540 21788
rect 19540 21732 19544 21788
rect 19480 21728 19544 21732
rect 19560 21788 19624 21792
rect 19560 21732 19564 21788
rect 19564 21732 19620 21788
rect 19620 21732 19624 21788
rect 19560 21728 19624 21732
rect 19640 21788 19704 21792
rect 19640 21732 19644 21788
rect 19644 21732 19700 21788
rect 19700 21732 19704 21788
rect 19640 21728 19704 21732
rect 19720 21788 19784 21792
rect 19720 21732 19724 21788
rect 19724 21732 19780 21788
rect 19780 21732 19784 21788
rect 19720 21728 19784 21732
rect 22508 21524 22572 21588
rect 5584 21244 5648 21248
rect 5584 21188 5588 21244
rect 5588 21188 5644 21244
rect 5644 21188 5648 21244
rect 5584 21184 5648 21188
rect 5664 21244 5728 21248
rect 5664 21188 5668 21244
rect 5668 21188 5724 21244
rect 5724 21188 5728 21244
rect 5664 21184 5728 21188
rect 5744 21244 5808 21248
rect 5744 21188 5748 21244
rect 5748 21188 5804 21244
rect 5804 21188 5808 21244
rect 5744 21184 5808 21188
rect 5824 21244 5888 21248
rect 5824 21188 5828 21244
rect 5828 21188 5884 21244
rect 5884 21188 5888 21244
rect 5824 21184 5888 21188
rect 14848 21244 14912 21248
rect 14848 21188 14852 21244
rect 14852 21188 14908 21244
rect 14908 21188 14912 21244
rect 14848 21184 14912 21188
rect 14928 21244 14992 21248
rect 14928 21188 14932 21244
rect 14932 21188 14988 21244
rect 14988 21188 14992 21244
rect 14928 21184 14992 21188
rect 15008 21244 15072 21248
rect 15008 21188 15012 21244
rect 15012 21188 15068 21244
rect 15068 21188 15072 21244
rect 15008 21184 15072 21188
rect 15088 21244 15152 21248
rect 15088 21188 15092 21244
rect 15092 21188 15148 21244
rect 15148 21188 15152 21244
rect 15088 21184 15152 21188
rect 24112 21244 24176 21248
rect 24112 21188 24116 21244
rect 24116 21188 24172 21244
rect 24172 21188 24176 21244
rect 24112 21184 24176 21188
rect 24192 21244 24256 21248
rect 24192 21188 24196 21244
rect 24196 21188 24252 21244
rect 24252 21188 24256 21244
rect 24192 21184 24256 21188
rect 24272 21244 24336 21248
rect 24272 21188 24276 21244
rect 24276 21188 24332 21244
rect 24332 21188 24336 21244
rect 24272 21184 24336 21188
rect 24352 21244 24416 21248
rect 24352 21188 24356 21244
rect 24356 21188 24412 21244
rect 24412 21188 24416 21244
rect 24352 21184 24416 21188
rect 10216 20700 10280 20704
rect 10216 20644 10220 20700
rect 10220 20644 10276 20700
rect 10276 20644 10280 20700
rect 10216 20640 10280 20644
rect 10296 20700 10360 20704
rect 10296 20644 10300 20700
rect 10300 20644 10356 20700
rect 10356 20644 10360 20700
rect 10296 20640 10360 20644
rect 10376 20700 10440 20704
rect 10376 20644 10380 20700
rect 10380 20644 10436 20700
rect 10436 20644 10440 20700
rect 10376 20640 10440 20644
rect 10456 20700 10520 20704
rect 10456 20644 10460 20700
rect 10460 20644 10516 20700
rect 10516 20644 10520 20700
rect 10456 20640 10520 20644
rect 19480 20700 19544 20704
rect 19480 20644 19484 20700
rect 19484 20644 19540 20700
rect 19540 20644 19544 20700
rect 19480 20640 19544 20644
rect 19560 20700 19624 20704
rect 19560 20644 19564 20700
rect 19564 20644 19620 20700
rect 19620 20644 19624 20700
rect 19560 20640 19624 20644
rect 19640 20700 19704 20704
rect 19640 20644 19644 20700
rect 19644 20644 19700 20700
rect 19700 20644 19704 20700
rect 19640 20640 19704 20644
rect 19720 20700 19784 20704
rect 19720 20644 19724 20700
rect 19724 20644 19780 20700
rect 19780 20644 19784 20700
rect 19720 20640 19784 20644
rect 27292 20360 27356 20364
rect 27292 20304 27342 20360
rect 27342 20304 27356 20360
rect 27292 20300 27356 20304
rect 5584 20156 5648 20160
rect 5584 20100 5588 20156
rect 5588 20100 5644 20156
rect 5644 20100 5648 20156
rect 5584 20096 5648 20100
rect 5664 20156 5728 20160
rect 5664 20100 5668 20156
rect 5668 20100 5724 20156
rect 5724 20100 5728 20156
rect 5664 20096 5728 20100
rect 5744 20156 5808 20160
rect 5744 20100 5748 20156
rect 5748 20100 5804 20156
rect 5804 20100 5808 20156
rect 5744 20096 5808 20100
rect 5824 20156 5888 20160
rect 5824 20100 5828 20156
rect 5828 20100 5884 20156
rect 5884 20100 5888 20156
rect 5824 20096 5888 20100
rect 14848 20156 14912 20160
rect 14848 20100 14852 20156
rect 14852 20100 14908 20156
rect 14908 20100 14912 20156
rect 14848 20096 14912 20100
rect 14928 20156 14992 20160
rect 14928 20100 14932 20156
rect 14932 20100 14988 20156
rect 14988 20100 14992 20156
rect 14928 20096 14992 20100
rect 15008 20156 15072 20160
rect 15008 20100 15012 20156
rect 15012 20100 15068 20156
rect 15068 20100 15072 20156
rect 15008 20096 15072 20100
rect 15088 20156 15152 20160
rect 15088 20100 15092 20156
rect 15092 20100 15148 20156
rect 15148 20100 15152 20156
rect 15088 20096 15152 20100
rect 24112 20156 24176 20160
rect 24112 20100 24116 20156
rect 24116 20100 24172 20156
rect 24172 20100 24176 20156
rect 24112 20096 24176 20100
rect 24192 20156 24256 20160
rect 24192 20100 24196 20156
rect 24196 20100 24252 20156
rect 24252 20100 24256 20156
rect 24192 20096 24256 20100
rect 24272 20156 24336 20160
rect 24272 20100 24276 20156
rect 24276 20100 24332 20156
rect 24332 20100 24336 20156
rect 24272 20096 24336 20100
rect 24352 20156 24416 20160
rect 24352 20100 24356 20156
rect 24356 20100 24412 20156
rect 24412 20100 24416 20156
rect 24352 20096 24416 20100
rect 10216 19612 10280 19616
rect 10216 19556 10220 19612
rect 10220 19556 10276 19612
rect 10276 19556 10280 19612
rect 10216 19552 10280 19556
rect 10296 19612 10360 19616
rect 10296 19556 10300 19612
rect 10300 19556 10356 19612
rect 10356 19556 10360 19612
rect 10296 19552 10360 19556
rect 10376 19612 10440 19616
rect 10376 19556 10380 19612
rect 10380 19556 10436 19612
rect 10436 19556 10440 19612
rect 10376 19552 10440 19556
rect 10456 19612 10520 19616
rect 10456 19556 10460 19612
rect 10460 19556 10516 19612
rect 10516 19556 10520 19612
rect 10456 19552 10520 19556
rect 19480 19612 19544 19616
rect 19480 19556 19484 19612
rect 19484 19556 19540 19612
rect 19540 19556 19544 19612
rect 19480 19552 19544 19556
rect 19560 19612 19624 19616
rect 19560 19556 19564 19612
rect 19564 19556 19620 19612
rect 19620 19556 19624 19612
rect 19560 19552 19624 19556
rect 19640 19612 19704 19616
rect 19640 19556 19644 19612
rect 19644 19556 19700 19612
rect 19700 19556 19704 19612
rect 19640 19552 19704 19556
rect 19720 19612 19784 19616
rect 19720 19556 19724 19612
rect 19724 19556 19780 19612
rect 19780 19556 19784 19612
rect 19720 19552 19784 19556
rect 5584 19068 5648 19072
rect 5584 19012 5588 19068
rect 5588 19012 5644 19068
rect 5644 19012 5648 19068
rect 5584 19008 5648 19012
rect 5664 19068 5728 19072
rect 5664 19012 5668 19068
rect 5668 19012 5724 19068
rect 5724 19012 5728 19068
rect 5664 19008 5728 19012
rect 5744 19068 5808 19072
rect 5744 19012 5748 19068
rect 5748 19012 5804 19068
rect 5804 19012 5808 19068
rect 5744 19008 5808 19012
rect 5824 19068 5888 19072
rect 5824 19012 5828 19068
rect 5828 19012 5884 19068
rect 5884 19012 5888 19068
rect 5824 19008 5888 19012
rect 14848 19068 14912 19072
rect 14848 19012 14852 19068
rect 14852 19012 14908 19068
rect 14908 19012 14912 19068
rect 14848 19008 14912 19012
rect 14928 19068 14992 19072
rect 14928 19012 14932 19068
rect 14932 19012 14988 19068
rect 14988 19012 14992 19068
rect 14928 19008 14992 19012
rect 15008 19068 15072 19072
rect 15008 19012 15012 19068
rect 15012 19012 15068 19068
rect 15068 19012 15072 19068
rect 15008 19008 15072 19012
rect 15088 19068 15152 19072
rect 15088 19012 15092 19068
rect 15092 19012 15148 19068
rect 15148 19012 15152 19068
rect 15088 19008 15152 19012
rect 24112 19068 24176 19072
rect 24112 19012 24116 19068
rect 24116 19012 24172 19068
rect 24172 19012 24176 19068
rect 24112 19008 24176 19012
rect 24192 19068 24256 19072
rect 24192 19012 24196 19068
rect 24196 19012 24252 19068
rect 24252 19012 24256 19068
rect 24192 19008 24256 19012
rect 24272 19068 24336 19072
rect 24272 19012 24276 19068
rect 24276 19012 24332 19068
rect 24332 19012 24336 19068
rect 24272 19008 24336 19012
rect 24352 19068 24416 19072
rect 24352 19012 24356 19068
rect 24356 19012 24412 19068
rect 24412 19012 24416 19068
rect 24352 19008 24416 19012
rect 10216 18524 10280 18528
rect 10216 18468 10220 18524
rect 10220 18468 10276 18524
rect 10276 18468 10280 18524
rect 10216 18464 10280 18468
rect 10296 18524 10360 18528
rect 10296 18468 10300 18524
rect 10300 18468 10356 18524
rect 10356 18468 10360 18524
rect 10296 18464 10360 18468
rect 10376 18524 10440 18528
rect 10376 18468 10380 18524
rect 10380 18468 10436 18524
rect 10436 18468 10440 18524
rect 10376 18464 10440 18468
rect 10456 18524 10520 18528
rect 10456 18468 10460 18524
rect 10460 18468 10516 18524
rect 10516 18468 10520 18524
rect 10456 18464 10520 18468
rect 19480 18524 19544 18528
rect 19480 18468 19484 18524
rect 19484 18468 19540 18524
rect 19540 18468 19544 18524
rect 19480 18464 19544 18468
rect 19560 18524 19624 18528
rect 19560 18468 19564 18524
rect 19564 18468 19620 18524
rect 19620 18468 19624 18524
rect 19560 18464 19624 18468
rect 19640 18524 19704 18528
rect 19640 18468 19644 18524
rect 19644 18468 19700 18524
rect 19700 18468 19704 18524
rect 19640 18464 19704 18468
rect 19720 18524 19784 18528
rect 19720 18468 19724 18524
rect 19724 18468 19780 18524
rect 19780 18468 19784 18524
rect 19720 18464 19784 18468
rect 5584 17980 5648 17984
rect 5584 17924 5588 17980
rect 5588 17924 5644 17980
rect 5644 17924 5648 17980
rect 5584 17920 5648 17924
rect 5664 17980 5728 17984
rect 5664 17924 5668 17980
rect 5668 17924 5724 17980
rect 5724 17924 5728 17980
rect 5664 17920 5728 17924
rect 5744 17980 5808 17984
rect 5744 17924 5748 17980
rect 5748 17924 5804 17980
rect 5804 17924 5808 17980
rect 5744 17920 5808 17924
rect 5824 17980 5888 17984
rect 5824 17924 5828 17980
rect 5828 17924 5884 17980
rect 5884 17924 5888 17980
rect 5824 17920 5888 17924
rect 14848 17980 14912 17984
rect 14848 17924 14852 17980
rect 14852 17924 14908 17980
rect 14908 17924 14912 17980
rect 14848 17920 14912 17924
rect 14928 17980 14992 17984
rect 14928 17924 14932 17980
rect 14932 17924 14988 17980
rect 14988 17924 14992 17980
rect 14928 17920 14992 17924
rect 15008 17980 15072 17984
rect 15008 17924 15012 17980
rect 15012 17924 15068 17980
rect 15068 17924 15072 17980
rect 15008 17920 15072 17924
rect 15088 17980 15152 17984
rect 15088 17924 15092 17980
rect 15092 17924 15148 17980
rect 15148 17924 15152 17980
rect 15088 17920 15152 17924
rect 24112 17980 24176 17984
rect 24112 17924 24116 17980
rect 24116 17924 24172 17980
rect 24172 17924 24176 17980
rect 24112 17920 24176 17924
rect 24192 17980 24256 17984
rect 24192 17924 24196 17980
rect 24196 17924 24252 17980
rect 24252 17924 24256 17980
rect 24192 17920 24256 17924
rect 24272 17980 24336 17984
rect 24272 17924 24276 17980
rect 24276 17924 24332 17980
rect 24332 17924 24336 17980
rect 24272 17920 24336 17924
rect 24352 17980 24416 17984
rect 24352 17924 24356 17980
rect 24356 17924 24412 17980
rect 24412 17924 24416 17980
rect 24352 17920 24416 17924
rect 10216 17436 10280 17440
rect 10216 17380 10220 17436
rect 10220 17380 10276 17436
rect 10276 17380 10280 17436
rect 10216 17376 10280 17380
rect 10296 17436 10360 17440
rect 10296 17380 10300 17436
rect 10300 17380 10356 17436
rect 10356 17380 10360 17436
rect 10296 17376 10360 17380
rect 10376 17436 10440 17440
rect 10376 17380 10380 17436
rect 10380 17380 10436 17436
rect 10436 17380 10440 17436
rect 10376 17376 10440 17380
rect 10456 17436 10520 17440
rect 10456 17380 10460 17436
rect 10460 17380 10516 17436
rect 10516 17380 10520 17436
rect 10456 17376 10520 17380
rect 19480 17436 19544 17440
rect 19480 17380 19484 17436
rect 19484 17380 19540 17436
rect 19540 17380 19544 17436
rect 19480 17376 19544 17380
rect 19560 17436 19624 17440
rect 19560 17380 19564 17436
rect 19564 17380 19620 17436
rect 19620 17380 19624 17436
rect 19560 17376 19624 17380
rect 19640 17436 19704 17440
rect 19640 17380 19644 17436
rect 19644 17380 19700 17436
rect 19700 17380 19704 17436
rect 19640 17376 19704 17380
rect 19720 17436 19784 17440
rect 19720 17380 19724 17436
rect 19724 17380 19780 17436
rect 19780 17380 19784 17436
rect 19720 17376 19784 17380
rect 5584 16892 5648 16896
rect 5584 16836 5588 16892
rect 5588 16836 5644 16892
rect 5644 16836 5648 16892
rect 5584 16832 5648 16836
rect 5664 16892 5728 16896
rect 5664 16836 5668 16892
rect 5668 16836 5724 16892
rect 5724 16836 5728 16892
rect 5664 16832 5728 16836
rect 5744 16892 5808 16896
rect 5744 16836 5748 16892
rect 5748 16836 5804 16892
rect 5804 16836 5808 16892
rect 5744 16832 5808 16836
rect 5824 16892 5888 16896
rect 5824 16836 5828 16892
rect 5828 16836 5884 16892
rect 5884 16836 5888 16892
rect 5824 16832 5888 16836
rect 14848 16892 14912 16896
rect 14848 16836 14852 16892
rect 14852 16836 14908 16892
rect 14908 16836 14912 16892
rect 14848 16832 14912 16836
rect 14928 16892 14992 16896
rect 14928 16836 14932 16892
rect 14932 16836 14988 16892
rect 14988 16836 14992 16892
rect 14928 16832 14992 16836
rect 15008 16892 15072 16896
rect 15008 16836 15012 16892
rect 15012 16836 15068 16892
rect 15068 16836 15072 16892
rect 15008 16832 15072 16836
rect 15088 16892 15152 16896
rect 15088 16836 15092 16892
rect 15092 16836 15148 16892
rect 15148 16836 15152 16892
rect 15088 16832 15152 16836
rect 24112 16892 24176 16896
rect 24112 16836 24116 16892
rect 24116 16836 24172 16892
rect 24172 16836 24176 16892
rect 24112 16832 24176 16836
rect 24192 16892 24256 16896
rect 24192 16836 24196 16892
rect 24196 16836 24252 16892
rect 24252 16836 24256 16892
rect 24192 16832 24256 16836
rect 24272 16892 24336 16896
rect 24272 16836 24276 16892
rect 24276 16836 24332 16892
rect 24332 16836 24336 16892
rect 24272 16832 24336 16836
rect 24352 16892 24416 16896
rect 24352 16836 24356 16892
rect 24356 16836 24412 16892
rect 24412 16836 24416 16892
rect 24352 16832 24416 16836
rect 10216 16348 10280 16352
rect 10216 16292 10220 16348
rect 10220 16292 10276 16348
rect 10276 16292 10280 16348
rect 10216 16288 10280 16292
rect 10296 16348 10360 16352
rect 10296 16292 10300 16348
rect 10300 16292 10356 16348
rect 10356 16292 10360 16348
rect 10296 16288 10360 16292
rect 10376 16348 10440 16352
rect 10376 16292 10380 16348
rect 10380 16292 10436 16348
rect 10436 16292 10440 16348
rect 10376 16288 10440 16292
rect 10456 16348 10520 16352
rect 10456 16292 10460 16348
rect 10460 16292 10516 16348
rect 10516 16292 10520 16348
rect 10456 16288 10520 16292
rect 19480 16348 19544 16352
rect 19480 16292 19484 16348
rect 19484 16292 19540 16348
rect 19540 16292 19544 16348
rect 19480 16288 19544 16292
rect 19560 16348 19624 16352
rect 19560 16292 19564 16348
rect 19564 16292 19620 16348
rect 19620 16292 19624 16348
rect 19560 16288 19624 16292
rect 19640 16348 19704 16352
rect 19640 16292 19644 16348
rect 19644 16292 19700 16348
rect 19700 16292 19704 16348
rect 19640 16288 19704 16292
rect 19720 16348 19784 16352
rect 19720 16292 19724 16348
rect 19724 16292 19780 16348
rect 19780 16292 19784 16348
rect 19720 16288 19784 16292
rect 5584 15804 5648 15808
rect 5584 15748 5588 15804
rect 5588 15748 5644 15804
rect 5644 15748 5648 15804
rect 5584 15744 5648 15748
rect 5664 15804 5728 15808
rect 5664 15748 5668 15804
rect 5668 15748 5724 15804
rect 5724 15748 5728 15804
rect 5664 15744 5728 15748
rect 5744 15804 5808 15808
rect 5744 15748 5748 15804
rect 5748 15748 5804 15804
rect 5804 15748 5808 15804
rect 5744 15744 5808 15748
rect 5824 15804 5888 15808
rect 5824 15748 5828 15804
rect 5828 15748 5884 15804
rect 5884 15748 5888 15804
rect 5824 15744 5888 15748
rect 14848 15804 14912 15808
rect 14848 15748 14852 15804
rect 14852 15748 14908 15804
rect 14908 15748 14912 15804
rect 14848 15744 14912 15748
rect 14928 15804 14992 15808
rect 14928 15748 14932 15804
rect 14932 15748 14988 15804
rect 14988 15748 14992 15804
rect 14928 15744 14992 15748
rect 15008 15804 15072 15808
rect 15008 15748 15012 15804
rect 15012 15748 15068 15804
rect 15068 15748 15072 15804
rect 15008 15744 15072 15748
rect 15088 15804 15152 15808
rect 15088 15748 15092 15804
rect 15092 15748 15148 15804
rect 15148 15748 15152 15804
rect 15088 15744 15152 15748
rect 24112 15804 24176 15808
rect 24112 15748 24116 15804
rect 24116 15748 24172 15804
rect 24172 15748 24176 15804
rect 24112 15744 24176 15748
rect 24192 15804 24256 15808
rect 24192 15748 24196 15804
rect 24196 15748 24252 15804
rect 24252 15748 24256 15804
rect 24192 15744 24256 15748
rect 24272 15804 24336 15808
rect 24272 15748 24276 15804
rect 24276 15748 24332 15804
rect 24332 15748 24336 15804
rect 24272 15744 24336 15748
rect 24352 15804 24416 15808
rect 24352 15748 24356 15804
rect 24356 15748 24412 15804
rect 24412 15748 24416 15804
rect 24352 15744 24416 15748
rect 10216 15260 10280 15264
rect 10216 15204 10220 15260
rect 10220 15204 10276 15260
rect 10276 15204 10280 15260
rect 10216 15200 10280 15204
rect 10296 15260 10360 15264
rect 10296 15204 10300 15260
rect 10300 15204 10356 15260
rect 10356 15204 10360 15260
rect 10296 15200 10360 15204
rect 10376 15260 10440 15264
rect 10376 15204 10380 15260
rect 10380 15204 10436 15260
rect 10436 15204 10440 15260
rect 10376 15200 10440 15204
rect 10456 15260 10520 15264
rect 10456 15204 10460 15260
rect 10460 15204 10516 15260
rect 10516 15204 10520 15260
rect 10456 15200 10520 15204
rect 19480 15260 19544 15264
rect 19480 15204 19484 15260
rect 19484 15204 19540 15260
rect 19540 15204 19544 15260
rect 19480 15200 19544 15204
rect 19560 15260 19624 15264
rect 19560 15204 19564 15260
rect 19564 15204 19620 15260
rect 19620 15204 19624 15260
rect 19560 15200 19624 15204
rect 19640 15260 19704 15264
rect 19640 15204 19644 15260
rect 19644 15204 19700 15260
rect 19700 15204 19704 15260
rect 19640 15200 19704 15204
rect 19720 15260 19784 15264
rect 19720 15204 19724 15260
rect 19724 15204 19780 15260
rect 19780 15204 19784 15260
rect 19720 15200 19784 15204
rect 5584 14716 5648 14720
rect 5584 14660 5588 14716
rect 5588 14660 5644 14716
rect 5644 14660 5648 14716
rect 5584 14656 5648 14660
rect 5664 14716 5728 14720
rect 5664 14660 5668 14716
rect 5668 14660 5724 14716
rect 5724 14660 5728 14716
rect 5664 14656 5728 14660
rect 5744 14716 5808 14720
rect 5744 14660 5748 14716
rect 5748 14660 5804 14716
rect 5804 14660 5808 14716
rect 5744 14656 5808 14660
rect 5824 14716 5888 14720
rect 5824 14660 5828 14716
rect 5828 14660 5884 14716
rect 5884 14660 5888 14716
rect 5824 14656 5888 14660
rect 14848 14716 14912 14720
rect 14848 14660 14852 14716
rect 14852 14660 14908 14716
rect 14908 14660 14912 14716
rect 14848 14656 14912 14660
rect 14928 14716 14992 14720
rect 14928 14660 14932 14716
rect 14932 14660 14988 14716
rect 14988 14660 14992 14716
rect 14928 14656 14992 14660
rect 15008 14716 15072 14720
rect 15008 14660 15012 14716
rect 15012 14660 15068 14716
rect 15068 14660 15072 14716
rect 15008 14656 15072 14660
rect 15088 14716 15152 14720
rect 15088 14660 15092 14716
rect 15092 14660 15148 14716
rect 15148 14660 15152 14716
rect 15088 14656 15152 14660
rect 24112 14716 24176 14720
rect 24112 14660 24116 14716
rect 24116 14660 24172 14716
rect 24172 14660 24176 14716
rect 24112 14656 24176 14660
rect 24192 14716 24256 14720
rect 24192 14660 24196 14716
rect 24196 14660 24252 14716
rect 24252 14660 24256 14716
rect 24192 14656 24256 14660
rect 24272 14716 24336 14720
rect 24272 14660 24276 14716
rect 24276 14660 24332 14716
rect 24332 14660 24336 14716
rect 24272 14656 24336 14660
rect 24352 14716 24416 14720
rect 24352 14660 24356 14716
rect 24356 14660 24412 14716
rect 24412 14660 24416 14716
rect 24352 14656 24416 14660
rect 10216 14172 10280 14176
rect 10216 14116 10220 14172
rect 10220 14116 10276 14172
rect 10276 14116 10280 14172
rect 10216 14112 10280 14116
rect 10296 14172 10360 14176
rect 10296 14116 10300 14172
rect 10300 14116 10356 14172
rect 10356 14116 10360 14172
rect 10296 14112 10360 14116
rect 10376 14172 10440 14176
rect 10376 14116 10380 14172
rect 10380 14116 10436 14172
rect 10436 14116 10440 14172
rect 10376 14112 10440 14116
rect 10456 14172 10520 14176
rect 10456 14116 10460 14172
rect 10460 14116 10516 14172
rect 10516 14116 10520 14172
rect 10456 14112 10520 14116
rect 19480 14172 19544 14176
rect 19480 14116 19484 14172
rect 19484 14116 19540 14172
rect 19540 14116 19544 14172
rect 19480 14112 19544 14116
rect 19560 14172 19624 14176
rect 19560 14116 19564 14172
rect 19564 14116 19620 14172
rect 19620 14116 19624 14172
rect 19560 14112 19624 14116
rect 19640 14172 19704 14176
rect 19640 14116 19644 14172
rect 19644 14116 19700 14172
rect 19700 14116 19704 14172
rect 19640 14112 19704 14116
rect 19720 14172 19784 14176
rect 19720 14116 19724 14172
rect 19724 14116 19780 14172
rect 19780 14116 19784 14172
rect 19720 14112 19784 14116
rect 27476 13908 27540 13972
rect 5584 13628 5648 13632
rect 5584 13572 5588 13628
rect 5588 13572 5644 13628
rect 5644 13572 5648 13628
rect 5584 13568 5648 13572
rect 5664 13628 5728 13632
rect 5664 13572 5668 13628
rect 5668 13572 5724 13628
rect 5724 13572 5728 13628
rect 5664 13568 5728 13572
rect 5744 13628 5808 13632
rect 5744 13572 5748 13628
rect 5748 13572 5804 13628
rect 5804 13572 5808 13628
rect 5744 13568 5808 13572
rect 5824 13628 5888 13632
rect 5824 13572 5828 13628
rect 5828 13572 5884 13628
rect 5884 13572 5888 13628
rect 5824 13568 5888 13572
rect 14848 13628 14912 13632
rect 14848 13572 14852 13628
rect 14852 13572 14908 13628
rect 14908 13572 14912 13628
rect 14848 13568 14912 13572
rect 14928 13628 14992 13632
rect 14928 13572 14932 13628
rect 14932 13572 14988 13628
rect 14988 13572 14992 13628
rect 14928 13568 14992 13572
rect 15008 13628 15072 13632
rect 15008 13572 15012 13628
rect 15012 13572 15068 13628
rect 15068 13572 15072 13628
rect 15008 13568 15072 13572
rect 15088 13628 15152 13632
rect 15088 13572 15092 13628
rect 15092 13572 15148 13628
rect 15148 13572 15152 13628
rect 15088 13568 15152 13572
rect 24112 13628 24176 13632
rect 24112 13572 24116 13628
rect 24116 13572 24172 13628
rect 24172 13572 24176 13628
rect 24112 13568 24176 13572
rect 24192 13628 24256 13632
rect 24192 13572 24196 13628
rect 24196 13572 24252 13628
rect 24252 13572 24256 13628
rect 24192 13568 24256 13572
rect 24272 13628 24336 13632
rect 24272 13572 24276 13628
rect 24276 13572 24332 13628
rect 24332 13572 24336 13628
rect 24272 13568 24336 13572
rect 24352 13628 24416 13632
rect 24352 13572 24356 13628
rect 24356 13572 24412 13628
rect 24412 13572 24416 13628
rect 24352 13568 24416 13572
rect 10216 13084 10280 13088
rect 10216 13028 10220 13084
rect 10220 13028 10276 13084
rect 10276 13028 10280 13084
rect 10216 13024 10280 13028
rect 10296 13084 10360 13088
rect 10296 13028 10300 13084
rect 10300 13028 10356 13084
rect 10356 13028 10360 13084
rect 10296 13024 10360 13028
rect 10376 13084 10440 13088
rect 10376 13028 10380 13084
rect 10380 13028 10436 13084
rect 10436 13028 10440 13084
rect 10376 13024 10440 13028
rect 10456 13084 10520 13088
rect 10456 13028 10460 13084
rect 10460 13028 10516 13084
rect 10516 13028 10520 13084
rect 10456 13024 10520 13028
rect 19480 13084 19544 13088
rect 19480 13028 19484 13084
rect 19484 13028 19540 13084
rect 19540 13028 19544 13084
rect 19480 13024 19544 13028
rect 19560 13084 19624 13088
rect 19560 13028 19564 13084
rect 19564 13028 19620 13084
rect 19620 13028 19624 13084
rect 19560 13024 19624 13028
rect 19640 13084 19704 13088
rect 19640 13028 19644 13084
rect 19644 13028 19700 13084
rect 19700 13028 19704 13084
rect 19640 13024 19704 13028
rect 19720 13084 19784 13088
rect 19720 13028 19724 13084
rect 19724 13028 19780 13084
rect 19780 13028 19784 13084
rect 19720 13024 19784 13028
rect 5584 12540 5648 12544
rect 5584 12484 5588 12540
rect 5588 12484 5644 12540
rect 5644 12484 5648 12540
rect 5584 12480 5648 12484
rect 5664 12540 5728 12544
rect 5664 12484 5668 12540
rect 5668 12484 5724 12540
rect 5724 12484 5728 12540
rect 5664 12480 5728 12484
rect 5744 12540 5808 12544
rect 5744 12484 5748 12540
rect 5748 12484 5804 12540
rect 5804 12484 5808 12540
rect 5744 12480 5808 12484
rect 5824 12540 5888 12544
rect 5824 12484 5828 12540
rect 5828 12484 5884 12540
rect 5884 12484 5888 12540
rect 5824 12480 5888 12484
rect 14848 12540 14912 12544
rect 14848 12484 14852 12540
rect 14852 12484 14908 12540
rect 14908 12484 14912 12540
rect 14848 12480 14912 12484
rect 14928 12540 14992 12544
rect 14928 12484 14932 12540
rect 14932 12484 14988 12540
rect 14988 12484 14992 12540
rect 14928 12480 14992 12484
rect 15008 12540 15072 12544
rect 15008 12484 15012 12540
rect 15012 12484 15068 12540
rect 15068 12484 15072 12540
rect 15008 12480 15072 12484
rect 15088 12540 15152 12544
rect 15088 12484 15092 12540
rect 15092 12484 15148 12540
rect 15148 12484 15152 12540
rect 15088 12480 15152 12484
rect 24112 12540 24176 12544
rect 24112 12484 24116 12540
rect 24116 12484 24172 12540
rect 24172 12484 24176 12540
rect 24112 12480 24176 12484
rect 24192 12540 24256 12544
rect 24192 12484 24196 12540
rect 24196 12484 24252 12540
rect 24252 12484 24256 12540
rect 24192 12480 24256 12484
rect 24272 12540 24336 12544
rect 24272 12484 24276 12540
rect 24276 12484 24332 12540
rect 24332 12484 24336 12540
rect 24272 12480 24336 12484
rect 24352 12540 24416 12544
rect 24352 12484 24356 12540
rect 24356 12484 24412 12540
rect 24412 12484 24416 12540
rect 24352 12480 24416 12484
rect 10216 11996 10280 12000
rect 10216 11940 10220 11996
rect 10220 11940 10276 11996
rect 10276 11940 10280 11996
rect 10216 11936 10280 11940
rect 10296 11996 10360 12000
rect 10296 11940 10300 11996
rect 10300 11940 10356 11996
rect 10356 11940 10360 11996
rect 10296 11936 10360 11940
rect 10376 11996 10440 12000
rect 10376 11940 10380 11996
rect 10380 11940 10436 11996
rect 10436 11940 10440 11996
rect 10376 11936 10440 11940
rect 10456 11996 10520 12000
rect 10456 11940 10460 11996
rect 10460 11940 10516 11996
rect 10516 11940 10520 11996
rect 10456 11936 10520 11940
rect 19480 11996 19544 12000
rect 19480 11940 19484 11996
rect 19484 11940 19540 11996
rect 19540 11940 19544 11996
rect 19480 11936 19544 11940
rect 19560 11996 19624 12000
rect 19560 11940 19564 11996
rect 19564 11940 19620 11996
rect 19620 11940 19624 11996
rect 19560 11936 19624 11940
rect 19640 11996 19704 12000
rect 19640 11940 19644 11996
rect 19644 11940 19700 11996
rect 19700 11940 19704 11996
rect 19640 11936 19704 11940
rect 19720 11996 19784 12000
rect 19720 11940 19724 11996
rect 19724 11940 19780 11996
rect 19780 11940 19784 11996
rect 19720 11936 19784 11940
rect 5584 11452 5648 11456
rect 5584 11396 5588 11452
rect 5588 11396 5644 11452
rect 5644 11396 5648 11452
rect 5584 11392 5648 11396
rect 5664 11452 5728 11456
rect 5664 11396 5668 11452
rect 5668 11396 5724 11452
rect 5724 11396 5728 11452
rect 5664 11392 5728 11396
rect 5744 11452 5808 11456
rect 5744 11396 5748 11452
rect 5748 11396 5804 11452
rect 5804 11396 5808 11452
rect 5744 11392 5808 11396
rect 5824 11452 5888 11456
rect 5824 11396 5828 11452
rect 5828 11396 5884 11452
rect 5884 11396 5888 11452
rect 5824 11392 5888 11396
rect 14848 11452 14912 11456
rect 14848 11396 14852 11452
rect 14852 11396 14908 11452
rect 14908 11396 14912 11452
rect 14848 11392 14912 11396
rect 14928 11452 14992 11456
rect 14928 11396 14932 11452
rect 14932 11396 14988 11452
rect 14988 11396 14992 11452
rect 14928 11392 14992 11396
rect 15008 11452 15072 11456
rect 15008 11396 15012 11452
rect 15012 11396 15068 11452
rect 15068 11396 15072 11452
rect 15008 11392 15072 11396
rect 15088 11452 15152 11456
rect 15088 11396 15092 11452
rect 15092 11396 15148 11452
rect 15148 11396 15152 11452
rect 15088 11392 15152 11396
rect 24112 11452 24176 11456
rect 24112 11396 24116 11452
rect 24116 11396 24172 11452
rect 24172 11396 24176 11452
rect 24112 11392 24176 11396
rect 24192 11452 24256 11456
rect 24192 11396 24196 11452
rect 24196 11396 24252 11452
rect 24252 11396 24256 11452
rect 24192 11392 24256 11396
rect 24272 11452 24336 11456
rect 24272 11396 24276 11452
rect 24276 11396 24332 11452
rect 24332 11396 24336 11452
rect 24272 11392 24336 11396
rect 24352 11452 24416 11456
rect 24352 11396 24356 11452
rect 24356 11396 24412 11452
rect 24412 11396 24416 11452
rect 24352 11392 24416 11396
rect 10216 10908 10280 10912
rect 10216 10852 10220 10908
rect 10220 10852 10276 10908
rect 10276 10852 10280 10908
rect 10216 10848 10280 10852
rect 10296 10908 10360 10912
rect 10296 10852 10300 10908
rect 10300 10852 10356 10908
rect 10356 10852 10360 10908
rect 10296 10848 10360 10852
rect 10376 10908 10440 10912
rect 10376 10852 10380 10908
rect 10380 10852 10436 10908
rect 10436 10852 10440 10908
rect 10376 10848 10440 10852
rect 10456 10908 10520 10912
rect 10456 10852 10460 10908
rect 10460 10852 10516 10908
rect 10516 10852 10520 10908
rect 10456 10848 10520 10852
rect 19480 10908 19544 10912
rect 19480 10852 19484 10908
rect 19484 10852 19540 10908
rect 19540 10852 19544 10908
rect 19480 10848 19544 10852
rect 19560 10908 19624 10912
rect 19560 10852 19564 10908
rect 19564 10852 19620 10908
rect 19620 10852 19624 10908
rect 19560 10848 19624 10852
rect 19640 10908 19704 10912
rect 19640 10852 19644 10908
rect 19644 10852 19700 10908
rect 19700 10852 19704 10908
rect 19640 10848 19704 10852
rect 19720 10908 19784 10912
rect 19720 10852 19724 10908
rect 19724 10852 19780 10908
rect 19780 10852 19784 10908
rect 19720 10848 19784 10852
rect 5584 10364 5648 10368
rect 5584 10308 5588 10364
rect 5588 10308 5644 10364
rect 5644 10308 5648 10364
rect 5584 10304 5648 10308
rect 5664 10364 5728 10368
rect 5664 10308 5668 10364
rect 5668 10308 5724 10364
rect 5724 10308 5728 10364
rect 5664 10304 5728 10308
rect 5744 10364 5808 10368
rect 5744 10308 5748 10364
rect 5748 10308 5804 10364
rect 5804 10308 5808 10364
rect 5744 10304 5808 10308
rect 5824 10364 5888 10368
rect 5824 10308 5828 10364
rect 5828 10308 5884 10364
rect 5884 10308 5888 10364
rect 5824 10304 5888 10308
rect 14848 10364 14912 10368
rect 14848 10308 14852 10364
rect 14852 10308 14908 10364
rect 14908 10308 14912 10364
rect 14848 10304 14912 10308
rect 14928 10364 14992 10368
rect 14928 10308 14932 10364
rect 14932 10308 14988 10364
rect 14988 10308 14992 10364
rect 14928 10304 14992 10308
rect 15008 10364 15072 10368
rect 15008 10308 15012 10364
rect 15012 10308 15068 10364
rect 15068 10308 15072 10364
rect 15008 10304 15072 10308
rect 15088 10364 15152 10368
rect 15088 10308 15092 10364
rect 15092 10308 15148 10364
rect 15148 10308 15152 10364
rect 15088 10304 15152 10308
rect 24112 10364 24176 10368
rect 24112 10308 24116 10364
rect 24116 10308 24172 10364
rect 24172 10308 24176 10364
rect 24112 10304 24176 10308
rect 24192 10364 24256 10368
rect 24192 10308 24196 10364
rect 24196 10308 24252 10364
rect 24252 10308 24256 10364
rect 24192 10304 24256 10308
rect 24272 10364 24336 10368
rect 24272 10308 24276 10364
rect 24276 10308 24332 10364
rect 24332 10308 24336 10364
rect 24272 10304 24336 10308
rect 24352 10364 24416 10368
rect 24352 10308 24356 10364
rect 24356 10308 24412 10364
rect 24412 10308 24416 10364
rect 24352 10304 24416 10308
rect 10216 9820 10280 9824
rect 10216 9764 10220 9820
rect 10220 9764 10276 9820
rect 10276 9764 10280 9820
rect 10216 9760 10280 9764
rect 10296 9820 10360 9824
rect 10296 9764 10300 9820
rect 10300 9764 10356 9820
rect 10356 9764 10360 9820
rect 10296 9760 10360 9764
rect 10376 9820 10440 9824
rect 10376 9764 10380 9820
rect 10380 9764 10436 9820
rect 10436 9764 10440 9820
rect 10376 9760 10440 9764
rect 10456 9820 10520 9824
rect 10456 9764 10460 9820
rect 10460 9764 10516 9820
rect 10516 9764 10520 9820
rect 10456 9760 10520 9764
rect 19480 9820 19544 9824
rect 19480 9764 19484 9820
rect 19484 9764 19540 9820
rect 19540 9764 19544 9820
rect 19480 9760 19544 9764
rect 19560 9820 19624 9824
rect 19560 9764 19564 9820
rect 19564 9764 19620 9820
rect 19620 9764 19624 9820
rect 19560 9760 19624 9764
rect 19640 9820 19704 9824
rect 19640 9764 19644 9820
rect 19644 9764 19700 9820
rect 19700 9764 19704 9820
rect 19640 9760 19704 9764
rect 19720 9820 19784 9824
rect 19720 9764 19724 9820
rect 19724 9764 19780 9820
rect 19780 9764 19784 9820
rect 19720 9760 19784 9764
rect 5584 9276 5648 9280
rect 5584 9220 5588 9276
rect 5588 9220 5644 9276
rect 5644 9220 5648 9276
rect 5584 9216 5648 9220
rect 5664 9276 5728 9280
rect 5664 9220 5668 9276
rect 5668 9220 5724 9276
rect 5724 9220 5728 9276
rect 5664 9216 5728 9220
rect 5744 9276 5808 9280
rect 5744 9220 5748 9276
rect 5748 9220 5804 9276
rect 5804 9220 5808 9276
rect 5744 9216 5808 9220
rect 5824 9276 5888 9280
rect 5824 9220 5828 9276
rect 5828 9220 5884 9276
rect 5884 9220 5888 9276
rect 5824 9216 5888 9220
rect 14848 9276 14912 9280
rect 14848 9220 14852 9276
rect 14852 9220 14908 9276
rect 14908 9220 14912 9276
rect 14848 9216 14912 9220
rect 14928 9276 14992 9280
rect 14928 9220 14932 9276
rect 14932 9220 14988 9276
rect 14988 9220 14992 9276
rect 14928 9216 14992 9220
rect 15008 9276 15072 9280
rect 15008 9220 15012 9276
rect 15012 9220 15068 9276
rect 15068 9220 15072 9276
rect 15008 9216 15072 9220
rect 15088 9276 15152 9280
rect 15088 9220 15092 9276
rect 15092 9220 15148 9276
rect 15148 9220 15152 9276
rect 15088 9216 15152 9220
rect 24112 9276 24176 9280
rect 24112 9220 24116 9276
rect 24116 9220 24172 9276
rect 24172 9220 24176 9276
rect 24112 9216 24176 9220
rect 24192 9276 24256 9280
rect 24192 9220 24196 9276
rect 24196 9220 24252 9276
rect 24252 9220 24256 9276
rect 24192 9216 24256 9220
rect 24272 9276 24336 9280
rect 24272 9220 24276 9276
rect 24276 9220 24332 9276
rect 24332 9220 24336 9276
rect 24272 9216 24336 9220
rect 24352 9276 24416 9280
rect 24352 9220 24356 9276
rect 24356 9220 24412 9276
rect 24412 9220 24416 9276
rect 24352 9216 24416 9220
rect 10216 8732 10280 8736
rect 10216 8676 10220 8732
rect 10220 8676 10276 8732
rect 10276 8676 10280 8732
rect 10216 8672 10280 8676
rect 10296 8732 10360 8736
rect 10296 8676 10300 8732
rect 10300 8676 10356 8732
rect 10356 8676 10360 8732
rect 10296 8672 10360 8676
rect 10376 8732 10440 8736
rect 10376 8676 10380 8732
rect 10380 8676 10436 8732
rect 10436 8676 10440 8732
rect 10376 8672 10440 8676
rect 10456 8732 10520 8736
rect 10456 8676 10460 8732
rect 10460 8676 10516 8732
rect 10516 8676 10520 8732
rect 10456 8672 10520 8676
rect 19480 8732 19544 8736
rect 19480 8676 19484 8732
rect 19484 8676 19540 8732
rect 19540 8676 19544 8732
rect 19480 8672 19544 8676
rect 19560 8732 19624 8736
rect 19560 8676 19564 8732
rect 19564 8676 19620 8732
rect 19620 8676 19624 8732
rect 19560 8672 19624 8676
rect 19640 8732 19704 8736
rect 19640 8676 19644 8732
rect 19644 8676 19700 8732
rect 19700 8676 19704 8732
rect 19640 8672 19704 8676
rect 19720 8732 19784 8736
rect 19720 8676 19724 8732
rect 19724 8676 19780 8732
rect 19780 8676 19784 8732
rect 19720 8672 19784 8676
rect 5584 8188 5648 8192
rect 5584 8132 5588 8188
rect 5588 8132 5644 8188
rect 5644 8132 5648 8188
rect 5584 8128 5648 8132
rect 5664 8188 5728 8192
rect 5664 8132 5668 8188
rect 5668 8132 5724 8188
rect 5724 8132 5728 8188
rect 5664 8128 5728 8132
rect 5744 8188 5808 8192
rect 5744 8132 5748 8188
rect 5748 8132 5804 8188
rect 5804 8132 5808 8188
rect 5744 8128 5808 8132
rect 5824 8188 5888 8192
rect 5824 8132 5828 8188
rect 5828 8132 5884 8188
rect 5884 8132 5888 8188
rect 5824 8128 5888 8132
rect 14848 8188 14912 8192
rect 14848 8132 14852 8188
rect 14852 8132 14908 8188
rect 14908 8132 14912 8188
rect 14848 8128 14912 8132
rect 14928 8188 14992 8192
rect 14928 8132 14932 8188
rect 14932 8132 14988 8188
rect 14988 8132 14992 8188
rect 14928 8128 14992 8132
rect 15008 8188 15072 8192
rect 15008 8132 15012 8188
rect 15012 8132 15068 8188
rect 15068 8132 15072 8188
rect 15008 8128 15072 8132
rect 15088 8188 15152 8192
rect 15088 8132 15092 8188
rect 15092 8132 15148 8188
rect 15148 8132 15152 8188
rect 15088 8128 15152 8132
rect 24112 8188 24176 8192
rect 24112 8132 24116 8188
rect 24116 8132 24172 8188
rect 24172 8132 24176 8188
rect 24112 8128 24176 8132
rect 24192 8188 24256 8192
rect 24192 8132 24196 8188
rect 24196 8132 24252 8188
rect 24252 8132 24256 8188
rect 24192 8128 24256 8132
rect 24272 8188 24336 8192
rect 24272 8132 24276 8188
rect 24276 8132 24332 8188
rect 24332 8132 24336 8188
rect 24272 8128 24336 8132
rect 24352 8188 24416 8192
rect 24352 8132 24356 8188
rect 24356 8132 24412 8188
rect 24412 8132 24416 8188
rect 24352 8128 24416 8132
rect 18644 7984 18708 7988
rect 18644 7928 18694 7984
rect 18694 7928 18708 7984
rect 18644 7924 18708 7928
rect 10216 7644 10280 7648
rect 10216 7588 10220 7644
rect 10220 7588 10276 7644
rect 10276 7588 10280 7644
rect 10216 7584 10280 7588
rect 10296 7644 10360 7648
rect 10296 7588 10300 7644
rect 10300 7588 10356 7644
rect 10356 7588 10360 7644
rect 10296 7584 10360 7588
rect 10376 7644 10440 7648
rect 10376 7588 10380 7644
rect 10380 7588 10436 7644
rect 10436 7588 10440 7644
rect 10376 7584 10440 7588
rect 10456 7644 10520 7648
rect 10456 7588 10460 7644
rect 10460 7588 10516 7644
rect 10516 7588 10520 7644
rect 10456 7584 10520 7588
rect 19480 7644 19544 7648
rect 19480 7588 19484 7644
rect 19484 7588 19540 7644
rect 19540 7588 19544 7644
rect 19480 7584 19544 7588
rect 19560 7644 19624 7648
rect 19560 7588 19564 7644
rect 19564 7588 19620 7644
rect 19620 7588 19624 7644
rect 19560 7584 19624 7588
rect 19640 7644 19704 7648
rect 19640 7588 19644 7644
rect 19644 7588 19700 7644
rect 19700 7588 19704 7644
rect 19640 7584 19704 7588
rect 19720 7644 19784 7648
rect 19720 7588 19724 7644
rect 19724 7588 19780 7644
rect 19780 7588 19784 7644
rect 19720 7584 19784 7588
rect 5584 7100 5648 7104
rect 5584 7044 5588 7100
rect 5588 7044 5644 7100
rect 5644 7044 5648 7100
rect 5584 7040 5648 7044
rect 5664 7100 5728 7104
rect 5664 7044 5668 7100
rect 5668 7044 5724 7100
rect 5724 7044 5728 7100
rect 5664 7040 5728 7044
rect 5744 7100 5808 7104
rect 5744 7044 5748 7100
rect 5748 7044 5804 7100
rect 5804 7044 5808 7100
rect 5744 7040 5808 7044
rect 5824 7100 5888 7104
rect 5824 7044 5828 7100
rect 5828 7044 5884 7100
rect 5884 7044 5888 7100
rect 5824 7040 5888 7044
rect 14848 7100 14912 7104
rect 14848 7044 14852 7100
rect 14852 7044 14908 7100
rect 14908 7044 14912 7100
rect 14848 7040 14912 7044
rect 14928 7100 14992 7104
rect 14928 7044 14932 7100
rect 14932 7044 14988 7100
rect 14988 7044 14992 7100
rect 14928 7040 14992 7044
rect 15008 7100 15072 7104
rect 15008 7044 15012 7100
rect 15012 7044 15068 7100
rect 15068 7044 15072 7100
rect 15008 7040 15072 7044
rect 15088 7100 15152 7104
rect 15088 7044 15092 7100
rect 15092 7044 15148 7100
rect 15148 7044 15152 7100
rect 15088 7040 15152 7044
rect 24112 7100 24176 7104
rect 24112 7044 24116 7100
rect 24116 7044 24172 7100
rect 24172 7044 24176 7100
rect 24112 7040 24176 7044
rect 24192 7100 24256 7104
rect 24192 7044 24196 7100
rect 24196 7044 24252 7100
rect 24252 7044 24256 7100
rect 24192 7040 24256 7044
rect 24272 7100 24336 7104
rect 24272 7044 24276 7100
rect 24276 7044 24332 7100
rect 24332 7044 24336 7100
rect 24272 7040 24336 7044
rect 24352 7100 24416 7104
rect 24352 7044 24356 7100
rect 24356 7044 24412 7100
rect 24412 7044 24416 7100
rect 24352 7040 24416 7044
rect 10216 6556 10280 6560
rect 10216 6500 10220 6556
rect 10220 6500 10276 6556
rect 10276 6500 10280 6556
rect 10216 6496 10280 6500
rect 10296 6556 10360 6560
rect 10296 6500 10300 6556
rect 10300 6500 10356 6556
rect 10356 6500 10360 6556
rect 10296 6496 10360 6500
rect 10376 6556 10440 6560
rect 10376 6500 10380 6556
rect 10380 6500 10436 6556
rect 10436 6500 10440 6556
rect 10376 6496 10440 6500
rect 10456 6556 10520 6560
rect 10456 6500 10460 6556
rect 10460 6500 10516 6556
rect 10516 6500 10520 6556
rect 10456 6496 10520 6500
rect 19480 6556 19544 6560
rect 19480 6500 19484 6556
rect 19484 6500 19540 6556
rect 19540 6500 19544 6556
rect 19480 6496 19544 6500
rect 19560 6556 19624 6560
rect 19560 6500 19564 6556
rect 19564 6500 19620 6556
rect 19620 6500 19624 6556
rect 19560 6496 19624 6500
rect 19640 6556 19704 6560
rect 19640 6500 19644 6556
rect 19644 6500 19700 6556
rect 19700 6500 19704 6556
rect 19640 6496 19704 6500
rect 19720 6556 19784 6560
rect 19720 6500 19724 6556
rect 19724 6500 19780 6556
rect 19780 6500 19784 6556
rect 19720 6496 19784 6500
rect 5584 6012 5648 6016
rect 5584 5956 5588 6012
rect 5588 5956 5644 6012
rect 5644 5956 5648 6012
rect 5584 5952 5648 5956
rect 5664 6012 5728 6016
rect 5664 5956 5668 6012
rect 5668 5956 5724 6012
rect 5724 5956 5728 6012
rect 5664 5952 5728 5956
rect 5744 6012 5808 6016
rect 5744 5956 5748 6012
rect 5748 5956 5804 6012
rect 5804 5956 5808 6012
rect 5744 5952 5808 5956
rect 5824 6012 5888 6016
rect 5824 5956 5828 6012
rect 5828 5956 5884 6012
rect 5884 5956 5888 6012
rect 5824 5952 5888 5956
rect 14848 6012 14912 6016
rect 14848 5956 14852 6012
rect 14852 5956 14908 6012
rect 14908 5956 14912 6012
rect 14848 5952 14912 5956
rect 14928 6012 14992 6016
rect 14928 5956 14932 6012
rect 14932 5956 14988 6012
rect 14988 5956 14992 6012
rect 14928 5952 14992 5956
rect 15008 6012 15072 6016
rect 15008 5956 15012 6012
rect 15012 5956 15068 6012
rect 15068 5956 15072 6012
rect 15008 5952 15072 5956
rect 15088 6012 15152 6016
rect 15088 5956 15092 6012
rect 15092 5956 15148 6012
rect 15148 5956 15152 6012
rect 15088 5952 15152 5956
rect 24112 6012 24176 6016
rect 24112 5956 24116 6012
rect 24116 5956 24172 6012
rect 24172 5956 24176 6012
rect 24112 5952 24176 5956
rect 24192 6012 24256 6016
rect 24192 5956 24196 6012
rect 24196 5956 24252 6012
rect 24252 5956 24256 6012
rect 24192 5952 24256 5956
rect 24272 6012 24336 6016
rect 24272 5956 24276 6012
rect 24276 5956 24332 6012
rect 24332 5956 24336 6012
rect 24272 5952 24336 5956
rect 24352 6012 24416 6016
rect 24352 5956 24356 6012
rect 24356 5956 24412 6012
rect 24412 5956 24416 6012
rect 24352 5952 24416 5956
rect 10216 5468 10280 5472
rect 10216 5412 10220 5468
rect 10220 5412 10276 5468
rect 10276 5412 10280 5468
rect 10216 5408 10280 5412
rect 10296 5468 10360 5472
rect 10296 5412 10300 5468
rect 10300 5412 10356 5468
rect 10356 5412 10360 5468
rect 10296 5408 10360 5412
rect 10376 5468 10440 5472
rect 10376 5412 10380 5468
rect 10380 5412 10436 5468
rect 10436 5412 10440 5468
rect 10376 5408 10440 5412
rect 10456 5468 10520 5472
rect 10456 5412 10460 5468
rect 10460 5412 10516 5468
rect 10516 5412 10520 5468
rect 10456 5408 10520 5412
rect 19480 5468 19544 5472
rect 19480 5412 19484 5468
rect 19484 5412 19540 5468
rect 19540 5412 19544 5468
rect 19480 5408 19544 5412
rect 19560 5468 19624 5472
rect 19560 5412 19564 5468
rect 19564 5412 19620 5468
rect 19620 5412 19624 5468
rect 19560 5408 19624 5412
rect 19640 5468 19704 5472
rect 19640 5412 19644 5468
rect 19644 5412 19700 5468
rect 19700 5412 19704 5468
rect 19640 5408 19704 5412
rect 19720 5468 19784 5472
rect 19720 5412 19724 5468
rect 19724 5412 19780 5468
rect 19780 5412 19784 5468
rect 19720 5408 19784 5412
rect 5584 4924 5648 4928
rect 5584 4868 5588 4924
rect 5588 4868 5644 4924
rect 5644 4868 5648 4924
rect 5584 4864 5648 4868
rect 5664 4924 5728 4928
rect 5664 4868 5668 4924
rect 5668 4868 5724 4924
rect 5724 4868 5728 4924
rect 5664 4864 5728 4868
rect 5744 4924 5808 4928
rect 5744 4868 5748 4924
rect 5748 4868 5804 4924
rect 5804 4868 5808 4924
rect 5744 4864 5808 4868
rect 5824 4924 5888 4928
rect 5824 4868 5828 4924
rect 5828 4868 5884 4924
rect 5884 4868 5888 4924
rect 5824 4864 5888 4868
rect 14848 4924 14912 4928
rect 14848 4868 14852 4924
rect 14852 4868 14908 4924
rect 14908 4868 14912 4924
rect 14848 4864 14912 4868
rect 14928 4924 14992 4928
rect 14928 4868 14932 4924
rect 14932 4868 14988 4924
rect 14988 4868 14992 4924
rect 14928 4864 14992 4868
rect 15008 4924 15072 4928
rect 15008 4868 15012 4924
rect 15012 4868 15068 4924
rect 15068 4868 15072 4924
rect 15008 4864 15072 4868
rect 15088 4924 15152 4928
rect 15088 4868 15092 4924
rect 15092 4868 15148 4924
rect 15148 4868 15152 4924
rect 15088 4864 15152 4868
rect 24112 4924 24176 4928
rect 24112 4868 24116 4924
rect 24116 4868 24172 4924
rect 24172 4868 24176 4924
rect 24112 4864 24176 4868
rect 24192 4924 24256 4928
rect 24192 4868 24196 4924
rect 24196 4868 24252 4924
rect 24252 4868 24256 4924
rect 24192 4864 24256 4868
rect 24272 4924 24336 4928
rect 24272 4868 24276 4924
rect 24276 4868 24332 4924
rect 24332 4868 24336 4924
rect 24272 4864 24336 4868
rect 24352 4924 24416 4928
rect 24352 4868 24356 4924
rect 24356 4868 24412 4924
rect 24412 4868 24416 4924
rect 24352 4864 24416 4868
rect 10216 4380 10280 4384
rect 10216 4324 10220 4380
rect 10220 4324 10276 4380
rect 10276 4324 10280 4380
rect 10216 4320 10280 4324
rect 10296 4380 10360 4384
rect 10296 4324 10300 4380
rect 10300 4324 10356 4380
rect 10356 4324 10360 4380
rect 10296 4320 10360 4324
rect 10376 4380 10440 4384
rect 10376 4324 10380 4380
rect 10380 4324 10436 4380
rect 10436 4324 10440 4380
rect 10376 4320 10440 4324
rect 10456 4380 10520 4384
rect 10456 4324 10460 4380
rect 10460 4324 10516 4380
rect 10516 4324 10520 4380
rect 10456 4320 10520 4324
rect 19480 4380 19544 4384
rect 19480 4324 19484 4380
rect 19484 4324 19540 4380
rect 19540 4324 19544 4380
rect 19480 4320 19544 4324
rect 19560 4380 19624 4384
rect 19560 4324 19564 4380
rect 19564 4324 19620 4380
rect 19620 4324 19624 4380
rect 19560 4320 19624 4324
rect 19640 4380 19704 4384
rect 19640 4324 19644 4380
rect 19644 4324 19700 4380
rect 19700 4324 19704 4380
rect 19640 4320 19704 4324
rect 19720 4380 19784 4384
rect 19720 4324 19724 4380
rect 19724 4324 19780 4380
rect 19780 4324 19784 4380
rect 19720 4320 19784 4324
rect 27292 3980 27356 4044
rect 5584 3836 5648 3840
rect 5584 3780 5588 3836
rect 5588 3780 5644 3836
rect 5644 3780 5648 3836
rect 5584 3776 5648 3780
rect 5664 3836 5728 3840
rect 5664 3780 5668 3836
rect 5668 3780 5724 3836
rect 5724 3780 5728 3836
rect 5664 3776 5728 3780
rect 5744 3836 5808 3840
rect 5744 3780 5748 3836
rect 5748 3780 5804 3836
rect 5804 3780 5808 3836
rect 5744 3776 5808 3780
rect 5824 3836 5888 3840
rect 5824 3780 5828 3836
rect 5828 3780 5884 3836
rect 5884 3780 5888 3836
rect 5824 3776 5888 3780
rect 14848 3836 14912 3840
rect 14848 3780 14852 3836
rect 14852 3780 14908 3836
rect 14908 3780 14912 3836
rect 14848 3776 14912 3780
rect 14928 3836 14992 3840
rect 14928 3780 14932 3836
rect 14932 3780 14988 3836
rect 14988 3780 14992 3836
rect 14928 3776 14992 3780
rect 15008 3836 15072 3840
rect 15008 3780 15012 3836
rect 15012 3780 15068 3836
rect 15068 3780 15072 3836
rect 15008 3776 15072 3780
rect 15088 3836 15152 3840
rect 15088 3780 15092 3836
rect 15092 3780 15148 3836
rect 15148 3780 15152 3836
rect 15088 3776 15152 3780
rect 24112 3836 24176 3840
rect 24112 3780 24116 3836
rect 24116 3780 24172 3836
rect 24172 3780 24176 3836
rect 24112 3776 24176 3780
rect 24192 3836 24256 3840
rect 24192 3780 24196 3836
rect 24196 3780 24252 3836
rect 24252 3780 24256 3836
rect 24192 3776 24256 3780
rect 24272 3836 24336 3840
rect 24272 3780 24276 3836
rect 24276 3780 24332 3836
rect 24332 3780 24336 3836
rect 24272 3776 24336 3780
rect 24352 3836 24416 3840
rect 24352 3780 24356 3836
rect 24356 3780 24412 3836
rect 24412 3780 24416 3836
rect 24352 3776 24416 3780
rect 10216 3292 10280 3296
rect 10216 3236 10220 3292
rect 10220 3236 10276 3292
rect 10276 3236 10280 3292
rect 10216 3232 10280 3236
rect 10296 3292 10360 3296
rect 10296 3236 10300 3292
rect 10300 3236 10356 3292
rect 10356 3236 10360 3292
rect 10296 3232 10360 3236
rect 10376 3292 10440 3296
rect 10376 3236 10380 3292
rect 10380 3236 10436 3292
rect 10436 3236 10440 3292
rect 10376 3232 10440 3236
rect 10456 3292 10520 3296
rect 10456 3236 10460 3292
rect 10460 3236 10516 3292
rect 10516 3236 10520 3292
rect 10456 3232 10520 3236
rect 19480 3292 19544 3296
rect 19480 3236 19484 3292
rect 19484 3236 19540 3292
rect 19540 3236 19544 3292
rect 19480 3232 19544 3236
rect 19560 3292 19624 3296
rect 19560 3236 19564 3292
rect 19564 3236 19620 3292
rect 19620 3236 19624 3292
rect 19560 3232 19624 3236
rect 19640 3292 19704 3296
rect 19640 3236 19644 3292
rect 19644 3236 19700 3292
rect 19700 3236 19704 3292
rect 19640 3232 19704 3236
rect 19720 3292 19784 3296
rect 19720 3236 19724 3292
rect 19724 3236 19780 3292
rect 19780 3236 19784 3292
rect 19720 3232 19784 3236
rect 5584 2748 5648 2752
rect 5584 2692 5588 2748
rect 5588 2692 5644 2748
rect 5644 2692 5648 2748
rect 5584 2688 5648 2692
rect 5664 2748 5728 2752
rect 5664 2692 5668 2748
rect 5668 2692 5724 2748
rect 5724 2692 5728 2748
rect 5664 2688 5728 2692
rect 5744 2748 5808 2752
rect 5744 2692 5748 2748
rect 5748 2692 5804 2748
rect 5804 2692 5808 2748
rect 5744 2688 5808 2692
rect 5824 2748 5888 2752
rect 5824 2692 5828 2748
rect 5828 2692 5884 2748
rect 5884 2692 5888 2748
rect 5824 2688 5888 2692
rect 14848 2748 14912 2752
rect 14848 2692 14852 2748
rect 14852 2692 14908 2748
rect 14908 2692 14912 2748
rect 14848 2688 14912 2692
rect 14928 2748 14992 2752
rect 14928 2692 14932 2748
rect 14932 2692 14988 2748
rect 14988 2692 14992 2748
rect 14928 2688 14992 2692
rect 15008 2748 15072 2752
rect 15008 2692 15012 2748
rect 15012 2692 15068 2748
rect 15068 2692 15072 2748
rect 15008 2688 15072 2692
rect 15088 2748 15152 2752
rect 15088 2692 15092 2748
rect 15092 2692 15148 2748
rect 15148 2692 15152 2748
rect 15088 2688 15152 2692
rect 24112 2748 24176 2752
rect 24112 2692 24116 2748
rect 24116 2692 24172 2748
rect 24172 2692 24176 2748
rect 24112 2688 24176 2692
rect 24192 2748 24256 2752
rect 24192 2692 24196 2748
rect 24196 2692 24252 2748
rect 24252 2692 24256 2748
rect 24192 2688 24256 2692
rect 24272 2748 24336 2752
rect 24272 2692 24276 2748
rect 24276 2692 24332 2748
rect 24332 2692 24336 2748
rect 24272 2688 24336 2692
rect 24352 2748 24416 2752
rect 24352 2692 24356 2748
rect 24356 2692 24412 2748
rect 24412 2692 24416 2748
rect 24352 2688 24416 2692
rect 10216 2204 10280 2208
rect 10216 2148 10220 2204
rect 10220 2148 10276 2204
rect 10276 2148 10280 2204
rect 10216 2144 10280 2148
rect 10296 2204 10360 2208
rect 10296 2148 10300 2204
rect 10300 2148 10356 2204
rect 10356 2148 10360 2204
rect 10296 2144 10360 2148
rect 10376 2204 10440 2208
rect 10376 2148 10380 2204
rect 10380 2148 10436 2204
rect 10436 2148 10440 2204
rect 10376 2144 10440 2148
rect 10456 2204 10520 2208
rect 10456 2148 10460 2204
rect 10460 2148 10516 2204
rect 10516 2148 10520 2204
rect 10456 2144 10520 2148
rect 19480 2204 19544 2208
rect 19480 2148 19484 2204
rect 19484 2148 19540 2204
rect 19540 2148 19544 2204
rect 19480 2144 19544 2148
rect 19560 2204 19624 2208
rect 19560 2148 19564 2204
rect 19564 2148 19620 2204
rect 19620 2148 19624 2204
rect 19560 2144 19624 2148
rect 19640 2204 19704 2208
rect 19640 2148 19644 2204
rect 19644 2148 19700 2204
rect 19700 2148 19704 2204
rect 19640 2144 19704 2148
rect 19720 2204 19784 2208
rect 19720 2148 19724 2204
rect 19724 2148 19780 2204
rect 19780 2148 19784 2204
rect 19720 2144 19784 2148
<< metal4 >>
rect 5576 47360 5896 47376
rect 5576 47296 5584 47360
rect 5648 47296 5664 47360
rect 5728 47296 5744 47360
rect 5808 47296 5824 47360
rect 5888 47296 5896 47360
rect 5576 46272 5896 47296
rect 5576 46208 5584 46272
rect 5648 46208 5664 46272
rect 5728 46208 5744 46272
rect 5808 46208 5824 46272
rect 5888 46208 5896 46272
rect 5576 45184 5896 46208
rect 5576 45120 5584 45184
rect 5648 45120 5664 45184
rect 5728 45120 5744 45184
rect 5808 45120 5824 45184
rect 5888 45120 5896 45184
rect 5576 44096 5896 45120
rect 5576 44032 5584 44096
rect 5648 44032 5664 44096
rect 5728 44032 5744 44096
rect 5808 44032 5824 44096
rect 5888 44032 5896 44096
rect 5576 43008 5896 44032
rect 5576 42944 5584 43008
rect 5648 42944 5664 43008
rect 5728 42944 5744 43008
rect 5808 42944 5824 43008
rect 5888 42944 5896 43008
rect 5576 41920 5896 42944
rect 5576 41856 5584 41920
rect 5648 41856 5664 41920
rect 5728 41856 5744 41920
rect 5808 41856 5824 41920
rect 5888 41856 5896 41920
rect 5576 40832 5896 41856
rect 5576 40768 5584 40832
rect 5648 40768 5664 40832
rect 5728 40768 5744 40832
rect 5808 40768 5824 40832
rect 5888 40768 5896 40832
rect 5576 39744 5896 40768
rect 5576 39680 5584 39744
rect 5648 39680 5664 39744
rect 5728 39680 5744 39744
rect 5808 39680 5824 39744
rect 5888 39680 5896 39744
rect 5576 38656 5896 39680
rect 5576 38592 5584 38656
rect 5648 38592 5664 38656
rect 5728 38592 5744 38656
rect 5808 38592 5824 38656
rect 5888 38592 5896 38656
rect 5576 37568 5896 38592
rect 5576 37504 5584 37568
rect 5648 37504 5664 37568
rect 5728 37504 5744 37568
rect 5808 37504 5824 37568
rect 5888 37504 5896 37568
rect 5576 36480 5896 37504
rect 5576 36416 5584 36480
rect 5648 36416 5664 36480
rect 5728 36416 5744 36480
rect 5808 36416 5824 36480
rect 5888 36416 5896 36480
rect 5576 35392 5896 36416
rect 5576 35328 5584 35392
rect 5648 35328 5664 35392
rect 5728 35328 5744 35392
rect 5808 35328 5824 35392
rect 5888 35328 5896 35392
rect 5576 34304 5896 35328
rect 5576 34240 5584 34304
rect 5648 34240 5664 34304
rect 5728 34240 5744 34304
rect 5808 34240 5824 34304
rect 5888 34240 5896 34304
rect 5576 33216 5896 34240
rect 5576 33152 5584 33216
rect 5648 33152 5664 33216
rect 5728 33152 5744 33216
rect 5808 33152 5824 33216
rect 5888 33152 5896 33216
rect 5576 32128 5896 33152
rect 5576 32064 5584 32128
rect 5648 32064 5664 32128
rect 5728 32064 5744 32128
rect 5808 32064 5824 32128
rect 5888 32064 5896 32128
rect 5576 31040 5896 32064
rect 5576 30976 5584 31040
rect 5648 30976 5664 31040
rect 5728 30976 5744 31040
rect 5808 30976 5824 31040
rect 5888 30976 5896 31040
rect 5576 29952 5896 30976
rect 5576 29888 5584 29952
rect 5648 29888 5664 29952
rect 5728 29888 5744 29952
rect 5808 29888 5824 29952
rect 5888 29888 5896 29952
rect 5576 28864 5896 29888
rect 5576 28800 5584 28864
rect 5648 28800 5664 28864
rect 5728 28800 5744 28864
rect 5808 28800 5824 28864
rect 5888 28800 5896 28864
rect 5576 27776 5896 28800
rect 5576 27712 5584 27776
rect 5648 27712 5664 27776
rect 5728 27712 5744 27776
rect 5808 27712 5824 27776
rect 5888 27712 5896 27776
rect 5576 26688 5896 27712
rect 5576 26624 5584 26688
rect 5648 26624 5664 26688
rect 5728 26624 5744 26688
rect 5808 26624 5824 26688
rect 5888 26624 5896 26688
rect 5576 25600 5896 26624
rect 5576 25536 5584 25600
rect 5648 25536 5664 25600
rect 5728 25536 5744 25600
rect 5808 25536 5824 25600
rect 5888 25536 5896 25600
rect 5576 24512 5896 25536
rect 5576 24448 5584 24512
rect 5648 24448 5664 24512
rect 5728 24448 5744 24512
rect 5808 24448 5824 24512
rect 5888 24448 5896 24512
rect 5576 23424 5896 24448
rect 5576 23360 5584 23424
rect 5648 23360 5664 23424
rect 5728 23360 5744 23424
rect 5808 23360 5824 23424
rect 5888 23360 5896 23424
rect 5576 22336 5896 23360
rect 5576 22272 5584 22336
rect 5648 22272 5664 22336
rect 5728 22272 5744 22336
rect 5808 22272 5824 22336
rect 5888 22272 5896 22336
rect 5576 21248 5896 22272
rect 5576 21184 5584 21248
rect 5648 21184 5664 21248
rect 5728 21184 5744 21248
rect 5808 21184 5824 21248
rect 5888 21184 5896 21248
rect 5576 20160 5896 21184
rect 5576 20096 5584 20160
rect 5648 20096 5664 20160
rect 5728 20096 5744 20160
rect 5808 20096 5824 20160
rect 5888 20096 5896 20160
rect 5576 19072 5896 20096
rect 5576 19008 5584 19072
rect 5648 19008 5664 19072
rect 5728 19008 5744 19072
rect 5808 19008 5824 19072
rect 5888 19008 5896 19072
rect 5576 17984 5896 19008
rect 5576 17920 5584 17984
rect 5648 17920 5664 17984
rect 5728 17920 5744 17984
rect 5808 17920 5824 17984
rect 5888 17920 5896 17984
rect 5576 16896 5896 17920
rect 5576 16832 5584 16896
rect 5648 16832 5664 16896
rect 5728 16832 5744 16896
rect 5808 16832 5824 16896
rect 5888 16832 5896 16896
rect 5576 15808 5896 16832
rect 5576 15744 5584 15808
rect 5648 15744 5664 15808
rect 5728 15744 5744 15808
rect 5808 15744 5824 15808
rect 5888 15744 5896 15808
rect 5576 14720 5896 15744
rect 5576 14656 5584 14720
rect 5648 14656 5664 14720
rect 5728 14656 5744 14720
rect 5808 14656 5824 14720
rect 5888 14656 5896 14720
rect 5576 13632 5896 14656
rect 5576 13568 5584 13632
rect 5648 13568 5664 13632
rect 5728 13568 5744 13632
rect 5808 13568 5824 13632
rect 5888 13568 5896 13632
rect 5576 12544 5896 13568
rect 5576 12480 5584 12544
rect 5648 12480 5664 12544
rect 5728 12480 5744 12544
rect 5808 12480 5824 12544
rect 5888 12480 5896 12544
rect 5576 11456 5896 12480
rect 5576 11392 5584 11456
rect 5648 11392 5664 11456
rect 5728 11392 5744 11456
rect 5808 11392 5824 11456
rect 5888 11392 5896 11456
rect 5576 10368 5896 11392
rect 5576 10304 5584 10368
rect 5648 10304 5664 10368
rect 5728 10304 5744 10368
rect 5808 10304 5824 10368
rect 5888 10304 5896 10368
rect 5576 9280 5896 10304
rect 5576 9216 5584 9280
rect 5648 9216 5664 9280
rect 5728 9216 5744 9280
rect 5808 9216 5824 9280
rect 5888 9216 5896 9280
rect 5576 8192 5896 9216
rect 5576 8128 5584 8192
rect 5648 8128 5664 8192
rect 5728 8128 5744 8192
rect 5808 8128 5824 8192
rect 5888 8128 5896 8192
rect 5576 7104 5896 8128
rect 5576 7040 5584 7104
rect 5648 7040 5664 7104
rect 5728 7040 5744 7104
rect 5808 7040 5824 7104
rect 5888 7040 5896 7104
rect 5576 6016 5896 7040
rect 5576 5952 5584 6016
rect 5648 5952 5664 6016
rect 5728 5952 5744 6016
rect 5808 5952 5824 6016
rect 5888 5952 5896 6016
rect 5576 4928 5896 5952
rect 5576 4864 5584 4928
rect 5648 4864 5664 4928
rect 5728 4864 5744 4928
rect 5808 4864 5824 4928
rect 5888 4864 5896 4928
rect 5576 3840 5896 4864
rect 5576 3776 5584 3840
rect 5648 3776 5664 3840
rect 5728 3776 5744 3840
rect 5808 3776 5824 3840
rect 5888 3776 5896 3840
rect 5576 2752 5896 3776
rect 5576 2688 5584 2752
rect 5648 2688 5664 2752
rect 5728 2688 5744 2752
rect 5808 2688 5824 2752
rect 5888 2688 5896 2752
rect 5576 2128 5896 2688
rect 10208 46816 10528 47376
rect 10208 46752 10216 46816
rect 10280 46752 10296 46816
rect 10360 46752 10376 46816
rect 10440 46752 10456 46816
rect 10520 46752 10528 46816
rect 10208 45728 10528 46752
rect 10208 45664 10216 45728
rect 10280 45664 10296 45728
rect 10360 45664 10376 45728
rect 10440 45664 10456 45728
rect 10520 45664 10528 45728
rect 10208 44640 10528 45664
rect 10208 44576 10216 44640
rect 10280 44576 10296 44640
rect 10360 44576 10376 44640
rect 10440 44576 10456 44640
rect 10520 44576 10528 44640
rect 10208 43552 10528 44576
rect 10208 43488 10216 43552
rect 10280 43488 10296 43552
rect 10360 43488 10376 43552
rect 10440 43488 10456 43552
rect 10520 43488 10528 43552
rect 10208 42464 10528 43488
rect 10208 42400 10216 42464
rect 10280 42400 10296 42464
rect 10360 42400 10376 42464
rect 10440 42400 10456 42464
rect 10520 42400 10528 42464
rect 10208 41376 10528 42400
rect 10208 41312 10216 41376
rect 10280 41312 10296 41376
rect 10360 41312 10376 41376
rect 10440 41312 10456 41376
rect 10520 41312 10528 41376
rect 10208 40288 10528 41312
rect 10208 40224 10216 40288
rect 10280 40224 10296 40288
rect 10360 40224 10376 40288
rect 10440 40224 10456 40288
rect 10520 40224 10528 40288
rect 10208 39200 10528 40224
rect 10208 39136 10216 39200
rect 10280 39136 10296 39200
rect 10360 39136 10376 39200
rect 10440 39136 10456 39200
rect 10520 39136 10528 39200
rect 10208 38112 10528 39136
rect 10208 38048 10216 38112
rect 10280 38048 10296 38112
rect 10360 38048 10376 38112
rect 10440 38048 10456 38112
rect 10520 38048 10528 38112
rect 10208 37024 10528 38048
rect 10208 36960 10216 37024
rect 10280 36960 10296 37024
rect 10360 36960 10376 37024
rect 10440 36960 10456 37024
rect 10520 36960 10528 37024
rect 10208 35936 10528 36960
rect 10208 35872 10216 35936
rect 10280 35872 10296 35936
rect 10360 35872 10376 35936
rect 10440 35872 10456 35936
rect 10520 35872 10528 35936
rect 10208 34848 10528 35872
rect 10208 34784 10216 34848
rect 10280 34784 10296 34848
rect 10360 34784 10376 34848
rect 10440 34784 10456 34848
rect 10520 34784 10528 34848
rect 10208 33760 10528 34784
rect 10208 33696 10216 33760
rect 10280 33696 10296 33760
rect 10360 33696 10376 33760
rect 10440 33696 10456 33760
rect 10520 33696 10528 33760
rect 10208 32672 10528 33696
rect 10208 32608 10216 32672
rect 10280 32608 10296 32672
rect 10360 32608 10376 32672
rect 10440 32608 10456 32672
rect 10520 32608 10528 32672
rect 10208 31584 10528 32608
rect 10208 31520 10216 31584
rect 10280 31520 10296 31584
rect 10360 31520 10376 31584
rect 10440 31520 10456 31584
rect 10520 31520 10528 31584
rect 10208 30496 10528 31520
rect 10208 30432 10216 30496
rect 10280 30432 10296 30496
rect 10360 30432 10376 30496
rect 10440 30432 10456 30496
rect 10520 30432 10528 30496
rect 10208 29408 10528 30432
rect 10208 29344 10216 29408
rect 10280 29344 10296 29408
rect 10360 29344 10376 29408
rect 10440 29344 10456 29408
rect 10520 29344 10528 29408
rect 10208 28320 10528 29344
rect 10208 28256 10216 28320
rect 10280 28256 10296 28320
rect 10360 28256 10376 28320
rect 10440 28256 10456 28320
rect 10520 28256 10528 28320
rect 10208 27232 10528 28256
rect 10208 27168 10216 27232
rect 10280 27168 10296 27232
rect 10360 27168 10376 27232
rect 10440 27168 10456 27232
rect 10520 27168 10528 27232
rect 10208 26144 10528 27168
rect 10208 26080 10216 26144
rect 10280 26080 10296 26144
rect 10360 26080 10376 26144
rect 10440 26080 10456 26144
rect 10520 26080 10528 26144
rect 10208 25056 10528 26080
rect 10208 24992 10216 25056
rect 10280 24992 10296 25056
rect 10360 24992 10376 25056
rect 10440 24992 10456 25056
rect 10520 24992 10528 25056
rect 10208 23968 10528 24992
rect 10208 23904 10216 23968
rect 10280 23904 10296 23968
rect 10360 23904 10376 23968
rect 10440 23904 10456 23968
rect 10520 23904 10528 23968
rect 10208 22880 10528 23904
rect 10208 22816 10216 22880
rect 10280 22816 10296 22880
rect 10360 22816 10376 22880
rect 10440 22816 10456 22880
rect 10520 22816 10528 22880
rect 10208 21792 10528 22816
rect 10208 21728 10216 21792
rect 10280 21728 10296 21792
rect 10360 21728 10376 21792
rect 10440 21728 10456 21792
rect 10520 21728 10528 21792
rect 10208 20704 10528 21728
rect 10208 20640 10216 20704
rect 10280 20640 10296 20704
rect 10360 20640 10376 20704
rect 10440 20640 10456 20704
rect 10520 20640 10528 20704
rect 10208 19616 10528 20640
rect 10208 19552 10216 19616
rect 10280 19552 10296 19616
rect 10360 19552 10376 19616
rect 10440 19552 10456 19616
rect 10520 19552 10528 19616
rect 10208 18528 10528 19552
rect 10208 18464 10216 18528
rect 10280 18464 10296 18528
rect 10360 18464 10376 18528
rect 10440 18464 10456 18528
rect 10520 18464 10528 18528
rect 10208 17440 10528 18464
rect 10208 17376 10216 17440
rect 10280 17376 10296 17440
rect 10360 17376 10376 17440
rect 10440 17376 10456 17440
rect 10520 17376 10528 17440
rect 10208 16352 10528 17376
rect 10208 16288 10216 16352
rect 10280 16288 10296 16352
rect 10360 16288 10376 16352
rect 10440 16288 10456 16352
rect 10520 16288 10528 16352
rect 10208 15264 10528 16288
rect 10208 15200 10216 15264
rect 10280 15200 10296 15264
rect 10360 15200 10376 15264
rect 10440 15200 10456 15264
rect 10520 15200 10528 15264
rect 10208 14176 10528 15200
rect 10208 14112 10216 14176
rect 10280 14112 10296 14176
rect 10360 14112 10376 14176
rect 10440 14112 10456 14176
rect 10520 14112 10528 14176
rect 10208 13088 10528 14112
rect 10208 13024 10216 13088
rect 10280 13024 10296 13088
rect 10360 13024 10376 13088
rect 10440 13024 10456 13088
rect 10520 13024 10528 13088
rect 10208 12000 10528 13024
rect 10208 11936 10216 12000
rect 10280 11936 10296 12000
rect 10360 11936 10376 12000
rect 10440 11936 10456 12000
rect 10520 11936 10528 12000
rect 10208 10912 10528 11936
rect 10208 10848 10216 10912
rect 10280 10848 10296 10912
rect 10360 10848 10376 10912
rect 10440 10848 10456 10912
rect 10520 10848 10528 10912
rect 10208 9824 10528 10848
rect 10208 9760 10216 9824
rect 10280 9760 10296 9824
rect 10360 9760 10376 9824
rect 10440 9760 10456 9824
rect 10520 9760 10528 9824
rect 10208 8736 10528 9760
rect 10208 8672 10216 8736
rect 10280 8672 10296 8736
rect 10360 8672 10376 8736
rect 10440 8672 10456 8736
rect 10520 8672 10528 8736
rect 10208 7648 10528 8672
rect 10208 7584 10216 7648
rect 10280 7584 10296 7648
rect 10360 7584 10376 7648
rect 10440 7584 10456 7648
rect 10520 7584 10528 7648
rect 10208 6560 10528 7584
rect 10208 6496 10216 6560
rect 10280 6496 10296 6560
rect 10360 6496 10376 6560
rect 10440 6496 10456 6560
rect 10520 6496 10528 6560
rect 10208 5472 10528 6496
rect 10208 5408 10216 5472
rect 10280 5408 10296 5472
rect 10360 5408 10376 5472
rect 10440 5408 10456 5472
rect 10520 5408 10528 5472
rect 10208 4384 10528 5408
rect 10208 4320 10216 4384
rect 10280 4320 10296 4384
rect 10360 4320 10376 4384
rect 10440 4320 10456 4384
rect 10520 4320 10528 4384
rect 10208 3296 10528 4320
rect 10208 3232 10216 3296
rect 10280 3232 10296 3296
rect 10360 3232 10376 3296
rect 10440 3232 10456 3296
rect 10520 3232 10528 3296
rect 10208 2208 10528 3232
rect 10208 2144 10216 2208
rect 10280 2144 10296 2208
rect 10360 2144 10376 2208
rect 10440 2144 10456 2208
rect 10520 2144 10528 2208
rect 10208 2128 10528 2144
rect 14840 47360 15160 47376
rect 14840 47296 14848 47360
rect 14912 47296 14928 47360
rect 14992 47296 15008 47360
rect 15072 47296 15088 47360
rect 15152 47296 15160 47360
rect 14840 46272 15160 47296
rect 14840 46208 14848 46272
rect 14912 46208 14928 46272
rect 14992 46208 15008 46272
rect 15072 46208 15088 46272
rect 15152 46208 15160 46272
rect 14840 45184 15160 46208
rect 14840 45120 14848 45184
rect 14912 45120 14928 45184
rect 14992 45120 15008 45184
rect 15072 45120 15088 45184
rect 15152 45120 15160 45184
rect 14840 44096 15160 45120
rect 14840 44032 14848 44096
rect 14912 44032 14928 44096
rect 14992 44032 15008 44096
rect 15072 44032 15088 44096
rect 15152 44032 15160 44096
rect 14840 43008 15160 44032
rect 14840 42944 14848 43008
rect 14912 42944 14928 43008
rect 14992 42944 15008 43008
rect 15072 42944 15088 43008
rect 15152 42944 15160 43008
rect 14840 41920 15160 42944
rect 14840 41856 14848 41920
rect 14912 41856 14928 41920
rect 14992 41856 15008 41920
rect 15072 41856 15088 41920
rect 15152 41856 15160 41920
rect 14840 40832 15160 41856
rect 14840 40768 14848 40832
rect 14912 40768 14928 40832
rect 14992 40768 15008 40832
rect 15072 40768 15088 40832
rect 15152 40768 15160 40832
rect 14840 39744 15160 40768
rect 14840 39680 14848 39744
rect 14912 39680 14928 39744
rect 14992 39680 15008 39744
rect 15072 39680 15088 39744
rect 15152 39680 15160 39744
rect 14840 38656 15160 39680
rect 14840 38592 14848 38656
rect 14912 38592 14928 38656
rect 14992 38592 15008 38656
rect 15072 38592 15088 38656
rect 15152 38592 15160 38656
rect 14840 37568 15160 38592
rect 14840 37504 14848 37568
rect 14912 37504 14928 37568
rect 14992 37504 15008 37568
rect 15072 37504 15088 37568
rect 15152 37504 15160 37568
rect 14840 36480 15160 37504
rect 14840 36416 14848 36480
rect 14912 36416 14928 36480
rect 14992 36416 15008 36480
rect 15072 36416 15088 36480
rect 15152 36416 15160 36480
rect 14840 35392 15160 36416
rect 14840 35328 14848 35392
rect 14912 35328 14928 35392
rect 14992 35328 15008 35392
rect 15072 35328 15088 35392
rect 15152 35328 15160 35392
rect 14840 34304 15160 35328
rect 19472 46816 19792 47376
rect 19472 46752 19480 46816
rect 19544 46752 19560 46816
rect 19624 46752 19640 46816
rect 19704 46752 19720 46816
rect 19784 46752 19792 46816
rect 19472 45728 19792 46752
rect 19472 45664 19480 45728
rect 19544 45664 19560 45728
rect 19624 45664 19640 45728
rect 19704 45664 19720 45728
rect 19784 45664 19792 45728
rect 19472 44640 19792 45664
rect 19472 44576 19480 44640
rect 19544 44576 19560 44640
rect 19624 44576 19640 44640
rect 19704 44576 19720 44640
rect 19784 44576 19792 44640
rect 19472 43552 19792 44576
rect 24104 47360 24424 47376
rect 24104 47296 24112 47360
rect 24176 47296 24192 47360
rect 24256 47296 24272 47360
rect 24336 47296 24352 47360
rect 24416 47296 24424 47360
rect 24104 46272 24424 47296
rect 24104 46208 24112 46272
rect 24176 46208 24192 46272
rect 24256 46208 24272 46272
rect 24336 46208 24352 46272
rect 24416 46208 24424 46272
rect 24104 45184 24424 46208
rect 24104 45120 24112 45184
rect 24176 45120 24192 45184
rect 24256 45120 24272 45184
rect 24336 45120 24352 45184
rect 24416 45120 24424 45184
rect 21955 44300 22021 44301
rect 21955 44236 21956 44300
rect 22020 44236 22021 44300
rect 21955 44235 22021 44236
rect 19472 43488 19480 43552
rect 19544 43488 19560 43552
rect 19624 43488 19640 43552
rect 19704 43488 19720 43552
rect 19784 43488 19792 43552
rect 19472 42464 19792 43488
rect 19472 42400 19480 42464
rect 19544 42400 19560 42464
rect 19624 42400 19640 42464
rect 19704 42400 19720 42464
rect 19784 42400 19792 42464
rect 19472 41376 19792 42400
rect 19472 41312 19480 41376
rect 19544 41312 19560 41376
rect 19624 41312 19640 41376
rect 19704 41312 19720 41376
rect 19784 41312 19792 41376
rect 19472 40288 19792 41312
rect 19472 40224 19480 40288
rect 19544 40224 19560 40288
rect 19624 40224 19640 40288
rect 19704 40224 19720 40288
rect 19784 40224 19792 40288
rect 19472 39200 19792 40224
rect 19472 39136 19480 39200
rect 19544 39136 19560 39200
rect 19624 39136 19640 39200
rect 19704 39136 19720 39200
rect 19784 39136 19792 39200
rect 19472 38112 19792 39136
rect 19472 38048 19480 38112
rect 19544 38048 19560 38112
rect 19624 38048 19640 38112
rect 19704 38048 19720 38112
rect 19784 38048 19792 38112
rect 19472 37024 19792 38048
rect 19472 36960 19480 37024
rect 19544 36960 19560 37024
rect 19624 36960 19640 37024
rect 19704 36960 19720 37024
rect 19784 36960 19792 37024
rect 19472 35936 19792 36960
rect 19472 35872 19480 35936
rect 19544 35872 19560 35936
rect 19624 35872 19640 35936
rect 19704 35872 19720 35936
rect 19784 35872 19792 35936
rect 18643 35188 18709 35189
rect 18643 35124 18644 35188
rect 18708 35124 18709 35188
rect 18643 35123 18709 35124
rect 14840 34240 14848 34304
rect 14912 34240 14928 34304
rect 14992 34240 15008 34304
rect 15072 34240 15088 34304
rect 15152 34240 15160 34304
rect 14840 33216 15160 34240
rect 14840 33152 14848 33216
rect 14912 33152 14928 33216
rect 14992 33152 15008 33216
rect 15072 33152 15088 33216
rect 15152 33152 15160 33216
rect 14840 32128 15160 33152
rect 14840 32064 14848 32128
rect 14912 32064 14928 32128
rect 14992 32064 15008 32128
rect 15072 32064 15088 32128
rect 15152 32064 15160 32128
rect 14840 31040 15160 32064
rect 14840 30976 14848 31040
rect 14912 30976 14928 31040
rect 14992 30976 15008 31040
rect 15072 30976 15088 31040
rect 15152 30976 15160 31040
rect 14840 29952 15160 30976
rect 14840 29888 14848 29952
rect 14912 29888 14928 29952
rect 14992 29888 15008 29952
rect 15072 29888 15088 29952
rect 15152 29888 15160 29952
rect 14840 28864 15160 29888
rect 14840 28800 14848 28864
rect 14912 28800 14928 28864
rect 14992 28800 15008 28864
rect 15072 28800 15088 28864
rect 15152 28800 15160 28864
rect 14840 27776 15160 28800
rect 14840 27712 14848 27776
rect 14912 27712 14928 27776
rect 14992 27712 15008 27776
rect 15072 27712 15088 27776
rect 15152 27712 15160 27776
rect 14840 26688 15160 27712
rect 14840 26624 14848 26688
rect 14912 26624 14928 26688
rect 14992 26624 15008 26688
rect 15072 26624 15088 26688
rect 15152 26624 15160 26688
rect 14840 25600 15160 26624
rect 14840 25536 14848 25600
rect 14912 25536 14928 25600
rect 14992 25536 15008 25600
rect 15072 25536 15088 25600
rect 15152 25536 15160 25600
rect 14840 24512 15160 25536
rect 14840 24448 14848 24512
rect 14912 24448 14928 24512
rect 14992 24448 15008 24512
rect 15072 24448 15088 24512
rect 15152 24448 15160 24512
rect 14840 23424 15160 24448
rect 14840 23360 14848 23424
rect 14912 23360 14928 23424
rect 14992 23360 15008 23424
rect 15072 23360 15088 23424
rect 15152 23360 15160 23424
rect 14840 22336 15160 23360
rect 14840 22272 14848 22336
rect 14912 22272 14928 22336
rect 14992 22272 15008 22336
rect 15072 22272 15088 22336
rect 15152 22272 15160 22336
rect 14840 21248 15160 22272
rect 14840 21184 14848 21248
rect 14912 21184 14928 21248
rect 14992 21184 15008 21248
rect 15072 21184 15088 21248
rect 15152 21184 15160 21248
rect 14840 20160 15160 21184
rect 14840 20096 14848 20160
rect 14912 20096 14928 20160
rect 14992 20096 15008 20160
rect 15072 20096 15088 20160
rect 15152 20096 15160 20160
rect 14840 19072 15160 20096
rect 14840 19008 14848 19072
rect 14912 19008 14928 19072
rect 14992 19008 15008 19072
rect 15072 19008 15088 19072
rect 15152 19008 15160 19072
rect 14840 17984 15160 19008
rect 14840 17920 14848 17984
rect 14912 17920 14928 17984
rect 14992 17920 15008 17984
rect 15072 17920 15088 17984
rect 15152 17920 15160 17984
rect 14840 16896 15160 17920
rect 14840 16832 14848 16896
rect 14912 16832 14928 16896
rect 14992 16832 15008 16896
rect 15072 16832 15088 16896
rect 15152 16832 15160 16896
rect 14840 15808 15160 16832
rect 14840 15744 14848 15808
rect 14912 15744 14928 15808
rect 14992 15744 15008 15808
rect 15072 15744 15088 15808
rect 15152 15744 15160 15808
rect 14840 14720 15160 15744
rect 14840 14656 14848 14720
rect 14912 14656 14928 14720
rect 14992 14656 15008 14720
rect 15072 14656 15088 14720
rect 15152 14656 15160 14720
rect 14840 13632 15160 14656
rect 14840 13568 14848 13632
rect 14912 13568 14928 13632
rect 14992 13568 15008 13632
rect 15072 13568 15088 13632
rect 15152 13568 15160 13632
rect 14840 12544 15160 13568
rect 14840 12480 14848 12544
rect 14912 12480 14928 12544
rect 14992 12480 15008 12544
rect 15072 12480 15088 12544
rect 15152 12480 15160 12544
rect 14840 11456 15160 12480
rect 14840 11392 14848 11456
rect 14912 11392 14928 11456
rect 14992 11392 15008 11456
rect 15072 11392 15088 11456
rect 15152 11392 15160 11456
rect 14840 10368 15160 11392
rect 14840 10304 14848 10368
rect 14912 10304 14928 10368
rect 14992 10304 15008 10368
rect 15072 10304 15088 10368
rect 15152 10304 15160 10368
rect 14840 9280 15160 10304
rect 14840 9216 14848 9280
rect 14912 9216 14928 9280
rect 14992 9216 15008 9280
rect 15072 9216 15088 9280
rect 15152 9216 15160 9280
rect 14840 8192 15160 9216
rect 14840 8128 14848 8192
rect 14912 8128 14928 8192
rect 14992 8128 15008 8192
rect 15072 8128 15088 8192
rect 15152 8128 15160 8192
rect 14840 7104 15160 8128
rect 18646 7989 18706 35123
rect 19472 34848 19792 35872
rect 19472 34784 19480 34848
rect 19544 34784 19560 34848
rect 19624 34784 19640 34848
rect 19704 34784 19720 34848
rect 19784 34784 19792 34848
rect 19472 33760 19792 34784
rect 21771 33964 21837 33965
rect 21771 33900 21772 33964
rect 21836 33900 21837 33964
rect 21771 33899 21837 33900
rect 19472 33696 19480 33760
rect 19544 33696 19560 33760
rect 19624 33696 19640 33760
rect 19704 33696 19720 33760
rect 19784 33696 19792 33760
rect 19472 32672 19792 33696
rect 19472 32608 19480 32672
rect 19544 32608 19560 32672
rect 19624 32608 19640 32672
rect 19704 32608 19720 32672
rect 19784 32608 19792 32672
rect 19472 31584 19792 32608
rect 19472 31520 19480 31584
rect 19544 31520 19560 31584
rect 19624 31520 19640 31584
rect 19704 31520 19720 31584
rect 19784 31520 19792 31584
rect 19472 30496 19792 31520
rect 19472 30432 19480 30496
rect 19544 30432 19560 30496
rect 19624 30432 19640 30496
rect 19704 30432 19720 30496
rect 19784 30432 19792 30496
rect 19472 29408 19792 30432
rect 19472 29344 19480 29408
rect 19544 29344 19560 29408
rect 19624 29344 19640 29408
rect 19704 29344 19720 29408
rect 19784 29344 19792 29408
rect 19472 28320 19792 29344
rect 19472 28256 19480 28320
rect 19544 28256 19560 28320
rect 19624 28256 19640 28320
rect 19704 28256 19720 28320
rect 19784 28256 19792 28320
rect 19472 27232 19792 28256
rect 19472 27168 19480 27232
rect 19544 27168 19560 27232
rect 19624 27168 19640 27232
rect 19704 27168 19720 27232
rect 19784 27168 19792 27232
rect 19472 26144 19792 27168
rect 19472 26080 19480 26144
rect 19544 26080 19560 26144
rect 19624 26080 19640 26144
rect 19704 26080 19720 26144
rect 19784 26080 19792 26144
rect 19472 25056 19792 26080
rect 19472 24992 19480 25056
rect 19544 24992 19560 25056
rect 19624 24992 19640 25056
rect 19704 24992 19720 25056
rect 19784 24992 19792 25056
rect 19472 23968 19792 24992
rect 19472 23904 19480 23968
rect 19544 23904 19560 23968
rect 19624 23904 19640 23968
rect 19704 23904 19720 23968
rect 19784 23904 19792 23968
rect 19472 22880 19792 23904
rect 21774 23493 21834 33899
rect 21958 24173 22018 44235
rect 24104 44096 24424 45120
rect 24104 44032 24112 44096
rect 24176 44032 24192 44096
rect 24256 44032 24272 44096
rect 24336 44032 24352 44096
rect 24416 44032 24424 44096
rect 24104 43008 24424 44032
rect 24104 42944 24112 43008
rect 24176 42944 24192 43008
rect 24256 42944 24272 43008
rect 24336 42944 24352 43008
rect 24416 42944 24424 43008
rect 24104 41920 24424 42944
rect 24104 41856 24112 41920
rect 24176 41856 24192 41920
rect 24256 41856 24272 41920
rect 24336 41856 24352 41920
rect 24416 41856 24424 41920
rect 24104 40832 24424 41856
rect 24104 40768 24112 40832
rect 24176 40768 24192 40832
rect 24256 40768 24272 40832
rect 24336 40768 24352 40832
rect 24416 40768 24424 40832
rect 24104 39744 24424 40768
rect 24104 39680 24112 39744
rect 24176 39680 24192 39744
rect 24256 39680 24272 39744
rect 24336 39680 24352 39744
rect 24416 39680 24424 39744
rect 24104 38656 24424 39680
rect 24104 38592 24112 38656
rect 24176 38592 24192 38656
rect 24256 38592 24272 38656
rect 24336 38592 24352 38656
rect 24416 38592 24424 38656
rect 24104 37568 24424 38592
rect 24104 37504 24112 37568
rect 24176 37504 24192 37568
rect 24256 37504 24272 37568
rect 24336 37504 24352 37568
rect 24416 37504 24424 37568
rect 24104 36480 24424 37504
rect 24104 36416 24112 36480
rect 24176 36416 24192 36480
rect 24256 36416 24272 36480
rect 24336 36416 24352 36480
rect 24416 36416 24424 36480
rect 24104 35392 24424 36416
rect 24104 35328 24112 35392
rect 24176 35328 24192 35392
rect 24256 35328 24272 35392
rect 24336 35328 24352 35392
rect 24416 35328 24424 35392
rect 24104 34304 24424 35328
rect 27475 34644 27541 34645
rect 27475 34580 27476 34644
rect 27540 34580 27541 34644
rect 27475 34579 27541 34580
rect 24104 34240 24112 34304
rect 24176 34240 24192 34304
rect 24256 34240 24272 34304
rect 24336 34240 24352 34304
rect 24416 34240 24424 34304
rect 24104 33216 24424 34240
rect 24104 33152 24112 33216
rect 24176 33152 24192 33216
rect 24256 33152 24272 33216
rect 24336 33152 24352 33216
rect 24416 33152 24424 33216
rect 22507 32332 22573 32333
rect 22507 32268 22508 32332
rect 22572 32268 22573 32332
rect 22507 32267 22573 32268
rect 21955 24172 22021 24173
rect 21955 24108 21956 24172
rect 22020 24108 22021 24172
rect 21955 24107 22021 24108
rect 21771 23492 21837 23493
rect 21771 23428 21772 23492
rect 21836 23428 21837 23492
rect 21771 23427 21837 23428
rect 19472 22816 19480 22880
rect 19544 22816 19560 22880
rect 19624 22816 19640 22880
rect 19704 22816 19720 22880
rect 19784 22816 19792 22880
rect 19472 21792 19792 22816
rect 19472 21728 19480 21792
rect 19544 21728 19560 21792
rect 19624 21728 19640 21792
rect 19704 21728 19720 21792
rect 19784 21728 19792 21792
rect 19472 20704 19792 21728
rect 22510 21589 22570 32267
rect 24104 32128 24424 33152
rect 24104 32064 24112 32128
rect 24176 32064 24192 32128
rect 24256 32064 24272 32128
rect 24336 32064 24352 32128
rect 24416 32064 24424 32128
rect 24104 31040 24424 32064
rect 24104 30976 24112 31040
rect 24176 30976 24192 31040
rect 24256 30976 24272 31040
rect 24336 30976 24352 31040
rect 24416 30976 24424 31040
rect 24104 29952 24424 30976
rect 24104 29888 24112 29952
rect 24176 29888 24192 29952
rect 24256 29888 24272 29952
rect 24336 29888 24352 29952
rect 24416 29888 24424 29952
rect 24104 28864 24424 29888
rect 24104 28800 24112 28864
rect 24176 28800 24192 28864
rect 24256 28800 24272 28864
rect 24336 28800 24352 28864
rect 24416 28800 24424 28864
rect 24104 27776 24424 28800
rect 24104 27712 24112 27776
rect 24176 27712 24192 27776
rect 24256 27712 24272 27776
rect 24336 27712 24352 27776
rect 24416 27712 24424 27776
rect 24104 26688 24424 27712
rect 24104 26624 24112 26688
rect 24176 26624 24192 26688
rect 24256 26624 24272 26688
rect 24336 26624 24352 26688
rect 24416 26624 24424 26688
rect 24104 25600 24424 26624
rect 24104 25536 24112 25600
rect 24176 25536 24192 25600
rect 24256 25536 24272 25600
rect 24336 25536 24352 25600
rect 24416 25536 24424 25600
rect 24104 24512 24424 25536
rect 24104 24448 24112 24512
rect 24176 24448 24192 24512
rect 24256 24448 24272 24512
rect 24336 24448 24352 24512
rect 24416 24448 24424 24512
rect 24104 23424 24424 24448
rect 24104 23360 24112 23424
rect 24176 23360 24192 23424
rect 24256 23360 24272 23424
rect 24336 23360 24352 23424
rect 24416 23360 24424 23424
rect 24104 22336 24424 23360
rect 24104 22272 24112 22336
rect 24176 22272 24192 22336
rect 24256 22272 24272 22336
rect 24336 22272 24352 22336
rect 24416 22272 24424 22336
rect 22507 21588 22573 21589
rect 22507 21524 22508 21588
rect 22572 21524 22573 21588
rect 22507 21523 22573 21524
rect 19472 20640 19480 20704
rect 19544 20640 19560 20704
rect 19624 20640 19640 20704
rect 19704 20640 19720 20704
rect 19784 20640 19792 20704
rect 19472 19616 19792 20640
rect 19472 19552 19480 19616
rect 19544 19552 19560 19616
rect 19624 19552 19640 19616
rect 19704 19552 19720 19616
rect 19784 19552 19792 19616
rect 19472 18528 19792 19552
rect 19472 18464 19480 18528
rect 19544 18464 19560 18528
rect 19624 18464 19640 18528
rect 19704 18464 19720 18528
rect 19784 18464 19792 18528
rect 19472 17440 19792 18464
rect 19472 17376 19480 17440
rect 19544 17376 19560 17440
rect 19624 17376 19640 17440
rect 19704 17376 19720 17440
rect 19784 17376 19792 17440
rect 19472 16352 19792 17376
rect 19472 16288 19480 16352
rect 19544 16288 19560 16352
rect 19624 16288 19640 16352
rect 19704 16288 19720 16352
rect 19784 16288 19792 16352
rect 19472 15264 19792 16288
rect 19472 15200 19480 15264
rect 19544 15200 19560 15264
rect 19624 15200 19640 15264
rect 19704 15200 19720 15264
rect 19784 15200 19792 15264
rect 19472 14176 19792 15200
rect 19472 14112 19480 14176
rect 19544 14112 19560 14176
rect 19624 14112 19640 14176
rect 19704 14112 19720 14176
rect 19784 14112 19792 14176
rect 19472 13088 19792 14112
rect 19472 13024 19480 13088
rect 19544 13024 19560 13088
rect 19624 13024 19640 13088
rect 19704 13024 19720 13088
rect 19784 13024 19792 13088
rect 19472 12000 19792 13024
rect 19472 11936 19480 12000
rect 19544 11936 19560 12000
rect 19624 11936 19640 12000
rect 19704 11936 19720 12000
rect 19784 11936 19792 12000
rect 19472 10912 19792 11936
rect 19472 10848 19480 10912
rect 19544 10848 19560 10912
rect 19624 10848 19640 10912
rect 19704 10848 19720 10912
rect 19784 10848 19792 10912
rect 19472 9824 19792 10848
rect 19472 9760 19480 9824
rect 19544 9760 19560 9824
rect 19624 9760 19640 9824
rect 19704 9760 19720 9824
rect 19784 9760 19792 9824
rect 19472 8736 19792 9760
rect 19472 8672 19480 8736
rect 19544 8672 19560 8736
rect 19624 8672 19640 8736
rect 19704 8672 19720 8736
rect 19784 8672 19792 8736
rect 18643 7988 18709 7989
rect 18643 7924 18644 7988
rect 18708 7924 18709 7988
rect 18643 7923 18709 7924
rect 14840 7040 14848 7104
rect 14912 7040 14928 7104
rect 14992 7040 15008 7104
rect 15072 7040 15088 7104
rect 15152 7040 15160 7104
rect 14840 6016 15160 7040
rect 14840 5952 14848 6016
rect 14912 5952 14928 6016
rect 14992 5952 15008 6016
rect 15072 5952 15088 6016
rect 15152 5952 15160 6016
rect 14840 4928 15160 5952
rect 14840 4864 14848 4928
rect 14912 4864 14928 4928
rect 14992 4864 15008 4928
rect 15072 4864 15088 4928
rect 15152 4864 15160 4928
rect 14840 3840 15160 4864
rect 14840 3776 14848 3840
rect 14912 3776 14928 3840
rect 14992 3776 15008 3840
rect 15072 3776 15088 3840
rect 15152 3776 15160 3840
rect 14840 2752 15160 3776
rect 14840 2688 14848 2752
rect 14912 2688 14928 2752
rect 14992 2688 15008 2752
rect 15072 2688 15088 2752
rect 15152 2688 15160 2752
rect 14840 2128 15160 2688
rect 19472 7648 19792 8672
rect 19472 7584 19480 7648
rect 19544 7584 19560 7648
rect 19624 7584 19640 7648
rect 19704 7584 19720 7648
rect 19784 7584 19792 7648
rect 19472 6560 19792 7584
rect 19472 6496 19480 6560
rect 19544 6496 19560 6560
rect 19624 6496 19640 6560
rect 19704 6496 19720 6560
rect 19784 6496 19792 6560
rect 19472 5472 19792 6496
rect 19472 5408 19480 5472
rect 19544 5408 19560 5472
rect 19624 5408 19640 5472
rect 19704 5408 19720 5472
rect 19784 5408 19792 5472
rect 19472 4384 19792 5408
rect 19472 4320 19480 4384
rect 19544 4320 19560 4384
rect 19624 4320 19640 4384
rect 19704 4320 19720 4384
rect 19784 4320 19792 4384
rect 19472 3296 19792 4320
rect 19472 3232 19480 3296
rect 19544 3232 19560 3296
rect 19624 3232 19640 3296
rect 19704 3232 19720 3296
rect 19784 3232 19792 3296
rect 19472 2208 19792 3232
rect 19472 2144 19480 2208
rect 19544 2144 19560 2208
rect 19624 2144 19640 2208
rect 19704 2144 19720 2208
rect 19784 2144 19792 2208
rect 19472 2128 19792 2144
rect 24104 21248 24424 22272
rect 24104 21184 24112 21248
rect 24176 21184 24192 21248
rect 24256 21184 24272 21248
rect 24336 21184 24352 21248
rect 24416 21184 24424 21248
rect 24104 20160 24424 21184
rect 27291 20364 27357 20365
rect 27291 20300 27292 20364
rect 27356 20300 27357 20364
rect 27291 20299 27357 20300
rect 24104 20096 24112 20160
rect 24176 20096 24192 20160
rect 24256 20096 24272 20160
rect 24336 20096 24352 20160
rect 24416 20096 24424 20160
rect 24104 19072 24424 20096
rect 24104 19008 24112 19072
rect 24176 19008 24192 19072
rect 24256 19008 24272 19072
rect 24336 19008 24352 19072
rect 24416 19008 24424 19072
rect 24104 17984 24424 19008
rect 24104 17920 24112 17984
rect 24176 17920 24192 17984
rect 24256 17920 24272 17984
rect 24336 17920 24352 17984
rect 24416 17920 24424 17984
rect 24104 16896 24424 17920
rect 24104 16832 24112 16896
rect 24176 16832 24192 16896
rect 24256 16832 24272 16896
rect 24336 16832 24352 16896
rect 24416 16832 24424 16896
rect 24104 15808 24424 16832
rect 24104 15744 24112 15808
rect 24176 15744 24192 15808
rect 24256 15744 24272 15808
rect 24336 15744 24352 15808
rect 24416 15744 24424 15808
rect 24104 14720 24424 15744
rect 24104 14656 24112 14720
rect 24176 14656 24192 14720
rect 24256 14656 24272 14720
rect 24336 14656 24352 14720
rect 24416 14656 24424 14720
rect 24104 13632 24424 14656
rect 24104 13568 24112 13632
rect 24176 13568 24192 13632
rect 24256 13568 24272 13632
rect 24336 13568 24352 13632
rect 24416 13568 24424 13632
rect 24104 12544 24424 13568
rect 24104 12480 24112 12544
rect 24176 12480 24192 12544
rect 24256 12480 24272 12544
rect 24336 12480 24352 12544
rect 24416 12480 24424 12544
rect 24104 11456 24424 12480
rect 24104 11392 24112 11456
rect 24176 11392 24192 11456
rect 24256 11392 24272 11456
rect 24336 11392 24352 11456
rect 24416 11392 24424 11456
rect 24104 10368 24424 11392
rect 24104 10304 24112 10368
rect 24176 10304 24192 10368
rect 24256 10304 24272 10368
rect 24336 10304 24352 10368
rect 24416 10304 24424 10368
rect 24104 9280 24424 10304
rect 24104 9216 24112 9280
rect 24176 9216 24192 9280
rect 24256 9216 24272 9280
rect 24336 9216 24352 9280
rect 24416 9216 24424 9280
rect 24104 8192 24424 9216
rect 24104 8128 24112 8192
rect 24176 8128 24192 8192
rect 24256 8128 24272 8192
rect 24336 8128 24352 8192
rect 24416 8128 24424 8192
rect 24104 7104 24424 8128
rect 24104 7040 24112 7104
rect 24176 7040 24192 7104
rect 24256 7040 24272 7104
rect 24336 7040 24352 7104
rect 24416 7040 24424 7104
rect 24104 6016 24424 7040
rect 24104 5952 24112 6016
rect 24176 5952 24192 6016
rect 24256 5952 24272 6016
rect 24336 5952 24352 6016
rect 24416 5952 24424 6016
rect 24104 4928 24424 5952
rect 24104 4864 24112 4928
rect 24176 4864 24192 4928
rect 24256 4864 24272 4928
rect 24336 4864 24352 4928
rect 24416 4864 24424 4928
rect 24104 3840 24424 4864
rect 27294 4045 27354 20299
rect 27478 13973 27538 34579
rect 27475 13972 27541 13973
rect 27475 13908 27476 13972
rect 27540 13908 27541 13972
rect 27475 13907 27541 13908
rect 27291 4044 27357 4045
rect 27291 3980 27292 4044
rect 27356 3980 27357 4044
rect 27291 3979 27357 3980
rect 24104 3776 24112 3840
rect 24176 3776 24192 3840
rect 24256 3776 24272 3840
rect 24336 3776 24352 3840
rect 24416 3776 24424 3840
rect 24104 2752 24424 3776
rect 24104 2688 24112 2752
rect 24176 2688 24192 2752
rect 24256 2688 24272 2752
rect 24336 2688 24352 2752
rect 24416 2688 24424 2752
rect 24104 2128 24424 2688
use sky130_fd_sc_hd__decap_12  FILLER_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 2484 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3128 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3772 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 4324 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 5060 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48
timestamp 1644511149
transform 1 0 5520 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_0_60
timestamp 1644511149
transform 1 0 6624 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_72
timestamp 1644511149
transform 1 0 7728 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_85
timestamp 1644511149
transform 1 0 8924 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_93
timestamp 1644511149
transform 1 0 9660 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_105
timestamp 1644511149
transform 1 0 10764 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_111 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 11316 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_113
timestamp 1644511149
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_125
timestamp 1644511149
transform 1 0 12604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_137
timestamp 1644511149
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_141
timestamp 1644511149
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_153
timestamp 1644511149
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_165
timestamp 1644511149
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_173
timestamp 1644511149
transform 1 0 17020 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_177
timestamp 1644511149
transform 1 0 17388 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_181
timestamp 1644511149
transform 1 0 17756 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_193
timestamp 1644511149
transform 1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_197
timestamp 1644511149
transform 1 0 19228 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_0_202
timestamp 1644511149
transform 1 0 19688 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_214
timestamp 1644511149
transform 1 0 20792 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_222
timestamp 1644511149
transform 1 0 21528 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_0_225
timestamp 1644511149
transform 1 0 21804 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_237
timestamp 1644511149
transform 1 0 22908 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_249
timestamp 1644511149
transform 1 0 24012 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_253
timestamp 1644511149
transform 1 0 24380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_276
timestamp 1644511149
transform 1 0 26496 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_281
timestamp 1644511149
transform 1 0 26956 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_293
timestamp 1644511149
transform 1 0 28060 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_1_3
timestamp 1644511149
transform 1 0 1380 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_27
timestamp 1644511149
transform 1 0 3588 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_52
timestamp 1644511149
transform 1 0 5888 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_78
timestamp 1644511149
transform 1 0 8280 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_103
timestamp 1644511149
transform 1 0 10580 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 1644511149
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_134
timestamp 1644511149
transform 1 0 13432 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_142
timestamp 1644511149
transform 1 0 14168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_164
timestamp 1644511149
transform 1 0 16192 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_190
timestamp 1644511149
transform 1 0 18584 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_198
timestamp 1644511149
transform 1 0 19320 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_220
timestamp 1644511149
transform 1 0 21344 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_228
timestamp 1644511149
transform 1 0 22080 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_240
timestamp 1644511149
transform 1 0 23184 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_245
timestamp 1644511149
transform 1 0 23644 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_270
timestamp 1644511149
transform 1 0 25944 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_278
timestamp 1644511149
transform 1 0 26680 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_284
timestamp 1644511149
transform 1 0 27232 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_291
timestamp 1644511149
transform 1 0 27876 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_2_6
timestamp 1644511149
transform 1 0 1656 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_13
timestamp 1644511149
transform 1 0 2300 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_17
timestamp 1644511149
transform 1 0 2668 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_21
timestamp 1644511149
transform 1 0 3036 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1644511149
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_29
timestamp 1644511149
transform 1 0 3772 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_36
timestamp 1644511149
transform 1 0 4416 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_2_65
timestamp 1644511149
transform 1 0 7084 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_72
timestamp 1644511149
transform 1 0 7728 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_76
timestamp 1644511149
transform 1 0 8096 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_80
timestamp 1644511149
transform 1 0 8464 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_85
timestamp 1644511149
transform 1 0 8924 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_108
timestamp 1644511149
transform 1 0 11040 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_115
timestamp 1644511149
transform 1 0 11684 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_2_126
timestamp 1644511149
transform 1 0 12696 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_133
timestamp 1644511149
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 1644511149
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_141
timestamp 1644511149
transform 1 0 14076 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_148
timestamp 1644511149
transform 1 0 14720 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_155
timestamp 1644511149
transform 1 0 15364 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_163
timestamp 1644511149
transform 1 0 16100 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_168
timestamp 1644511149
transform 1 0 16560 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_175
timestamp 1644511149
transform 1 0 17204 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_183
timestamp 1644511149
transform 1 0 17940 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_188
timestamp 1644511149
transform 1 0 18400 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_197
timestamp 1644511149
transform 1 0 19228 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_2_203
timestamp 1644511149
transform 1 0 19780 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_211
timestamp 1644511149
transform 1 0 20516 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_215
timestamp 1644511149
transform 1 0 20884 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_240
timestamp 1644511149
transform 1 0 23184 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_256
timestamp 1644511149
transform 1 0 24656 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_262
timestamp 1644511149
transform 1 0 25208 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_266
timestamp 1644511149
transform 1 0 25576 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_2_295
timestamp 1644511149
transform 1 0 28244 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_3
timestamp 1644511149
transform 1 0 1380 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_8
timestamp 1644511149
transform 1 0 1840 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_15
timestamp 1644511149
transform 1 0 2484 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_40
timestamp 1644511149
transform 1 0 4784 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_44
timestamp 1644511149
transform 1 0 5152 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_48
timestamp 1644511149
transform 1 0 5520 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_3_60
timestamp 1644511149
transform 1 0 6624 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_66
timestamp 1644511149
transform 1 0 7176 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_70
timestamp 1644511149
transform 1 0 7544 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_82
timestamp 1644511149
transform 1 0 8648 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_3_91
timestamp 1644511149
transform 1 0 9476 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_3_99
timestamp 1644511149
transform 1 0 10212 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp 1644511149
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1644511149
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_113
timestamp 1644511149
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_125
timestamp 1644511149
transform 1 0 12604 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_150
timestamp 1644511149
transform 1 0 14904 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_162
timestamp 1644511149
transform 1 0 16008 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_3_169
timestamp 1644511149
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_3_181
timestamp 1644511149
transform 1 0 17756 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_3_205
timestamp 1644511149
transform 1 0 19964 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_213
timestamp 1644511149
transform 1 0 20700 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_217
timestamp 1644511149
transform 1 0 21068 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_223
timestamp 1644511149
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_228
timestamp 1644511149
transform 1 0 22080 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_240
timestamp 1644511149
transform 1 0 23184 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_252
timestamp 1644511149
transform 1 0 24288 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_264
timestamp 1644511149
transform 1 0 25392 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_272
timestamp 1644511149
transform 1 0 26128 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_276
timestamp 1644511149
transform 1 0 26496 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_284
timestamp 1644511149
transform 1 0 27232 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_290
timestamp 1644511149
transform 1 0 27784 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_294
timestamp 1644511149
transform 1 0 28152 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_298
timestamp 1644511149
transform 1 0 28520 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_24
timestamp 1644511149
transform 1 0 3312 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_29
timestamp 1644511149
transform 1 0 3772 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_35
timestamp 1644511149
transform 1 0 4324 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_57
timestamp 1644511149
transform 1 0 6348 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_69
timestamp 1644511149
transform 1 0 7452 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_81
timestamp 1644511149
transform 1 0 8556 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_85
timestamp 1644511149
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_97
timestamp 1644511149
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_109
timestamp 1644511149
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_121
timestamp 1644511149
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp 1644511149
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1644511149
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_141
timestamp 1644511149
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_153
timestamp 1644511149
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_165
timestamp 1644511149
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_177
timestamp 1644511149
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_189
timestamp 1644511149
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 1644511149
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_197
timestamp 1644511149
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_209
timestamp 1644511149
transform 1 0 20332 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_234
timestamp 1644511149
transform 1 0 22632 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_246
timestamp 1644511149
transform 1 0 23736 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_4_253
timestamp 1644511149
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_265
timestamp 1644511149
transform 1 0 25484 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_273
timestamp 1644511149
transform 1 0 26220 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_295
timestamp 1644511149
transform 1 0 28244 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_3
timestamp 1644511149
transform 1 0 1380 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_7
timestamp 1644511149
transform 1 0 1748 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_11
timestamp 1644511149
transform 1 0 2116 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_36
timestamp 1644511149
transform 1 0 4416 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_5_43
timestamp 1644511149
transform 1 0 5060 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1644511149
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_57
timestamp 1644511149
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_69
timestamp 1644511149
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_81
timestamp 1644511149
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_93
timestamp 1644511149
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 1644511149
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1644511149
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_113
timestamp 1644511149
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_125
timestamp 1644511149
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_137
timestamp 1644511149
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_149
timestamp 1644511149
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp 1644511149
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1644511149
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_169
timestamp 1644511149
transform 1 0 16652 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_177
timestamp 1644511149
transform 1 0 17388 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_183
timestamp 1644511149
transform 1 0 17940 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_195
timestamp 1644511149
transform 1 0 19044 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_207
timestamp 1644511149
transform 1 0 20148 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_219
timestamp 1644511149
transform 1 0 21252 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_223
timestamp 1644511149
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_225
timestamp 1644511149
transform 1 0 21804 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_233
timestamp 1644511149
transform 1 0 22540 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_240
timestamp 1644511149
transform 1 0 23184 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_252
timestamp 1644511149
transform 1 0 24288 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_264
timestamp 1644511149
transform 1 0 25392 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_276
timestamp 1644511149
transform 1 0 26496 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_281
timestamp 1644511149
transform 1 0 26956 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_285
timestamp 1644511149
transform 1 0 27324 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_289
timestamp 1644511149
transform 1 0 27692 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_297
timestamp 1644511149
transform 1 0 28428 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_3
timestamp 1644511149
transform 1 0 1380 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_6_14
timestamp 1644511149
transform 1 0 2392 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_21
timestamp 1644511149
transform 1 0 3036 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1644511149
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_29
timestamp 1644511149
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_41
timestamp 1644511149
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_53
timestamp 1644511149
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_65
timestamp 1644511149
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 1644511149
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1644511149
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_85
timestamp 1644511149
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_97
timestamp 1644511149
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_109
timestamp 1644511149
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_121
timestamp 1644511149
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1644511149
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1644511149
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_141
timestamp 1644511149
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_153
timestamp 1644511149
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_165
timestamp 1644511149
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_177
timestamp 1644511149
transform 1 0 17388 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_185
timestamp 1644511149
transform 1 0 18124 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_192
timestamp 1644511149
transform 1 0 18768 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_197
timestamp 1644511149
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_209
timestamp 1644511149
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_221
timestamp 1644511149
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_233
timestamp 1644511149
transform 1 0 22540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_245
timestamp 1644511149
transform 1 0 23644 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp 1644511149
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_253
timestamp 1644511149
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_265
timestamp 1644511149
transform 1 0 25484 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_273
timestamp 1644511149
transform 1 0 26220 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_295
timestamp 1644511149
transform 1 0 28244 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_3
timestamp 1644511149
transform 1 0 1380 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_7
timestamp 1644511149
transform 1 0 1748 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_7_32
timestamp 1644511149
transform 1 0 4048 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_44
timestamp 1644511149
transform 1 0 5152 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_57
timestamp 1644511149
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_69
timestamp 1644511149
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_81
timestamp 1644511149
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_93
timestamp 1644511149
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 1644511149
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1644511149
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_113
timestamp 1644511149
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_125
timestamp 1644511149
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_137
timestamp 1644511149
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_149
timestamp 1644511149
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_161
timestamp 1644511149
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1644511149
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_169
timestamp 1644511149
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_181
timestamp 1644511149
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_193
timestamp 1644511149
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_205
timestamp 1644511149
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_217
timestamp 1644511149
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp 1644511149
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_225
timestamp 1644511149
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_237
timestamp 1644511149
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_249
timestamp 1644511149
transform 1 0 24012 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_261
timestamp 1644511149
transform 1 0 25116 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_273
timestamp 1644511149
transform 1 0 26220 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_279
timestamp 1644511149
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_281
timestamp 1644511149
transform 1 0 26956 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_285
timestamp 1644511149
transform 1 0 27324 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_292
timestamp 1644511149
transform 1 0 27968 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_298
timestamp 1644511149
transform 1 0 28520 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_3
timestamp 1644511149
transform 1 0 1380 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_7
timestamp 1644511149
transform 1 0 1748 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_11
timestamp 1644511149
transform 1 0 2116 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_23
timestamp 1644511149
transform 1 0 3220 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1644511149
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_32
timestamp 1644511149
transform 1 0 4048 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_44
timestamp 1644511149
transform 1 0 5152 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_56
timestamp 1644511149
transform 1 0 6256 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_68
timestamp 1644511149
transform 1 0 7360 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_80
timestamp 1644511149
transform 1 0 8464 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_85
timestamp 1644511149
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_97
timestamp 1644511149
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_109
timestamp 1644511149
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_121
timestamp 1644511149
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_133
timestamp 1644511149
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1644511149
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_141
timestamp 1644511149
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_153
timestamp 1644511149
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_165
timestamp 1644511149
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_177
timestamp 1644511149
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_189
timestamp 1644511149
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1644511149
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_197
timestamp 1644511149
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_209
timestamp 1644511149
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_221
timestamp 1644511149
transform 1 0 21436 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_233
timestamp 1644511149
transform 1 0 22540 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_245
timestamp 1644511149
transform 1 0 23644 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_251
timestamp 1644511149
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_253
timestamp 1644511149
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_265
timestamp 1644511149
transform 1 0 25484 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_273
timestamp 1644511149
transform 1 0 26220 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_295
timestamp 1644511149
transform 1 0 28244 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_3
timestamp 1644511149
transform 1 0 1380 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_25
timestamp 1644511149
transform 1 0 3404 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_50
timestamp 1644511149
transform 1 0 5704 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_9_57
timestamp 1644511149
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_69
timestamp 1644511149
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_81
timestamp 1644511149
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_93
timestamp 1644511149
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_105
timestamp 1644511149
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1644511149
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_113
timestamp 1644511149
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_125
timestamp 1644511149
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_137
timestamp 1644511149
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_149
timestamp 1644511149
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_161
timestamp 1644511149
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1644511149
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_169
timestamp 1644511149
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_181
timestamp 1644511149
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_193
timestamp 1644511149
transform 1 0 18860 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_205
timestamp 1644511149
transform 1 0 19964 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_217
timestamp 1644511149
transform 1 0 21068 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_223
timestamp 1644511149
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_225
timestamp 1644511149
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_237
timestamp 1644511149
transform 1 0 22908 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_249
timestamp 1644511149
transform 1 0 24012 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_9_276
timestamp 1644511149
transform 1 0 26496 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_284
timestamp 1644511149
transform 1 0 27232 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_290
timestamp 1644511149
transform 1 0 27784 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_294
timestamp 1644511149
transform 1 0 28152 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_298
timestamp 1644511149
transform 1 0 28520 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_3
timestamp 1644511149
transform 1 0 1380 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_7
timestamp 1644511149
transform 1 0 1748 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_11
timestamp 1644511149
transform 1 0 2116 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_19
timestamp 1644511149
transform 1 0 2852 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_23
timestamp 1644511149
transform 1 0 3220 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1644511149
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_32
timestamp 1644511149
transform 1 0 4048 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_39
timestamp 1644511149
transform 1 0 4692 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_51
timestamp 1644511149
transform 1 0 5796 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_63
timestamp 1644511149
transform 1 0 6900 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_75
timestamp 1644511149
transform 1 0 8004 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1644511149
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_85
timestamp 1644511149
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_97
timestamp 1644511149
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_109
timestamp 1644511149
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_121
timestamp 1644511149
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_133
timestamp 1644511149
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1644511149
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_141
timestamp 1644511149
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_153
timestamp 1644511149
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_165
timestamp 1644511149
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_177
timestamp 1644511149
transform 1 0 17388 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_189
timestamp 1644511149
transform 1 0 18492 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_195
timestamp 1644511149
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_197
timestamp 1644511149
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_209
timestamp 1644511149
transform 1 0 20332 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_221
timestamp 1644511149
transform 1 0 21436 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_233
timestamp 1644511149
transform 1 0 22540 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_245
timestamp 1644511149
transform 1 0 23644 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_251
timestamp 1644511149
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_253
timestamp 1644511149
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_10_265
timestamp 1644511149
transform 1 0 25484 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_270
timestamp 1644511149
transform 1 0 25944 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_295
timestamp 1644511149
transform 1 0 28244 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_3
timestamp 1644511149
transform 1 0 1380 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_11_8
timestamp 1644511149
transform 1 0 1840 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_41
timestamp 1644511149
transform 1 0 4876 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_11_53
timestamp 1644511149
transform 1 0 5980 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_57
timestamp 1644511149
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_69
timestamp 1644511149
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_81
timestamp 1644511149
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_93
timestamp 1644511149
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_105
timestamp 1644511149
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1644511149
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_113
timestamp 1644511149
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_125
timestamp 1644511149
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_137
timestamp 1644511149
transform 1 0 13708 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_149
timestamp 1644511149
transform 1 0 14812 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_161
timestamp 1644511149
transform 1 0 15916 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp 1644511149
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_169
timestamp 1644511149
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_181
timestamp 1644511149
transform 1 0 17756 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_193
timestamp 1644511149
transform 1 0 18860 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_205
timestamp 1644511149
transform 1 0 19964 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_217
timestamp 1644511149
transform 1 0 21068 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_223
timestamp 1644511149
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_225
timestamp 1644511149
transform 1 0 21804 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_237
timestamp 1644511149
transform 1 0 22908 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_249
timestamp 1644511149
transform 1 0 24012 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_11_276
timestamp 1644511149
transform 1 0 26496 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_281
timestamp 1644511149
transform 1 0 26956 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_286
timestamp 1644511149
transform 1 0 27416 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_293
timestamp 1644511149
transform 1 0 28060 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_12_24
timestamp 1644511149
transform 1 0 3312 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_12_29
timestamp 1644511149
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_41
timestamp 1644511149
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_53
timestamp 1644511149
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_65
timestamp 1644511149
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 1644511149
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1644511149
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_85
timestamp 1644511149
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_97
timestamp 1644511149
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_109
timestamp 1644511149
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_121
timestamp 1644511149
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_133
timestamp 1644511149
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1644511149
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_141
timestamp 1644511149
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_153
timestamp 1644511149
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_165
timestamp 1644511149
transform 1 0 16284 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_177
timestamp 1644511149
transform 1 0 17388 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_189
timestamp 1644511149
transform 1 0 18492 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_195
timestamp 1644511149
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_197
timestamp 1644511149
transform 1 0 19228 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_209
timestamp 1644511149
transform 1 0 20332 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_221
timestamp 1644511149
transform 1 0 21436 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_233
timestamp 1644511149
transform 1 0 22540 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_245
timestamp 1644511149
transform 1 0 23644 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_251
timestamp 1644511149
transform 1 0 24196 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_253
timestamp 1644511149
transform 1 0 24380 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_257
timestamp 1644511149
transform 1 0 24748 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_264
timestamp 1644511149
transform 1 0 25392 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_272
timestamp 1644511149
transform 1 0 26128 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_295
timestamp 1644511149
transform 1 0 28244 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_3
timestamp 1644511149
transform 1 0 1380 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_13_30
timestamp 1644511149
transform 1 0 3864 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_42
timestamp 1644511149
transform 1 0 4968 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_54
timestamp 1644511149
transform 1 0 6072 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_13_57
timestamp 1644511149
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_69
timestamp 1644511149
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_81
timestamp 1644511149
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_93
timestamp 1644511149
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_105
timestamp 1644511149
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1644511149
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_113
timestamp 1644511149
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_125
timestamp 1644511149
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_137
timestamp 1644511149
transform 1 0 13708 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_149
timestamp 1644511149
transform 1 0 14812 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_161
timestamp 1644511149
transform 1 0 15916 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 1644511149
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_169
timestamp 1644511149
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_181
timestamp 1644511149
transform 1 0 17756 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_193
timestamp 1644511149
transform 1 0 18860 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_205
timestamp 1644511149
transform 1 0 19964 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_217
timestamp 1644511149
transform 1 0 21068 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_223
timestamp 1644511149
transform 1 0 21620 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_225
timestamp 1644511149
transform 1 0 21804 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_237
timestamp 1644511149
transform 1 0 22908 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_249
timestamp 1644511149
transform 1 0 24012 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_13_276
timestamp 1644511149
transform 1 0 26496 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_281
timestamp 1644511149
transform 1 0 26956 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_285
timestamp 1644511149
transform 1 0 27324 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_292
timestamp 1644511149
transform 1 0 27968 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_298
timestamp 1644511149
transform 1 0 28520 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_3
timestamp 1644511149
transform 1 0 1380 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_8
timestamp 1644511149
transform 1 0 1840 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_15
timestamp 1644511149
transform 1 0 2484 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_22
timestamp 1644511149
transform 1 0 3128 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_14_29
timestamp 1644511149
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_41
timestamp 1644511149
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_53
timestamp 1644511149
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_65
timestamp 1644511149
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp 1644511149
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1644511149
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_85
timestamp 1644511149
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_97
timestamp 1644511149
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_109
timestamp 1644511149
transform 1 0 11132 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_121
timestamp 1644511149
transform 1 0 12236 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_133
timestamp 1644511149
transform 1 0 13340 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1644511149
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_141
timestamp 1644511149
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_153
timestamp 1644511149
transform 1 0 15180 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_165
timestamp 1644511149
transform 1 0 16284 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_169
timestamp 1644511149
transform 1 0 16652 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_179
timestamp 1644511149
transform 1 0 17572 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_191
timestamp 1644511149
transform 1 0 18676 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_195
timestamp 1644511149
transform 1 0 19044 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_197
timestamp 1644511149
transform 1 0 19228 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_209
timestamp 1644511149
transform 1 0 20332 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_221
timestamp 1644511149
transform 1 0 21436 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_233
timestamp 1644511149
transform 1 0 22540 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_245
timestamp 1644511149
transform 1 0 23644 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_251
timestamp 1644511149
transform 1 0 24196 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_253
timestamp 1644511149
transform 1 0 24380 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_257
timestamp 1644511149
transform 1 0 24748 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_282
timestamp 1644511149
transform 1 0 27048 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_289
timestamp 1644511149
transform 1 0 27692 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_297
timestamp 1644511149
transform 1 0 28428 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_3
timestamp 1644511149
transform 1 0 1380 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_7
timestamp 1644511149
transform 1 0 1748 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_19
timestamp 1644511149
transform 1 0 2852 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_31
timestamp 1644511149
transform 1 0 3956 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_43
timestamp 1644511149
transform 1 0 5060 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1644511149
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_57
timestamp 1644511149
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_69
timestamp 1644511149
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_81
timestamp 1644511149
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_93
timestamp 1644511149
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_105
timestamp 1644511149
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1644511149
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_113
timestamp 1644511149
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_125
timestamp 1644511149
transform 1 0 12604 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_137
timestamp 1644511149
transform 1 0 13708 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_149
timestamp 1644511149
transform 1 0 14812 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_164
timestamp 1644511149
transform 1 0 16192 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_15_185
timestamp 1644511149
transform 1 0 18124 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_197
timestamp 1644511149
transform 1 0 19228 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_205
timestamp 1644511149
transform 1 0 19964 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_15_216
timestamp 1644511149
transform 1 0 20976 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_15_225
timestamp 1644511149
transform 1 0 21804 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_237
timestamp 1644511149
transform 1 0 22908 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_249
timestamp 1644511149
transform 1 0 24012 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_15_276
timestamp 1644511149
transform 1 0 26496 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_281
timestamp 1644511149
transform 1 0 26956 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_285
timestamp 1644511149
transform 1 0 27324 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_292
timestamp 1644511149
transform 1 0 27968 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_298
timestamp 1644511149
transform 1 0 28520 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_3
timestamp 1644511149
transform 1 0 1380 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_16_10
timestamp 1644511149
transform 1 0 2024 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_22
timestamp 1644511149
transform 1 0 3128 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_16_29
timestamp 1644511149
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_41
timestamp 1644511149
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_53
timestamp 1644511149
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_65
timestamp 1644511149
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp 1644511149
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1644511149
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_85
timestamp 1644511149
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_97
timestamp 1644511149
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_109
timestamp 1644511149
transform 1 0 11132 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_121
timestamp 1644511149
transform 1 0 12236 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_133
timestamp 1644511149
transform 1 0 13340 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 1644511149
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_141
timestamp 1644511149
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_153
timestamp 1644511149
transform 1 0 15180 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_16_159
timestamp 1644511149
transform 1 0 15732 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_16_170
timestamp 1644511149
transform 1 0 16744 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_16_192
timestamp 1644511149
transform 1 0 18768 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_197
timestamp 1644511149
transform 1 0 19228 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_214
timestamp 1644511149
transform 1 0 20792 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_16_221
timestamp 1644511149
transform 1 0 21436 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_233
timestamp 1644511149
transform 1 0 22540 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_245
timestamp 1644511149
transform 1 0 23644 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_251
timestamp 1644511149
transform 1 0 24196 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_253
timestamp 1644511149
transform 1 0 24380 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_265
timestamp 1644511149
transform 1 0 25484 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_270
timestamp 1644511149
transform 1 0 25944 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_295
timestamp 1644511149
transform 1 0 28244 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_3
timestamp 1644511149
transform 1 0 1380 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_25
timestamp 1644511149
transform 1 0 3404 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_37
timestamp 1644511149
transform 1 0 4508 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_49
timestamp 1644511149
transform 1 0 5612 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1644511149
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_57
timestamp 1644511149
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_69
timestamp 1644511149
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_81
timestamp 1644511149
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_93
timestamp 1644511149
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_105
timestamp 1644511149
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1644511149
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_113
timestamp 1644511149
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_125
timestamp 1644511149
transform 1 0 12604 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_137
timestamp 1644511149
transform 1 0 13708 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_149
timestamp 1644511149
transform 1 0 14812 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_161
timestamp 1644511149
transform 1 0 15916 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_167
timestamp 1644511149
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_169
timestamp 1644511149
transform 1 0 16652 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_175
timestamp 1644511149
transform 1 0 17204 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_182
timestamp 1644511149
transform 1 0 17848 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_190
timestamp 1644511149
transform 1 0 18584 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_197
timestamp 1644511149
transform 1 0 19228 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_206
timestamp 1644511149
transform 1 0 20056 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_215
timestamp 1644511149
transform 1 0 20884 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_223
timestamp 1644511149
transform 1 0 21620 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_225
timestamp 1644511149
transform 1 0 21804 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_233
timestamp 1644511149
transform 1 0 22540 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_239
timestamp 1644511149
transform 1 0 23092 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_252
timestamp 1644511149
transform 1 0 24288 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_17_261
timestamp 1644511149
transform 1 0 25116 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_265
timestamp 1644511149
transform 1 0 25484 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_271
timestamp 1644511149
transform 1 0 26036 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_279
timestamp 1644511149
transform 1 0 26772 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_281
timestamp 1644511149
transform 1 0 26956 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_286
timestamp 1644511149
transform 1 0 27416 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_293
timestamp 1644511149
transform 1 0 28060 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_3
timestamp 1644511149
transform 1 0 1380 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_7
timestamp 1644511149
transform 1 0 1748 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_19
timestamp 1644511149
transform 1 0 2852 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1644511149
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_29
timestamp 1644511149
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_41
timestamp 1644511149
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_53
timestamp 1644511149
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_65
timestamp 1644511149
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_77
timestamp 1644511149
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1644511149
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_85
timestamp 1644511149
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_97
timestamp 1644511149
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_109
timestamp 1644511149
transform 1 0 11132 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_121
timestamp 1644511149
transform 1 0 12236 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_133
timestamp 1644511149
transform 1 0 13340 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_139
timestamp 1644511149
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_141
timestamp 1644511149
transform 1 0 14076 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_153
timestamp 1644511149
transform 1 0 15180 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_18_160
timestamp 1644511149
transform 1 0 15824 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_18_172
timestamp 1644511149
transform 1 0 16928 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_178
timestamp 1644511149
transform 1 0 17480 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_190
timestamp 1644511149
transform 1 0 18584 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_18_200
timestamp 1644511149
transform 1 0 19504 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_212
timestamp 1644511149
transform 1 0 20608 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_216
timestamp 1644511149
transform 1 0 20976 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_220
timestamp 1644511149
transform 1 0 21344 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_248
timestamp 1644511149
transform 1 0 23920 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_253
timestamp 1644511149
transform 1 0 24380 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_276
timestamp 1644511149
transform 1 0 26496 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_284
timestamp 1644511149
transform 1 0 27232 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_291
timestamp 1644511149
transform 1 0 27876 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_3
timestamp 1644511149
transform 1 0 1380 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_19_8
timestamp 1644511149
transform 1 0 1840 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_20
timestamp 1644511149
transform 1 0 2944 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_32
timestamp 1644511149
transform 1 0 4048 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_44
timestamp 1644511149
transform 1 0 5152 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_57
timestamp 1644511149
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_69
timestamp 1644511149
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_81
timestamp 1644511149
transform 1 0 8556 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_93
timestamp 1644511149
transform 1 0 9660 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_105
timestamp 1644511149
transform 1 0 10764 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1644511149
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_113
timestamp 1644511149
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_125
timestamp 1644511149
transform 1 0 12604 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_137
timestamp 1644511149
transform 1 0 13708 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_145
timestamp 1644511149
transform 1 0 14444 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_164
timestamp 1644511149
transform 1 0 16192 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_169
timestamp 1644511149
transform 1 0 16652 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_175
timestamp 1644511149
transform 1 0 17204 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_181
timestamp 1644511149
transform 1 0 17756 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_193
timestamp 1644511149
transform 1 0 18860 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_205
timestamp 1644511149
transform 1 0 19964 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_213
timestamp 1644511149
transform 1 0 20700 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_219
timestamp 1644511149
transform 1 0 21252 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_223
timestamp 1644511149
transform 1 0 21620 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_241
timestamp 1644511149
transform 1 0 23276 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_247
timestamp 1644511149
transform 1 0 23828 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_257
timestamp 1644511149
transform 1 0 24748 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_265
timestamp 1644511149
transform 1 0 25484 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_276
timestamp 1644511149
transform 1 0 26496 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_288
timestamp 1644511149
transform 1 0 27600 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_295
timestamp 1644511149
transform 1 0 28244 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_3
timestamp 1644511149
transform 1 0 1380 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_7
timestamp 1644511149
transform 1 0 1748 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_11
timestamp 1644511149
transform 1 0 2116 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_23
timestamp 1644511149
transform 1 0 3220 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1644511149
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_29
timestamp 1644511149
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_41
timestamp 1644511149
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_53
timestamp 1644511149
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_65
timestamp 1644511149
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_77
timestamp 1644511149
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1644511149
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_85
timestamp 1644511149
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_97
timestamp 1644511149
transform 1 0 10028 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_109
timestamp 1644511149
transform 1 0 11132 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_121
timestamp 1644511149
transform 1 0 12236 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_133
timestamp 1644511149
transform 1 0 13340 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_139
timestamp 1644511149
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_144
timestamp 1644511149
transform 1 0 14352 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_152
timestamp 1644511149
transform 1 0 15088 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_160
timestamp 1644511149
transform 1 0 15824 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_167
timestamp 1644511149
transform 1 0 16468 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_171
timestamp 1644511149
transform 1 0 16836 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_188
timestamp 1644511149
transform 1 0 18400 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_20_197
timestamp 1644511149
transform 1 0 19228 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_203
timestamp 1644511149
transform 1 0 19780 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_207
timestamp 1644511149
transform 1 0 20148 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_215
timestamp 1644511149
transform 1 0 20884 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_226
timestamp 1644511149
transform 1 0 21896 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_20_240
timestamp 1644511149
transform 1 0 23184 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_253
timestamp 1644511149
transform 1 0 24380 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_260
timestamp 1644511149
transform 1 0 25024 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_270
timestamp 1644511149
transform 1 0 25944 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_295
timestamp 1644511149
transform 1 0 28244 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_3
timestamp 1644511149
transform 1 0 1380 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_25
timestamp 1644511149
transform 1 0 3404 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_37
timestamp 1644511149
transform 1 0 4508 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_49
timestamp 1644511149
transform 1 0 5612 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1644511149
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_57
timestamp 1644511149
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_69
timestamp 1644511149
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_81
timestamp 1644511149
transform 1 0 8556 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_93
timestamp 1644511149
transform 1 0 9660 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_105
timestamp 1644511149
transform 1 0 10764 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 1644511149
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_113
timestamp 1644511149
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_125
timestamp 1644511149
transform 1 0 12604 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_21_149
timestamp 1644511149
transform 1 0 14812 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_21_160
timestamp 1644511149
transform 1 0 15824 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_21_169
timestamp 1644511149
transform 1 0 16652 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_178
timestamp 1644511149
transform 1 0 17480 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_185
timestamp 1644511149
transform 1 0 18124 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_189
timestamp 1644511149
transform 1 0 18492 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_193
timestamp 1644511149
transform 1 0 18860 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_199
timestamp 1644511149
transform 1 0 19412 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_216
timestamp 1644511149
transform 1 0 20976 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_21_225
timestamp 1644511149
transform 1 0 21804 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_237
timestamp 1644511149
transform 1 0 22908 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_21_244
timestamp 1644511149
transform 1 0 23552 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_21_256
timestamp 1644511149
transform 1 0 24656 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_264
timestamp 1644511149
transform 1 0 25392 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_271
timestamp 1644511149
transform 1 0 26036 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_279
timestamp 1644511149
transform 1 0 26772 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_286
timestamp 1644511149
transform 1 0 27416 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_293
timestamp 1644511149
transform 1 0 28060 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_22_24
timestamp 1644511149
transform 1 0 3312 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_29
timestamp 1644511149
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_41
timestamp 1644511149
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_53
timestamp 1644511149
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_65
timestamp 1644511149
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_77
timestamp 1644511149
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1644511149
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_85
timestamp 1644511149
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_97
timestamp 1644511149
transform 1 0 10028 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_109
timestamp 1644511149
transform 1 0 11132 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_121
timestamp 1644511149
transform 1 0 12236 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_133
timestamp 1644511149
transform 1 0 13340 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_139
timestamp 1644511149
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_141
timestamp 1644511149
transform 1 0 14076 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_149
timestamp 1644511149
transform 1 0 14812 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_157
timestamp 1644511149
transform 1 0 15548 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_164
timestamp 1644511149
transform 1 0 16192 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_176
timestamp 1644511149
transform 1 0 17296 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_188
timestamp 1644511149
transform 1 0 18400 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_22_197
timestamp 1644511149
transform 1 0 19228 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_22_208
timestamp 1644511149
transform 1 0 20240 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_22_232
timestamp 1644511149
transform 1 0 22448 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_241
timestamp 1644511149
transform 1 0 23276 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_249
timestamp 1644511149
transform 1 0 24012 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_262
timestamp 1644511149
transform 1 0 25208 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_270
timestamp 1644511149
transform 1 0 25944 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_295
timestamp 1644511149
transform 1 0 28244 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_3
timestamp 1644511149
transform 1 0 1380 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_10
timestamp 1644511149
transform 1 0 2024 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_14
timestamp 1644511149
transform 1 0 2392 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_36
timestamp 1644511149
transform 1 0 4416 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_48
timestamp 1644511149
transform 1 0 5520 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_23_57
timestamp 1644511149
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_69
timestamp 1644511149
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_81
timestamp 1644511149
transform 1 0 8556 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_93
timestamp 1644511149
transform 1 0 9660 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_105
timestamp 1644511149
transform 1 0 10764 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp 1644511149
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_113
timestamp 1644511149
transform 1 0 11500 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_117
timestamp 1644511149
transform 1 0 11868 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_134
timestamp 1644511149
transform 1 0 13432 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_146
timestamp 1644511149
transform 1 0 14536 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_150
timestamp 1644511149
transform 1 0 14904 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_154
timestamp 1644511149
transform 1 0 15272 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_166
timestamp 1644511149
transform 1 0 16376 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_23_169
timestamp 1644511149
transform 1 0 16652 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_181
timestamp 1644511149
transform 1 0 17756 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_199
timestamp 1644511149
transform 1 0 19412 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_23_216
timestamp 1644511149
transform 1 0 20976 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_225
timestamp 1644511149
transform 1 0 21804 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_231
timestamp 1644511149
transform 1 0 22356 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_251
timestamp 1644511149
transform 1 0 24196 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_23_269
timestamp 1644511149
transform 1 0 25852 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_276
timestamp 1644511149
transform 1 0 26496 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_288
timestamp 1644511149
transform 1 0 27600 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_295
timestamp 1644511149
transform 1 0 28244 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_3
timestamp 1644511149
transform 1 0 1380 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_7
timestamp 1644511149
transform 1 0 1748 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_19
timestamp 1644511149
transform 1 0 2852 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1644511149
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_32
timestamp 1644511149
transform 1 0 4048 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_44
timestamp 1644511149
transform 1 0 5152 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_56
timestamp 1644511149
transform 1 0 6256 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_68
timestamp 1644511149
transform 1 0 7360 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_80
timestamp 1644511149
transform 1 0 8464 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_85
timestamp 1644511149
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_97
timestamp 1644511149
transform 1 0 10028 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_109
timestamp 1644511149
transform 1 0 11132 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_117
timestamp 1644511149
transform 1 0 11868 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_123
timestamp 1644511149
transform 1 0 12420 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_130
timestamp 1644511149
transform 1 0 13064 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_138
timestamp 1644511149
transform 1 0 13800 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_147
timestamp 1644511149
transform 1 0 14628 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_154
timestamp 1644511149
transform 1 0 15272 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_161
timestamp 1644511149
transform 1 0 15916 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_179
timestamp 1644511149
transform 1 0 17572 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_192
timestamp 1644511149
transform 1 0 18768 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_204
timestamp 1644511149
transform 1 0 19872 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_214
timestamp 1644511149
transform 1 0 20792 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_226
timestamp 1644511149
transform 1 0 21896 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_232
timestamp 1644511149
transform 1 0 22448 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_242
timestamp 1644511149
transform 1 0 23368 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_250
timestamp 1644511149
transform 1 0 24104 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_253
timestamp 1644511149
transform 1 0 24380 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_258
timestamp 1644511149
transform 1 0 24840 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_270
timestamp 1644511149
transform 1 0 25944 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_295
timestamp 1644511149
transform 1 0 28244 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_25_3
timestamp 1644511149
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_18
timestamp 1644511149
transform 1 0 2760 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_30
timestamp 1644511149
transform 1 0 3864 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_42
timestamp 1644511149
transform 1 0 4968 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_54
timestamp 1644511149
transform 1 0 6072 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_25_57
timestamp 1644511149
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_69
timestamp 1644511149
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_81
timestamp 1644511149
transform 1 0 8556 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_93
timestamp 1644511149
transform 1 0 9660 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_105
timestamp 1644511149
transform 1 0 10764 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp 1644511149
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_113
timestamp 1644511149
transform 1 0 11500 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_121
timestamp 1644511149
transform 1 0 12236 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_131
timestamp 1644511149
transform 1 0 13156 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_143
timestamp 1644511149
transform 1 0 14260 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_151
timestamp 1644511149
transform 1 0 14996 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_25_159
timestamp 1644511149
transform 1 0 15732 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_167
timestamp 1644511149
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_169
timestamp 1644511149
transform 1 0 16652 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_173
timestamp 1644511149
transform 1 0 17020 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_180
timestamp 1644511149
transform 1 0 17664 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_192
timestamp 1644511149
transform 1 0 18768 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_25_204
timestamp 1644511149
transform 1 0 19872 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_216
timestamp 1644511149
transform 1 0 20976 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_25_225
timestamp 1644511149
transform 1 0 21804 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_237
timestamp 1644511149
transform 1 0 22908 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_249
timestamp 1644511149
transform 1 0 24012 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_257
timestamp 1644511149
transform 1 0 24748 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_261
timestamp 1644511149
transform 1 0 25116 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_272
timestamp 1644511149
transform 1 0 26128 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_25_285
timestamp 1644511149
transform 1 0 27324 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_25_295
timestamp 1644511149
transform 1 0 28244 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_3
timestamp 1644511149
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_15
timestamp 1644511149
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1644511149
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_29
timestamp 1644511149
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_41
timestamp 1644511149
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_53
timestamp 1644511149
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_65
timestamp 1644511149
transform 1 0 7084 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_77
timestamp 1644511149
transform 1 0 8188 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 1644511149
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_85
timestamp 1644511149
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_97
timestamp 1644511149
transform 1 0 10028 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_109
timestamp 1644511149
transform 1 0 11132 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_121
timestamp 1644511149
transform 1 0 12236 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_133
timestamp 1644511149
transform 1 0 13340 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_139
timestamp 1644511149
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_148
timestamp 1644511149
transform 1 0 14720 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_152
timestamp 1644511149
transform 1 0 15088 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_160
timestamp 1644511149
transform 1 0 15824 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_180
timestamp 1644511149
transform 1 0 17664 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_189
timestamp 1644511149
transform 1 0 18492 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_195
timestamp 1644511149
transform 1 0 19044 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_200
timestamp 1644511149
transform 1 0 19504 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_26_212
timestamp 1644511149
transform 1 0 20608 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_220
timestamp 1644511149
transform 1 0 21344 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_232
timestamp 1644511149
transform 1 0 22448 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_247
timestamp 1644511149
transform 1 0 23828 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_251
timestamp 1644511149
transform 1 0 24196 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_253
timestamp 1644511149
transform 1 0 24380 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_257
timestamp 1644511149
transform 1 0 24748 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_261
timestamp 1644511149
transform 1 0 25116 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_268
timestamp 1644511149
transform 1 0 25760 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_26_295
timestamp 1644511149
transform 1 0 28244 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_3
timestamp 1644511149
transform 1 0 1380 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_27_8
timestamp 1644511149
transform 1 0 1840 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_20
timestamp 1644511149
transform 1 0 2944 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_32
timestamp 1644511149
transform 1 0 4048 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_44
timestamp 1644511149
transform 1 0 5152 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_57
timestamp 1644511149
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_69
timestamp 1644511149
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_81
timestamp 1644511149
transform 1 0 8556 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_93
timestamp 1644511149
transform 1 0 9660 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_105
timestamp 1644511149
transform 1 0 10764 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_111
timestamp 1644511149
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_113
timestamp 1644511149
transform 1 0 11500 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_27_130
timestamp 1644511149
transform 1 0 13064 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_140
timestamp 1644511149
transform 1 0 13984 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_152
timestamp 1644511149
transform 1 0 15088 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_27_162
timestamp 1644511149
transform 1 0 16008 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_27_174
timestamp 1644511149
transform 1 0 17112 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_186
timestamp 1644511149
transform 1 0 18216 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_198
timestamp 1644511149
transform 1 0 19320 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_206
timestamp 1644511149
transform 1 0 20056 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_210
timestamp 1644511149
transform 1 0 20424 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_220
timestamp 1644511149
transform 1 0 21344 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_27_231
timestamp 1644511149
transform 1 0 22356 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_252
timestamp 1644511149
transform 1 0 24288 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_264
timestamp 1644511149
transform 1 0 25392 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_27_273
timestamp 1644511149
transform 1 0 26220 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_279
timestamp 1644511149
transform 1 0 26772 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_288
timestamp 1644511149
transform 1 0 27600 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_295
timestamp 1644511149
transform 1 0 28244 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_24
timestamp 1644511149
transform 1 0 3312 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_29
timestamp 1644511149
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_41
timestamp 1644511149
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_53
timestamp 1644511149
transform 1 0 5980 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_65
timestamp 1644511149
transform 1 0 7084 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_77
timestamp 1644511149
transform 1 0 8188 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_83
timestamp 1644511149
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_85
timestamp 1644511149
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_97
timestamp 1644511149
transform 1 0 10028 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_109
timestamp 1644511149
transform 1 0 11132 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_113
timestamp 1644511149
transform 1 0 11500 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_133
timestamp 1644511149
transform 1 0 13340 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_139
timestamp 1644511149
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_150
timestamp 1644511149
transform 1 0 14904 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_28_158
timestamp 1644511149
transform 1 0 15640 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_168
timestamp 1644511149
transform 1 0 16560 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_175
timestamp 1644511149
transform 1 0 17204 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_191
timestamp 1644511149
transform 1 0 18676 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_195
timestamp 1644511149
transform 1 0 19044 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_28_197
timestamp 1644511149
transform 1 0 19228 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_28_219
timestamp 1644511149
transform 1 0 21252 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_28_243
timestamp 1644511149
transform 1 0 23460 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_251
timestamp 1644511149
transform 1 0 24196 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_269
timestamp 1644511149
transform 1 0 25852 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_273
timestamp 1644511149
transform 1 0 26220 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_295
timestamp 1644511149
transform 1 0 28244 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_29_6
timestamp 1644511149
transform 1 0 1656 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_18
timestamp 1644511149
transform 1 0 2760 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_30
timestamp 1644511149
transform 1 0 3864 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_42
timestamp 1644511149
transform 1 0 4968 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_54
timestamp 1644511149
transform 1 0 6072 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_29_57
timestamp 1644511149
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_69
timestamp 1644511149
transform 1 0 7452 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_81
timestamp 1644511149
transform 1 0 8556 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_93
timestamp 1644511149
transform 1 0 9660 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_105
timestamp 1644511149
transform 1 0 10764 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_111
timestamp 1644511149
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_29_113
timestamp 1644511149
transform 1 0 11500 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_119
timestamp 1644511149
transform 1 0 12052 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_29_125
timestamp 1644511149
transform 1 0 12604 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_131
timestamp 1644511149
transform 1 0 13156 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_138
timestamp 1644511149
transform 1 0 13800 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_29_150
timestamp 1644511149
transform 1 0 14904 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_162
timestamp 1644511149
transform 1 0 16008 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_29_174
timestamp 1644511149
transform 1 0 17112 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_182
timestamp 1644511149
transform 1 0 17848 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_29_200
timestamp 1644511149
transform 1 0 19504 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_218
timestamp 1644511149
transform 1 0 21160 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_29_231
timestamp 1644511149
transform 1 0 22356 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_241
timestamp 1644511149
transform 1 0 23276 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_250
timestamp 1644511149
transform 1 0 24104 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_258
timestamp 1644511149
transform 1 0 24840 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_29_269
timestamp 1644511149
transform 1 0 25852 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_277
timestamp 1644511149
transform 1 0 26588 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_284
timestamp 1644511149
transform 1 0 27232 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_288
timestamp 1644511149
transform 1 0 27600 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_29_292
timestamp 1644511149
transform 1 0 27968 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_298
timestamp 1644511149
transform 1 0 28520 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_3
timestamp 1644511149
transform 1 0 1380 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_10
timestamp 1644511149
transform 1 0 2024 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_17
timestamp 1644511149
transform 1 0 2668 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_30_25
timestamp 1644511149
transform 1 0 3404 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_30_29
timestamp 1644511149
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_41
timestamp 1644511149
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_53
timestamp 1644511149
transform 1 0 5980 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_65
timestamp 1644511149
transform 1 0 7084 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_77
timestamp 1644511149
transform 1 0 8188 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_83
timestamp 1644511149
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_85
timestamp 1644511149
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_97
timestamp 1644511149
transform 1 0 10028 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_109
timestamp 1644511149
transform 1 0 11132 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_121
timestamp 1644511149
transform 1 0 12236 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_133
timestamp 1644511149
transform 1 0 13340 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_139
timestamp 1644511149
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_141
timestamp 1644511149
transform 1 0 14076 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_153
timestamp 1644511149
transform 1 0 15180 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_170
timestamp 1644511149
transform 1 0 16744 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_181
timestamp 1644511149
transform 1 0 17756 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_188
timestamp 1644511149
transform 1 0 18400 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_30_197
timestamp 1644511149
transform 1 0 19228 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_209
timestamp 1644511149
transform 1 0 20332 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_30_221
timestamp 1644511149
transform 1 0 21436 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_225
timestamp 1644511149
transform 1 0 21804 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_232
timestamp 1644511149
transform 1 0 22448 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_244
timestamp 1644511149
transform 1 0 23552 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_30_253
timestamp 1644511149
transform 1 0 24380 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_265
timestamp 1644511149
transform 1 0 25484 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_273
timestamp 1644511149
transform 1 0 26220 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_295
timestamp 1644511149
transform 1 0 28244 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_24
timestamp 1644511149
transform 1 0 3312 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_36
timestamp 1644511149
transform 1 0 4416 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_48
timestamp 1644511149
transform 1 0 5520 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_31_57
timestamp 1644511149
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_69
timestamp 1644511149
transform 1 0 7452 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_81
timestamp 1644511149
transform 1 0 8556 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_93
timestamp 1644511149
transform 1 0 9660 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_105
timestamp 1644511149
transform 1 0 10764 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_111
timestamp 1644511149
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_113
timestamp 1644511149
transform 1 0 11500 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_125
timestamp 1644511149
transform 1 0 12604 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_137
timestamp 1644511149
transform 1 0 13708 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_145
timestamp 1644511149
transform 1 0 14444 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_31_151
timestamp 1644511149
transform 1 0 14996 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_163
timestamp 1644511149
transform 1 0 16100 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_167
timestamp 1644511149
transform 1 0 16468 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_31_169
timestamp 1644511149
transform 1 0 16652 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_177
timestamp 1644511149
transform 1 0 17388 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_185
timestamp 1644511149
transform 1 0 18124 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_197
timestamp 1644511149
transform 1 0 19228 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_31_209
timestamp 1644511149
transform 1 0 20332 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_214
timestamp 1644511149
transform 1 0 20792 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_222
timestamp 1644511149
transform 1 0 21528 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_31_225
timestamp 1644511149
transform 1 0 21804 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_237
timestamp 1644511149
transform 1 0 22908 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_31_249
timestamp 1644511149
transform 1 0 24012 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_257
timestamp 1644511149
transform 1 0 24748 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_264
timestamp 1644511149
transform 1 0 25392 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_272
timestamp 1644511149
transform 1 0 26128 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_276
timestamp 1644511149
transform 1 0 26496 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_31_281
timestamp 1644511149
transform 1 0 26956 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_287
timestamp 1644511149
transform 1 0 27508 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_294
timestamp 1644511149
transform 1 0 28152 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_298
timestamp 1644511149
transform 1 0 28520 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_3
timestamp 1644511149
transform 1 0 1380 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_7
timestamp 1644511149
transform 1 0 1748 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_14
timestamp 1644511149
transform 1 0 2392 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_21
timestamp 1644511149
transform 1 0 3036 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1644511149
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_29
timestamp 1644511149
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_41
timestamp 1644511149
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_53
timestamp 1644511149
transform 1 0 5980 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_65
timestamp 1644511149
transform 1 0 7084 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_77
timestamp 1644511149
transform 1 0 8188 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_83
timestamp 1644511149
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_85
timestamp 1644511149
transform 1 0 8924 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_97
timestamp 1644511149
transform 1 0 10028 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_109
timestamp 1644511149
transform 1 0 11132 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_130
timestamp 1644511149
transform 1 0 13064 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_138
timestamp 1644511149
transform 1 0 13800 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_32_141
timestamp 1644511149
transform 1 0 14076 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_145
timestamp 1644511149
transform 1 0 14444 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_154
timestamp 1644511149
transform 1 0 15272 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_162
timestamp 1644511149
transform 1 0 16008 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_32_174
timestamp 1644511149
transform 1 0 17112 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_182
timestamp 1644511149
transform 1 0 17848 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_190
timestamp 1644511149
transform 1 0 18584 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_32_197
timestamp 1644511149
transform 1 0 19228 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_32_205
timestamp 1644511149
transform 1 0 19964 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_213
timestamp 1644511149
transform 1 0 20700 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_217
timestamp 1644511149
transform 1 0 21068 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_222
timestamp 1644511149
transform 1 0 21528 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_226
timestamp 1644511149
transform 1 0 21896 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_233
timestamp 1644511149
transform 1 0 22540 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_239
timestamp 1644511149
transform 1 0 23092 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_245
timestamp 1644511149
transform 1 0 23644 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_251
timestamp 1644511149
transform 1 0 24196 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_253
timestamp 1644511149
transform 1 0 24380 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_270
timestamp 1644511149
transform 1 0 25944 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_295
timestamp 1644511149
transform 1 0 28244 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_3
timestamp 1644511149
transform 1 0 1380 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_11
timestamp 1644511149
transform 1 0 2116 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_33_34
timestamp 1644511149
transform 1 0 4232 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_46
timestamp 1644511149
transform 1 0 5336 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_54
timestamp 1644511149
transform 1 0 6072 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_33_57
timestamp 1644511149
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_69
timestamp 1644511149
transform 1 0 7452 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_81
timestamp 1644511149
transform 1 0 8556 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_93
timestamp 1644511149
transform 1 0 9660 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_105
timestamp 1644511149
transform 1 0 10764 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_111
timestamp 1644511149
transform 1 0 11316 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_113
timestamp 1644511149
transform 1 0 11500 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_117
timestamp 1644511149
transform 1 0 11868 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_134
timestamp 1644511149
transform 1 0 13432 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_154
timestamp 1644511149
transform 1 0 15272 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_163
timestamp 1644511149
transform 1 0 16100 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_167
timestamp 1644511149
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_169
timestamp 1644511149
transform 1 0 16652 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_177
timestamp 1644511149
transform 1 0 17388 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_185
timestamp 1644511149
transform 1 0 18124 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_193
timestamp 1644511149
transform 1 0 18860 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_201
timestamp 1644511149
transform 1 0 19596 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_218
timestamp 1644511149
transform 1 0 21160 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_33_225
timestamp 1644511149
transform 1 0 21804 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_229
timestamp 1644511149
transform 1 0 22172 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_239
timestamp 1644511149
transform 1 0 23092 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_259
timestamp 1644511149
transform 1 0 24932 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_263
timestamp 1644511149
transform 1 0 25300 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_273
timestamp 1644511149
transform 1 0 26220 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_279
timestamp 1644511149
transform 1 0 26772 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_281
timestamp 1644511149
transform 1 0 26956 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_286
timestamp 1644511149
transform 1 0 27416 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_290
timestamp 1644511149
transform 1 0 27784 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_294
timestamp 1644511149
transform 1 0 28152 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_298
timestamp 1644511149
transform 1 0 28520 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_24
timestamp 1644511149
transform 1 0 3312 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_34_29
timestamp 1644511149
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_41
timestamp 1644511149
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_53
timestamp 1644511149
transform 1 0 5980 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_65
timestamp 1644511149
transform 1 0 7084 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_77
timestamp 1644511149
transform 1 0 8188 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_83
timestamp 1644511149
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_85
timestamp 1644511149
transform 1 0 8924 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_97
timestamp 1644511149
transform 1 0 10028 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_109
timestamp 1644511149
transform 1 0 11132 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_117
timestamp 1644511149
transform 1 0 11868 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_124
timestamp 1644511149
transform 1 0 12512 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_131
timestamp 1644511149
transform 1 0 13156 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_139
timestamp 1644511149
transform 1 0 13892 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_144
timestamp 1644511149
transform 1 0 14352 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_148
timestamp 1644511149
transform 1 0 14720 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_154
timestamp 1644511149
transform 1 0 15272 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_161
timestamp 1644511149
transform 1 0 15916 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_169
timestamp 1644511149
transform 1 0 16652 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_34_175
timestamp 1644511149
transform 1 0 17204 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_181
timestamp 1644511149
transform 1 0 17756 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_34_188
timestamp 1644511149
transform 1 0 18400 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_34_204
timestamp 1644511149
transform 1 0 19872 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_212
timestamp 1644511149
transform 1 0 20608 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_217
timestamp 1644511149
transform 1 0 21068 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_237
timestamp 1644511149
transform 1 0 22908 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_244
timestamp 1644511149
transform 1 0 23552 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_34_253
timestamp 1644511149
transform 1 0 24380 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_266
timestamp 1644511149
transform 1 0 25576 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_34_295
timestamp 1644511149
transform 1 0 28244 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_3
timestamp 1644511149
transform 1 0 1380 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_35_12
timestamp 1644511149
transform 1 0 2208 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_24
timestamp 1644511149
transform 1 0 3312 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_36
timestamp 1644511149
transform 1 0 4416 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_48
timestamp 1644511149
transform 1 0 5520 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_35_57
timestamp 1644511149
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_69
timestamp 1644511149
transform 1 0 7452 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_81
timestamp 1644511149
transform 1 0 8556 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_93
timestamp 1644511149
transform 1 0 9660 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_105
timestamp 1644511149
transform 1 0 10764 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_111
timestamp 1644511149
transform 1 0 11316 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_113
timestamp 1644511149
transform 1 0 11500 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_125
timestamp 1644511149
transform 1 0 12604 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_137
timestamp 1644511149
transform 1 0 13708 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_35_149
timestamp 1644511149
transform 1 0 14812 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_35_158
timestamp 1644511149
transform 1 0 15640 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_166
timestamp 1644511149
transform 1 0 16376 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_169
timestamp 1644511149
transform 1 0 16652 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_173
timestamp 1644511149
transform 1 0 17020 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_178
timestamp 1644511149
transform 1 0 17480 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_189
timestamp 1644511149
transform 1 0 18492 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_197
timestamp 1644511149
transform 1 0 19228 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_205
timestamp 1644511149
transform 1 0 19964 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_213
timestamp 1644511149
transform 1 0 20700 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_220
timestamp 1644511149
transform 1 0 21344 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_35_231
timestamp 1644511149
transform 1 0 22356 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_243
timestamp 1644511149
transform 1 0 23460 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_247
timestamp 1644511149
transform 1 0 23828 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_251
timestamp 1644511149
transform 1 0 24196 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_276
timestamp 1644511149
transform 1 0 26496 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_281
timestamp 1644511149
transform 1 0 26956 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_35_290
timestamp 1644511149
transform 1 0 27784 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_298
timestamp 1644511149
transform 1 0 28520 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_3
timestamp 1644511149
transform 1 0 1380 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_36_8
timestamp 1644511149
transform 1 0 1840 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_20
timestamp 1644511149
transform 1 0 2944 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_36_29
timestamp 1644511149
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_41
timestamp 1644511149
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_53
timestamp 1644511149
transform 1 0 5980 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_65
timestamp 1644511149
transform 1 0 7084 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_77
timestamp 1644511149
transform 1 0 8188 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_83
timestamp 1644511149
transform 1 0 8740 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_85
timestamp 1644511149
transform 1 0 8924 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_97
timestamp 1644511149
transform 1 0 10028 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_109
timestamp 1644511149
transform 1 0 11132 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_121
timestamp 1644511149
transform 1 0 12236 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_133
timestamp 1644511149
transform 1 0 13340 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_139
timestamp 1644511149
transform 1 0 13892 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_144
timestamp 1644511149
transform 1 0 14352 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_156
timestamp 1644511149
transform 1 0 15456 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_168
timestamp 1644511149
transform 1 0 16560 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_180
timestamp 1644511149
transform 1 0 17664 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_192
timestamp 1644511149
transform 1 0 18768 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_197
timestamp 1644511149
transform 1 0 19228 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_201
timestamp 1644511149
transform 1 0 19596 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_206
timestamp 1644511149
transform 1 0 20056 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_36_217
timestamp 1644511149
transform 1 0 21068 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_229
timestamp 1644511149
transform 1 0 22172 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_36_238
timestamp 1644511149
transform 1 0 23000 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_244
timestamp 1644511149
transform 1 0 23552 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_248
timestamp 1644511149
transform 1 0 23920 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_256
timestamp 1644511149
transform 1 0 24656 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_266
timestamp 1644511149
transform 1 0 25576 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_36_295
timestamp 1644511149
transform 1 0 28244 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_37_3
timestamp 1644511149
transform 1 0 1380 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_15
timestamp 1644511149
transform 1 0 2484 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_27
timestamp 1644511149
transform 1 0 3588 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_39
timestamp 1644511149
transform 1 0 4692 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_51
timestamp 1644511149
transform 1 0 5796 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_55
timestamp 1644511149
transform 1 0 6164 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_57
timestamp 1644511149
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_69
timestamp 1644511149
transform 1 0 7452 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_81
timestamp 1644511149
transform 1 0 8556 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_93
timestamp 1644511149
transform 1 0 9660 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_105
timestamp 1644511149
transform 1 0 10764 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_111
timestamp 1644511149
transform 1 0 11316 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_113
timestamp 1644511149
transform 1 0 11500 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_37_121
timestamp 1644511149
transform 1 0 12236 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_37_129
timestamp 1644511149
transform 1 0 12972 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_37_149
timestamp 1644511149
transform 1 0 14812 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_161
timestamp 1644511149
transform 1 0 15916 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_167
timestamp 1644511149
transform 1 0 16468 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_169
timestamp 1644511149
transform 1 0 16652 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_181
timestamp 1644511149
transform 1 0 17756 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_196
timestamp 1644511149
transform 1 0 19136 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_204
timestamp 1644511149
transform 1 0 19872 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_37_209
timestamp 1644511149
transform 1 0 20332 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_37_221
timestamp 1644511149
transform 1 0 21436 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_37_230
timestamp 1644511149
transform 1 0 22264 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_37_252
timestamp 1644511149
transform 1 0 24288 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_258
timestamp 1644511149
transform 1 0 24840 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_275
timestamp 1644511149
transform 1 0 26404 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_279
timestamp 1644511149
transform 1 0 26772 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_284
timestamp 1644511149
transform 1 0 27232 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_288
timestamp 1644511149
transform 1 0 27600 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_37_292
timestamp 1644511149
transform 1 0 27968 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_298
timestamp 1644511149
transform 1 0 28520 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_3
timestamp 1644511149
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_15
timestamp 1644511149
transform 1 0 2484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 1644511149
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_29
timestamp 1644511149
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_41
timestamp 1644511149
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_53
timestamp 1644511149
transform 1 0 5980 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_65
timestamp 1644511149
transform 1 0 7084 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_77
timestamp 1644511149
transform 1 0 8188 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_83
timestamp 1644511149
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_85
timestamp 1644511149
transform 1 0 8924 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_97
timestamp 1644511149
transform 1 0 10028 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_109
timestamp 1644511149
transform 1 0 11132 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_38_117
timestamp 1644511149
transform 1 0 11868 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_38_136
timestamp 1644511149
transform 1 0 13616 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_38_141
timestamp 1644511149
transform 1 0 14076 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_38_153
timestamp 1644511149
transform 1 0 15180 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_162
timestamp 1644511149
transform 1 0 16008 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_172
timestamp 1644511149
transform 1 0 16928 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_181
timestamp 1644511149
transform 1 0 17756 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_189
timestamp 1644511149
transform 1 0 18492 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_195
timestamp 1644511149
transform 1 0 19044 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_38_205
timestamp 1644511149
transform 1 0 19964 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_211
timestamp 1644511149
transform 1 0 20516 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_217
timestamp 1644511149
transform 1 0 21068 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_226
timestamp 1644511149
transform 1 0 21896 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_235
timestamp 1644511149
transform 1 0 22724 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_248
timestamp 1644511149
transform 1 0 23920 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_253
timestamp 1644511149
transform 1 0 24380 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_259
timestamp 1644511149
transform 1 0 24932 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_267
timestamp 1644511149
transform 1 0 25668 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_283
timestamp 1644511149
transform 1 0 27140 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_38_294
timestamp 1644511149
transform 1 0 28152 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_298
timestamp 1644511149
transform 1 0 28520 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_3
timestamp 1644511149
transform 1 0 1380 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_15
timestamp 1644511149
transform 1 0 2484 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_27
timestamp 1644511149
transform 1 0 3588 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_43
timestamp 1644511149
transform 1 0 5060 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_39_55
timestamp 1644511149
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_57
timestamp 1644511149
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_69
timestamp 1644511149
transform 1 0 7452 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_81
timestamp 1644511149
transform 1 0 8556 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_93
timestamp 1644511149
transform 1 0 9660 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_105
timestamp 1644511149
transform 1 0 10764 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_111
timestamp 1644511149
transform 1 0 11316 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_113
timestamp 1644511149
transform 1 0 11500 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_39_130
timestamp 1644511149
transform 1 0 13064 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_142
timestamp 1644511149
transform 1 0 14168 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_39_164
timestamp 1644511149
transform 1 0 16192 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_169
timestamp 1644511149
transform 1 0 16652 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_173
timestamp 1644511149
transform 1 0 17020 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_180
timestamp 1644511149
transform 1 0 17664 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_188
timestamp 1644511149
transform 1 0 18400 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_39_205
timestamp 1644511149
transform 1 0 19964 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_211
timestamp 1644511149
transform 1 0 20516 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_219
timestamp 1644511149
transform 1 0 21252 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_223
timestamp 1644511149
transform 1 0 21620 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_230
timestamp 1644511149
transform 1 0 22264 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_39_238
timestamp 1644511149
transform 1 0 23000 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_250
timestamp 1644511149
transform 1 0 24104 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_39_262
timestamp 1644511149
transform 1 0 25208 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_276
timestamp 1644511149
transform 1 0 26496 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_281
timestamp 1644511149
transform 1 0 26956 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_291
timestamp 1644511149
transform 1 0 27876 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_40_6
timestamp 1644511149
transform 1 0 1656 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_18
timestamp 1644511149
transform 1 0 2760 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_26
timestamp 1644511149
transform 1 0 3496 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_40_29
timestamp 1644511149
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_50
timestamp 1644511149
transform 1 0 5704 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_62
timestamp 1644511149
transform 1 0 6808 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_74
timestamp 1644511149
transform 1 0 7912 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_82
timestamp 1644511149
transform 1 0 8648 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_40_85
timestamp 1644511149
transform 1 0 8924 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_97
timestamp 1644511149
transform 1 0 10028 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_109
timestamp 1644511149
transform 1 0 11132 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_40_117
timestamp 1644511149
transform 1 0 11868 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_40_123
timestamp 1644511149
transform 1 0 12420 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_135
timestamp 1644511149
transform 1 0 13524 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_139
timestamp 1644511149
transform 1 0 13892 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_40_141
timestamp 1644511149
transform 1 0 14076 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_40_149
timestamp 1644511149
transform 1 0 14812 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_40_155
timestamp 1644511149
transform 1 0 15364 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_164
timestamp 1644511149
transform 1 0 16192 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_174
timestamp 1644511149
transform 1 0 17112 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_180
timestamp 1644511149
transform 1 0 17664 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_191
timestamp 1644511149
transform 1 0 18676 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_195
timestamp 1644511149
transform 1 0 19044 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_197
timestamp 1644511149
transform 1 0 19228 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_215
timestamp 1644511149
transform 1 0 20884 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_222
timestamp 1644511149
transform 1 0 21528 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_228
timestamp 1644511149
transform 1 0 22080 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_233
timestamp 1644511149
transform 1 0 22540 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_245
timestamp 1644511149
transform 1 0 23644 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_251
timestamp 1644511149
transform 1 0 24196 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_253
timestamp 1644511149
transform 1 0 24380 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_257
timestamp 1644511149
transform 1 0 24748 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_270
timestamp 1644511149
transform 1 0 25944 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_295
timestamp 1644511149
transform 1 0 28244 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_41_3
timestamp 1644511149
transform 1 0 1380 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_41_9
timestamp 1644511149
transform 1 0 1932 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_21
timestamp 1644511149
transform 1 0 3036 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_29
timestamp 1644511149
transform 1 0 3772 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_36
timestamp 1644511149
transform 1 0 4416 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_52
timestamp 1644511149
transform 1 0 5888 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_41_63
timestamp 1644511149
transform 1 0 6900 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_75
timestamp 1644511149
transform 1 0 8004 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_87
timestamp 1644511149
transform 1 0 9108 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_99
timestamp 1644511149
transform 1 0 10212 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_41_111
timestamp 1644511149
transform 1 0 11316 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_113
timestamp 1644511149
transform 1 0 11500 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_41_125
timestamp 1644511149
transform 1 0 12604 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_135
timestamp 1644511149
transform 1 0 13524 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_147
timestamp 1644511149
transform 1 0 14628 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_153
timestamp 1644511149
transform 1 0 15180 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_157
timestamp 1644511149
transform 1 0 15548 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_41_165
timestamp 1644511149
transform 1 0 16284 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_41_175
timestamp 1644511149
transform 1 0 17204 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_185
timestamp 1644511149
transform 1 0 18124 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_41_196
timestamp 1644511149
transform 1 0 19136 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_220
timestamp 1644511149
transform 1 0 21344 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_41_235
timestamp 1644511149
transform 1 0 22724 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_247
timestamp 1644511149
transform 1 0 23828 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_41_276
timestamp 1644511149
transform 1 0 26496 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_285
timestamp 1644511149
transform 1 0 27324 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_41_292
timestamp 1644511149
transform 1 0 27968 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_298
timestamp 1644511149
transform 1 0 28520 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_24
timestamp 1644511149
transform 1 0 3312 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_42_29
timestamp 1644511149
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_50
timestamp 1644511149
transform 1 0 5704 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_62
timestamp 1644511149
transform 1 0 6808 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_74
timestamp 1644511149
transform 1 0 7912 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_82
timestamp 1644511149
transform 1 0 8648 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_42_85
timestamp 1644511149
transform 1 0 8924 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_97
timestamp 1644511149
transform 1 0 10028 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_109
timestamp 1644511149
transform 1 0 11132 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_42_117
timestamp 1644511149
transform 1 0 11868 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_42_136
timestamp 1644511149
transform 1 0 13616 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_141
timestamp 1644511149
transform 1 0 14076 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_149
timestamp 1644511149
transform 1 0 14812 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_42_155
timestamp 1644511149
transform 1 0 15364 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_42_168
timestamp 1644511149
transform 1 0 16560 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_180
timestamp 1644511149
transform 1 0 17664 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_192
timestamp 1644511149
transform 1 0 18768 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_42_197
timestamp 1644511149
transform 1 0 19228 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_209
timestamp 1644511149
transform 1 0 20332 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_221
timestamp 1644511149
transform 1 0 21436 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_225
timestamp 1644511149
transform 1 0 21804 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_230
timestamp 1644511149
transform 1 0 22264 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_241
timestamp 1644511149
transform 1 0 23276 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_248
timestamp 1644511149
transform 1 0 23920 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_269
timestamp 1644511149
transform 1 0 25852 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_273
timestamp 1644511149
transform 1 0 26220 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_295
timestamp 1644511149
transform 1 0 28244 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_3
timestamp 1644511149
transform 1 0 1380 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_7
timestamp 1644511149
transform 1 0 1748 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_19
timestamp 1644511149
transform 1 0 2852 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_31
timestamp 1644511149
transform 1 0 3956 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_43
timestamp 1644511149
transform 1 0 5060 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_43_55
timestamp 1644511149
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_57
timestamp 1644511149
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_69
timestamp 1644511149
transform 1 0 7452 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_81
timestamp 1644511149
transform 1 0 8556 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_93
timestamp 1644511149
transform 1 0 9660 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_105
timestamp 1644511149
transform 1 0 10764 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_111
timestamp 1644511149
transform 1 0 11316 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_113
timestamp 1644511149
transform 1 0 11500 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_43_121
timestamp 1644511149
transform 1 0 12236 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_43_129
timestamp 1644511149
transform 1 0 12972 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_136
timestamp 1644511149
transform 1 0 13616 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_43_156
timestamp 1644511149
transform 1 0 15456 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_169
timestamp 1644511149
transform 1 0 16652 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_177
timestamp 1644511149
transform 1 0 17388 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_43_186
timestamp 1644511149
transform 1 0 18216 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_194
timestamp 1644511149
transform 1 0 18952 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_198
timestamp 1644511149
transform 1 0 19320 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_210
timestamp 1644511149
transform 1 0 20424 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_43_222
timestamp 1644511149
transform 1 0 21528 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_225
timestamp 1644511149
transform 1 0 21804 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_229
timestamp 1644511149
transform 1 0 22172 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_235
timestamp 1644511149
transform 1 0 22724 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_247
timestamp 1644511149
transform 1 0 23828 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_255
timestamp 1644511149
transform 1 0 24564 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_43_262
timestamp 1644511149
transform 1 0 25208 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_274
timestamp 1644511149
transform 1 0 26312 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_43_281
timestamp 1644511149
transform 1 0 26956 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_43_290
timestamp 1644511149
transform 1 0 27784 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_298
timestamp 1644511149
transform 1 0 28520 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_3
timestamp 1644511149
transform 1 0 1380 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_15
timestamp 1644511149
transform 1 0 2484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_27
timestamp 1644511149
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_29
timestamp 1644511149
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_41
timestamp 1644511149
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_53
timestamp 1644511149
transform 1 0 5980 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_65
timestamp 1644511149
transform 1 0 7084 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_77
timestamp 1644511149
transform 1 0 8188 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_83
timestamp 1644511149
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_85
timestamp 1644511149
transform 1 0 8924 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_97
timestamp 1644511149
transform 1 0 10028 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_109
timestamp 1644511149
transform 1 0 11132 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_121
timestamp 1644511149
transform 1 0 12236 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_133
timestamp 1644511149
transform 1 0 13340 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_139
timestamp 1644511149
transform 1 0 13892 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_141
timestamp 1644511149
transform 1 0 14076 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_145
timestamp 1644511149
transform 1 0 14444 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_44_149
timestamp 1644511149
transform 1 0 14812 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_44_161
timestamp 1644511149
transform 1 0 15916 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_173
timestamp 1644511149
transform 1 0 17020 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_177
timestamp 1644511149
transform 1 0 17388 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_184
timestamp 1644511149
transform 1 0 18032 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_201
timestamp 1644511149
transform 1 0 19596 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_208
timestamp 1644511149
transform 1 0 20240 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_44_216
timestamp 1644511149
transform 1 0 20976 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_44_226
timestamp 1644511149
transform 1 0 21896 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_236
timestamp 1644511149
transform 1 0 22816 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_44_246
timestamp 1644511149
transform 1 0 23736 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_44_269
timestamp 1644511149
transform 1 0 25852 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_44_281
timestamp 1644511149
transform 1 0 26956 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_44_287
timestamp 1644511149
transform 1 0 27508 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_294
timestamp 1644511149
transform 1 0 28152 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_298
timestamp 1644511149
transform 1 0 28520 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_3
timestamp 1644511149
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_15
timestamp 1644511149
transform 1 0 2484 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_27
timestamp 1644511149
transform 1 0 3588 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_39
timestamp 1644511149
transform 1 0 4692 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_51
timestamp 1644511149
transform 1 0 5796 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_55
timestamp 1644511149
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_57
timestamp 1644511149
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_69
timestamp 1644511149
transform 1 0 7452 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_81
timestamp 1644511149
transform 1 0 8556 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_93
timestamp 1644511149
transform 1 0 9660 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_105
timestamp 1644511149
transform 1 0 10764 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_111
timestamp 1644511149
transform 1 0 11316 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_113
timestamp 1644511149
transform 1 0 11500 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_125
timestamp 1644511149
transform 1 0 12604 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_137
timestamp 1644511149
transform 1 0 13708 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_149
timestamp 1644511149
transform 1 0 14812 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_157
timestamp 1644511149
transform 1 0 15548 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_164
timestamp 1644511149
transform 1 0 16192 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_172
timestamp 1644511149
transform 1 0 16928 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_182
timestamp 1644511149
transform 1 0 17848 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_189
timestamp 1644511149
transform 1 0 18492 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_209
timestamp 1644511149
transform 1 0 20332 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_45_217
timestamp 1644511149
transform 1 0 21068 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_223
timestamp 1644511149
transform 1 0 21620 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_45_229
timestamp 1644511149
transform 1 0 22172 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_45_238
timestamp 1644511149
transform 1 0 23000 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_250
timestamp 1644511149
transform 1 0 24104 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_262
timestamp 1644511149
transform 1 0 25208 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_274
timestamp 1644511149
transform 1 0 26312 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_45_281
timestamp 1644511149
transform 1 0 26956 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_287
timestamp 1644511149
transform 1 0 27508 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_291
timestamp 1644511149
transform 1 0 27876 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_46_3
timestamp 1644511149
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_15
timestamp 1644511149
transform 1 0 2484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_27
timestamp 1644511149
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_29
timestamp 1644511149
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_41
timestamp 1644511149
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_53
timestamp 1644511149
transform 1 0 5980 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_65
timestamp 1644511149
transform 1 0 7084 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_77
timestamp 1644511149
transform 1 0 8188 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_83
timestamp 1644511149
transform 1 0 8740 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_85
timestamp 1644511149
transform 1 0 8924 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_97
timestamp 1644511149
transform 1 0 10028 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_109
timestamp 1644511149
transform 1 0 11132 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_121
timestamp 1644511149
transform 1 0 12236 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_136
timestamp 1644511149
transform 1 0 13616 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_141
timestamp 1644511149
transform 1 0 14076 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_46_151
timestamp 1644511149
transform 1 0 14996 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_157
timestamp 1644511149
transform 1 0 15548 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_174
timestamp 1644511149
transform 1 0 17112 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_188
timestamp 1644511149
transform 1 0 18400 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_46_197
timestamp 1644511149
transform 1 0 19228 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_204
timestamp 1644511149
transform 1 0 19872 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_215
timestamp 1644511149
transform 1 0 20884 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_224
timestamp 1644511149
transform 1 0 21712 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_46_232
timestamp 1644511149
transform 1 0 22448 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_46_244
timestamp 1644511149
transform 1 0 23552 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_46_253
timestamp 1644511149
transform 1 0 24380 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_265
timestamp 1644511149
transform 1 0 25484 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_273
timestamp 1644511149
transform 1 0 26220 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_295
timestamp 1644511149
transform 1 0 28244 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_47_6
timestamp 1644511149
transform 1 0 1656 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_18
timestamp 1644511149
transform 1 0 2760 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_30
timestamp 1644511149
transform 1 0 3864 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_42
timestamp 1644511149
transform 1 0 4968 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_47_54
timestamp 1644511149
transform 1 0 6072 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_47_57
timestamp 1644511149
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_69
timestamp 1644511149
transform 1 0 7452 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_81
timestamp 1644511149
transform 1 0 8556 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_93
timestamp 1644511149
transform 1 0 9660 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_105
timestamp 1644511149
transform 1 0 10764 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_111
timestamp 1644511149
transform 1 0 11316 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_113
timestamp 1644511149
transform 1 0 11500 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_125
timestamp 1644511149
transform 1 0 12604 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_47_149
timestamp 1644511149
transform 1 0 14812 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_47_157
timestamp 1644511149
transform 1 0 15548 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_164
timestamp 1644511149
transform 1 0 16192 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_172
timestamp 1644511149
transform 1 0 16928 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_176
timestamp 1644511149
transform 1 0 17296 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_183
timestamp 1644511149
transform 1 0 17940 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_193
timestamp 1644511149
transform 1 0 18860 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_203
timestamp 1644511149
transform 1 0 19780 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_47_215
timestamp 1644511149
transform 1 0 20884 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_223
timestamp 1644511149
transform 1 0 21620 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_47_225
timestamp 1644511149
transform 1 0 21804 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_47_232
timestamp 1644511149
transform 1 0 22448 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_47_246
timestamp 1644511149
transform 1 0 23736 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_47_266
timestamp 1644511149
transform 1 0 25576 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_47_278
timestamp 1644511149
transform 1 0 26680 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_47_281
timestamp 1644511149
transform 1 0 26956 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_47_287
timestamp 1644511149
transform 1 0 27508 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_294
timestamp 1644511149
transform 1 0 28152 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_298
timestamp 1644511149
transform 1 0 28520 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_3
timestamp 1644511149
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_15
timestamp 1644511149
transform 1 0 2484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 1644511149
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_29
timestamp 1644511149
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_41
timestamp 1644511149
transform 1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_53
timestamp 1644511149
transform 1 0 5980 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_65
timestamp 1644511149
transform 1 0 7084 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_77
timestamp 1644511149
transform 1 0 8188 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_83
timestamp 1644511149
transform 1 0 8740 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_85
timestamp 1644511149
transform 1 0 8924 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_97
timestamp 1644511149
transform 1 0 10028 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_109
timestamp 1644511149
transform 1 0 11132 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_121
timestamp 1644511149
transform 1 0 12236 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_133
timestamp 1644511149
transform 1 0 13340 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_139
timestamp 1644511149
transform 1 0 13892 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_48_141
timestamp 1644511149
transform 1 0 14076 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_147
timestamp 1644511149
transform 1 0 14628 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_159
timestamp 1644511149
transform 1 0 15732 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_171
timestamp 1644511149
transform 1 0 16836 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_175
timestamp 1644511149
transform 1 0 17204 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_182
timestamp 1644511149
transform 1 0 17848 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_48_194
timestamp 1644511149
transform 1 0 18952 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_48_197
timestamp 1644511149
transform 1 0 19228 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_209
timestamp 1644511149
transform 1 0 20332 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_48_221
timestamp 1644511149
transform 1 0 21436 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_227
timestamp 1644511149
transform 1 0 21988 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_231
timestamp 1644511149
transform 1 0 22356 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_235
timestamp 1644511149
transform 1 0 22724 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_48_245
timestamp 1644511149
transform 1 0 23644 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_251
timestamp 1644511149
transform 1 0 24196 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_253
timestamp 1644511149
transform 1 0 24380 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_265
timestamp 1644511149
transform 1 0 25484 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_273
timestamp 1644511149
transform 1 0 26220 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_295
timestamp 1644511149
transform 1 0 28244 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_49_3
timestamp 1644511149
transform 1 0 1380 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_15
timestamp 1644511149
transform 1 0 2484 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_27
timestamp 1644511149
transform 1 0 3588 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_39
timestamp 1644511149
transform 1 0 4692 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_51
timestamp 1644511149
transform 1 0 5796 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_55
timestamp 1644511149
transform 1 0 6164 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_57
timestamp 1644511149
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_69
timestamp 1644511149
transform 1 0 7452 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_81
timestamp 1644511149
transform 1 0 8556 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_93
timestamp 1644511149
transform 1 0 9660 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_105
timestamp 1644511149
transform 1 0 10764 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_111
timestamp 1644511149
transform 1 0 11316 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_113
timestamp 1644511149
transform 1 0 11500 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_125
timestamp 1644511149
transform 1 0 12604 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_137
timestamp 1644511149
transform 1 0 13708 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_149
timestamp 1644511149
transform 1 0 14812 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_161
timestamp 1644511149
transform 1 0 15916 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_167
timestamp 1644511149
transform 1 0 16468 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_169
timestamp 1644511149
transform 1 0 16652 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_181
timestamp 1644511149
transform 1 0 17756 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_193
timestamp 1644511149
transform 1 0 18860 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_205
timestamp 1644511149
transform 1 0 19964 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_217
timestamp 1644511149
transform 1 0 21068 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_223
timestamp 1644511149
transform 1 0 21620 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_225
timestamp 1644511149
transform 1 0 21804 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_237
timestamp 1644511149
transform 1 0 22908 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_249
timestamp 1644511149
transform 1 0 24012 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_261
timestamp 1644511149
transform 1 0 25116 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_273
timestamp 1644511149
transform 1 0 26220 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_279
timestamp 1644511149
transform 1 0 26772 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_49_281
timestamp 1644511149
transform 1 0 26956 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_286
timestamp 1644511149
transform 1 0 27416 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_49_293
timestamp 1644511149
transform 1 0 28060 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_50_3
timestamp 1644511149
transform 1 0 1380 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_15
timestamp 1644511149
transform 1 0 2484 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_27
timestamp 1644511149
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_29
timestamp 1644511149
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_41
timestamp 1644511149
transform 1 0 4876 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_53
timestamp 1644511149
transform 1 0 5980 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_65
timestamp 1644511149
transform 1 0 7084 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_77
timestamp 1644511149
transform 1 0 8188 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_83
timestamp 1644511149
transform 1 0 8740 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_85
timestamp 1644511149
transform 1 0 8924 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_97
timestamp 1644511149
transform 1 0 10028 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_109
timestamp 1644511149
transform 1 0 11132 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_121
timestamp 1644511149
transform 1 0 12236 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_133
timestamp 1644511149
transform 1 0 13340 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_139
timestamp 1644511149
transform 1 0 13892 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_50_141
timestamp 1644511149
transform 1 0 14076 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_147
timestamp 1644511149
transform 1 0 14628 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_157
timestamp 1644511149
transform 1 0 15548 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_50_165
timestamp 1644511149
transform 1 0 16284 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_50_187
timestamp 1644511149
transform 1 0 18308 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_195
timestamp 1644511149
transform 1 0 19044 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_50_213
timestamp 1644511149
transform 1 0 20700 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_221
timestamp 1644511149
transform 1 0 21436 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_229
timestamp 1644511149
transform 1 0 22172 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_236
timestamp 1644511149
transform 1 0 22816 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_248
timestamp 1644511149
transform 1 0 23920 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_269
timestamp 1644511149
transform 1 0 25852 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_273
timestamp 1644511149
transform 1 0 26220 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_295
timestamp 1644511149
transform 1 0 28244 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_51_6
timestamp 1644511149
transform 1 0 1656 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_18
timestamp 1644511149
transform 1 0 2760 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_30
timestamp 1644511149
transform 1 0 3864 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_42
timestamp 1644511149
transform 1 0 4968 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_51_54
timestamp 1644511149
transform 1 0 6072 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_51_57
timestamp 1644511149
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_69
timestamp 1644511149
transform 1 0 7452 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_81
timestamp 1644511149
transform 1 0 8556 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_93
timestamp 1644511149
transform 1 0 9660 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_105
timestamp 1644511149
transform 1 0 10764 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_111
timestamp 1644511149
transform 1 0 11316 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_113
timestamp 1644511149
transform 1 0 11500 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_125
timestamp 1644511149
transform 1 0 12604 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_137
timestamp 1644511149
transform 1 0 13708 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_51_145
timestamp 1644511149
transform 1 0 14444 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_164
timestamp 1644511149
transform 1 0 16192 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_172
timestamp 1644511149
transform 1 0 16928 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_51_185
timestamp 1644511149
transform 1 0 18124 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_193
timestamp 1644511149
transform 1 0 18860 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_198
timestamp 1644511149
transform 1 0 19320 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_206
timestamp 1644511149
transform 1 0 20056 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_51_218
timestamp 1644511149
transform 1 0 21160 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_51_233
timestamp 1644511149
transform 1 0 22540 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_51_241
timestamp 1644511149
transform 1 0 23276 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_253
timestamp 1644511149
transform 1 0 24380 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_257
timestamp 1644511149
transform 1 0 24748 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_275
timestamp 1644511149
transform 1 0 26404 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_279
timestamp 1644511149
transform 1 0 26772 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_51_284
timestamp 1644511149
transform 1 0 27232 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_51_293
timestamp 1644511149
transform 1 0 28060 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_52_3
timestamp 1644511149
transform 1 0 1380 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_15
timestamp 1644511149
transform 1 0 2484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_27
timestamp 1644511149
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_29
timestamp 1644511149
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_41
timestamp 1644511149
transform 1 0 4876 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_53
timestamp 1644511149
transform 1 0 5980 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_65
timestamp 1644511149
transform 1 0 7084 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_77
timestamp 1644511149
transform 1 0 8188 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_83
timestamp 1644511149
transform 1 0 8740 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_85
timestamp 1644511149
transform 1 0 8924 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_97
timestamp 1644511149
transform 1 0 10028 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_109
timestamp 1644511149
transform 1 0 11132 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_121
timestamp 1644511149
transform 1 0 12236 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_133
timestamp 1644511149
transform 1 0 13340 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_139
timestamp 1644511149
transform 1 0 13892 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_52_141
timestamp 1644511149
transform 1 0 14076 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_52_152
timestamp 1644511149
transform 1 0 15088 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_52_159
timestamp 1644511149
transform 1 0 15732 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_171
timestamp 1644511149
transform 1 0 16836 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_177
timestamp 1644511149
transform 1 0 17388 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_189
timestamp 1644511149
transform 1 0 18492 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_195
timestamp 1644511149
transform 1 0 19044 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_52_201
timestamp 1644511149
transform 1 0 19596 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_52_211
timestamp 1644511149
transform 1 0 20516 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_220
timestamp 1644511149
transform 1 0 21344 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_52_228
timestamp 1644511149
transform 1 0 22080 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_240
timestamp 1644511149
transform 1 0 23184 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_253
timestamp 1644511149
transform 1 0 24380 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_52_262
timestamp 1644511149
transform 1 0 25208 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_295
timestamp 1644511149
transform 1 0 28244 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_3
timestamp 1644511149
transform 1 0 1380 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_53_10
timestamp 1644511149
transform 1 0 2024 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_22
timestamp 1644511149
transform 1 0 3128 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_34
timestamp 1644511149
transform 1 0 4232 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_46
timestamp 1644511149
transform 1 0 5336 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_54
timestamp 1644511149
transform 1 0 6072 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_53_57
timestamp 1644511149
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_69
timestamp 1644511149
transform 1 0 7452 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_81
timestamp 1644511149
transform 1 0 8556 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_93
timestamp 1644511149
transform 1 0 9660 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_105
timestamp 1644511149
transform 1 0 10764 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_111
timestamp 1644511149
transform 1 0 11316 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_113
timestamp 1644511149
transform 1 0 11500 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_125
timestamp 1644511149
transform 1 0 12604 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_137
timestamp 1644511149
transform 1 0 13708 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_149
timestamp 1644511149
transform 1 0 14812 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_161
timestamp 1644511149
transform 1 0 15916 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_167
timestamp 1644511149
transform 1 0 16468 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_53_169
timestamp 1644511149
transform 1 0 16652 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_53_176
timestamp 1644511149
transform 1 0 17296 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_184
timestamp 1644511149
transform 1 0 18032 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_53_202
timestamp 1644511149
transform 1 0 19688 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_214
timestamp 1644511149
transform 1 0 20792 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_222
timestamp 1644511149
transform 1 0 21528 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_228
timestamp 1644511149
transform 1 0 22080 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_232
timestamp 1644511149
transform 1 0 22448 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_249
timestamp 1644511149
transform 1 0 24012 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_261
timestamp 1644511149
transform 1 0 25116 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_273
timestamp 1644511149
transform 1 0 26220 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_279
timestamp 1644511149
transform 1 0 26772 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_53_281
timestamp 1644511149
transform 1 0 26956 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_53_289
timestamp 1644511149
transform 1 0 27692 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_53_293
timestamp 1644511149
transform 1 0 28060 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_54_24
timestamp 1644511149
transform 1 0 3312 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_54_29
timestamp 1644511149
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_41
timestamp 1644511149
transform 1 0 4876 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_53
timestamp 1644511149
transform 1 0 5980 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_65
timestamp 1644511149
transform 1 0 7084 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_77
timestamp 1644511149
transform 1 0 8188 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_83
timestamp 1644511149
transform 1 0 8740 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_85
timestamp 1644511149
transform 1 0 8924 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_97
timestamp 1644511149
transform 1 0 10028 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_109
timestamp 1644511149
transform 1 0 11132 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_121
timestamp 1644511149
transform 1 0 12236 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_133
timestamp 1644511149
transform 1 0 13340 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_139
timestamp 1644511149
transform 1 0 13892 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_141
timestamp 1644511149
transform 1 0 14076 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_153
timestamp 1644511149
transform 1 0 15180 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_54_165
timestamp 1644511149
transform 1 0 16284 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_170
timestamp 1644511149
transform 1 0 16744 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_54_183
timestamp 1644511149
transform 1 0 17940 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_54_192
timestamp 1644511149
transform 1 0 18768 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_202
timestamp 1644511149
transform 1 0 19688 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_54_209
timestamp 1644511149
transform 1 0 20332 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_54_221
timestamp 1644511149
transform 1 0 21436 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_225
timestamp 1644511149
transform 1 0 21804 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_54_233
timestamp 1644511149
transform 1 0 22540 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_54_241
timestamp 1644511149
transform 1 0 23276 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_54_246
timestamp 1644511149
transform 1 0 23736 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_54_253
timestamp 1644511149
transform 1 0 24380 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_265
timestamp 1644511149
transform 1 0 25484 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_287
timestamp 1644511149
transform 1 0 27508 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_294
timestamp 1644511149
transform 1 0 28152 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_298
timestamp 1644511149
transform 1 0 28520 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_55_3
timestamp 1644511149
transform 1 0 1380 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_7
timestamp 1644511149
transform 1 0 1748 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_19
timestamp 1644511149
transform 1 0 2852 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_31
timestamp 1644511149
transform 1 0 3956 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_43
timestamp 1644511149
transform 1 0 5060 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_55_55
timestamp 1644511149
transform 1 0 6164 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_57
timestamp 1644511149
transform 1 0 6348 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_69
timestamp 1644511149
transform 1 0 7452 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_81
timestamp 1644511149
transform 1 0 8556 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_93
timestamp 1644511149
transform 1 0 9660 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_105
timestamp 1644511149
transform 1 0 10764 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_111
timestamp 1644511149
transform 1 0 11316 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_113
timestamp 1644511149
transform 1 0 11500 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_125
timestamp 1644511149
transform 1 0 12604 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_137
timestamp 1644511149
transform 1 0 13708 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_149
timestamp 1644511149
transform 1 0 14812 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_161
timestamp 1644511149
transform 1 0 15916 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_167
timestamp 1644511149
transform 1 0 16468 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_185
timestamp 1644511149
transform 1 0 18124 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_197
timestamp 1644511149
transform 1 0 19228 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_55_210
timestamp 1644511149
transform 1 0 20424 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_219
timestamp 1644511149
transform 1 0 21252 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_223
timestamp 1644511149
transform 1 0 21620 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_232
timestamp 1644511149
transform 1 0 22448 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_244
timestamp 1644511149
transform 1 0 23552 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_55_252
timestamp 1644511149
transform 1 0 24288 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_55_276
timestamp 1644511149
transform 1 0 26496 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_284
timestamp 1644511149
transform 1 0 27232 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_288
timestamp 1644511149
transform 1 0 27600 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_55_292
timestamp 1644511149
transform 1 0 27968 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_298
timestamp 1644511149
transform 1 0 28520 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_3
timestamp 1644511149
transform 1 0 1380 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_15
timestamp 1644511149
transform 1 0 2484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_27
timestamp 1644511149
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_29
timestamp 1644511149
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_41
timestamp 1644511149
transform 1 0 4876 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_53
timestamp 1644511149
transform 1 0 5980 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_65
timestamp 1644511149
transform 1 0 7084 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_77
timestamp 1644511149
transform 1 0 8188 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_83
timestamp 1644511149
transform 1 0 8740 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_85
timestamp 1644511149
transform 1 0 8924 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_97
timestamp 1644511149
transform 1 0 10028 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_109
timestamp 1644511149
transform 1 0 11132 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_121
timestamp 1644511149
transform 1 0 12236 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_133
timestamp 1644511149
transform 1 0 13340 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_139
timestamp 1644511149
transform 1 0 13892 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_141
timestamp 1644511149
transform 1 0 14076 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_153
timestamp 1644511149
transform 1 0 15180 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_165
timestamp 1644511149
transform 1 0 16284 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_177
timestamp 1644511149
transform 1 0 17388 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_189
timestamp 1644511149
transform 1 0 18492 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_195
timestamp 1644511149
transform 1 0 19044 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_197
timestamp 1644511149
transform 1 0 19228 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_201
timestamp 1644511149
transform 1 0 19596 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_210
timestamp 1644511149
transform 1 0 20424 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_222
timestamp 1644511149
transform 1 0 21528 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_56_230
timestamp 1644511149
transform 1 0 22264 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_239
timestamp 1644511149
transform 1 0 23092 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_247
timestamp 1644511149
transform 1 0 23828 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_251
timestamp 1644511149
transform 1 0 24196 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_253
timestamp 1644511149
transform 1 0 24380 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_56_265
timestamp 1644511149
transform 1 0 25484 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_56_270
timestamp 1644511149
transform 1 0 25944 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_295
timestamp 1644511149
transform 1 0 28244 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_57_3
timestamp 1644511149
transform 1 0 1380 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_15
timestamp 1644511149
transform 1 0 2484 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_27
timestamp 1644511149
transform 1 0 3588 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_39
timestamp 1644511149
transform 1 0 4692 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_51
timestamp 1644511149
transform 1 0 5796 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_55
timestamp 1644511149
transform 1 0 6164 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_57
timestamp 1644511149
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_69
timestamp 1644511149
transform 1 0 7452 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_81
timestamp 1644511149
transform 1 0 8556 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_93
timestamp 1644511149
transform 1 0 9660 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_105
timestamp 1644511149
transform 1 0 10764 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_111
timestamp 1644511149
transform 1 0 11316 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_113
timestamp 1644511149
transform 1 0 11500 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_125
timestamp 1644511149
transform 1 0 12604 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_137
timestamp 1644511149
transform 1 0 13708 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_149
timestamp 1644511149
transform 1 0 14812 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_161
timestamp 1644511149
transform 1 0 15916 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_167
timestamp 1644511149
transform 1 0 16468 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_169
timestamp 1644511149
transform 1 0 16652 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_57_181
timestamp 1644511149
transform 1 0 17756 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_199
timestamp 1644511149
transform 1 0 19412 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_57_210
timestamp 1644511149
transform 1 0 20424 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_57_222
timestamp 1644511149
transform 1 0 21528 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_57_225
timestamp 1644511149
transform 1 0 21804 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_231
timestamp 1644511149
transform 1 0 22356 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_236
timestamp 1644511149
transform 1 0 22816 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_57_256
timestamp 1644511149
transform 1 0 24656 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_57_264
timestamp 1644511149
transform 1 0 25392 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_269
timestamp 1644511149
transform 1 0 25852 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_276
timestamp 1644511149
transform 1 0 26496 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_281
timestamp 1644511149
transform 1 0 26956 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_285
timestamp 1644511149
transform 1 0 27324 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_295
timestamp 1644511149
transform 1 0 28244 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_58_3
timestamp 1644511149
transform 1 0 1380 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_18
timestamp 1644511149
transform 1 0 2760 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_58_26
timestamp 1644511149
transform 1 0 3496 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_58_29
timestamp 1644511149
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_41
timestamp 1644511149
transform 1 0 4876 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_53
timestamp 1644511149
transform 1 0 5980 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_65
timestamp 1644511149
transform 1 0 7084 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_77
timestamp 1644511149
transform 1 0 8188 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_83
timestamp 1644511149
transform 1 0 8740 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_85
timestamp 1644511149
transform 1 0 8924 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_97
timestamp 1644511149
transform 1 0 10028 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_109
timestamp 1644511149
transform 1 0 11132 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_121
timestamp 1644511149
transform 1 0 12236 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_133
timestamp 1644511149
transform 1 0 13340 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_139
timestamp 1644511149
transform 1 0 13892 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_141
timestamp 1644511149
transform 1 0 14076 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_153
timestamp 1644511149
transform 1 0 15180 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_165
timestamp 1644511149
transform 1 0 16284 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_177
timestamp 1644511149
transform 1 0 17388 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_189
timestamp 1644511149
transform 1 0 18492 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_195
timestamp 1644511149
transform 1 0 19044 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_58_200
timestamp 1644511149
transform 1 0 19504 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_206
timestamp 1644511149
transform 1 0 20056 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_214
timestamp 1644511149
transform 1 0 20792 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_218
timestamp 1644511149
transform 1 0 21160 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_223
timestamp 1644511149
transform 1 0 21620 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_235
timestamp 1644511149
transform 1 0 22724 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_58_248
timestamp 1644511149
transform 1 0 23920 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_257
timestamp 1644511149
transform 1 0 24748 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_269
timestamp 1644511149
transform 1 0 25852 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_273
timestamp 1644511149
transform 1 0 26220 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_295
timestamp 1644511149
transform 1 0 28244 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_3
timestamp 1644511149
transform 1 0 1380 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_59_28
timestamp 1644511149
transform 1 0 3680 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_40
timestamp 1644511149
transform 1 0 4784 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_52
timestamp 1644511149
transform 1 0 5888 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_59_57
timestamp 1644511149
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_69
timestamp 1644511149
transform 1 0 7452 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_81
timestamp 1644511149
transform 1 0 8556 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_93
timestamp 1644511149
transform 1 0 9660 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_105
timestamp 1644511149
transform 1 0 10764 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_111
timestamp 1644511149
transform 1 0 11316 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_113
timestamp 1644511149
transform 1 0 11500 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_125
timestamp 1644511149
transform 1 0 12604 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_137
timestamp 1644511149
transform 1 0 13708 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_149
timestamp 1644511149
transform 1 0 14812 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_161
timestamp 1644511149
transform 1 0 15916 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_167
timestamp 1644511149
transform 1 0 16468 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_169
timestamp 1644511149
transform 1 0 16652 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_59_181
timestamp 1644511149
transform 1 0 17756 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_59_192
timestamp 1644511149
transform 1 0 18768 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_204
timestamp 1644511149
transform 1 0 19872 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_59_220
timestamp 1644511149
transform 1 0 21344 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_59_230
timestamp 1644511149
transform 1 0 22264 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_242
timestamp 1644511149
transform 1 0 23368 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_254
timestamp 1644511149
transform 1 0 24472 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_59_276
timestamp 1644511149
transform 1 0 26496 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_59_290
timestamp 1644511149
transform 1 0 27784 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_59_298
timestamp 1644511149
transform 1 0 28520 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_24
timestamp 1644511149
transform 1 0 3312 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_60_29
timestamp 1644511149
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_41
timestamp 1644511149
transform 1 0 4876 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_53
timestamp 1644511149
transform 1 0 5980 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_65
timestamp 1644511149
transform 1 0 7084 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_77
timestamp 1644511149
transform 1 0 8188 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_83
timestamp 1644511149
transform 1 0 8740 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_85
timestamp 1644511149
transform 1 0 8924 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_97
timestamp 1644511149
transform 1 0 10028 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_109
timestamp 1644511149
transform 1 0 11132 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_121
timestamp 1644511149
transform 1 0 12236 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_133
timestamp 1644511149
transform 1 0 13340 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_139
timestamp 1644511149
transform 1 0 13892 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_141
timestamp 1644511149
transform 1 0 14076 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_153
timestamp 1644511149
transform 1 0 15180 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_165
timestamp 1644511149
transform 1 0 16284 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_177
timestamp 1644511149
transform 1 0 17388 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_60_192
timestamp 1644511149
transform 1 0 18768 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_197
timestamp 1644511149
transform 1 0 19228 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_204
timestamp 1644511149
transform 1 0 19872 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_213
timestamp 1644511149
transform 1 0 20700 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_60_222
timestamp 1644511149
transform 1 0 21528 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_60_230
timestamp 1644511149
transform 1 0 22264 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_60_240
timestamp 1644511149
transform 1 0 23184 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_60_253
timestamp 1644511149
transform 1 0 24380 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_60_265
timestamp 1644511149
transform 1 0 25484 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_285
timestamp 1644511149
transform 1 0 27324 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_295
timestamp 1644511149
transform 1 0 28244 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_3
timestamp 1644511149
transform 1 0 1380 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_7
timestamp 1644511149
transform 1 0 1748 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_61_14
timestamp 1644511149
transform 1 0 2392 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_26
timestamp 1644511149
transform 1 0 3496 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_38
timestamp 1644511149
transform 1 0 4600 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_50
timestamp 1644511149
transform 1 0 5704 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_61_57
timestamp 1644511149
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_69
timestamp 1644511149
transform 1 0 7452 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_81
timestamp 1644511149
transform 1 0 8556 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_93
timestamp 1644511149
transform 1 0 9660 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_105
timestamp 1644511149
transform 1 0 10764 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_111
timestamp 1644511149
transform 1 0 11316 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_113
timestamp 1644511149
transform 1 0 11500 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_125
timestamp 1644511149
transform 1 0 12604 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_137
timestamp 1644511149
transform 1 0 13708 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_149
timestamp 1644511149
transform 1 0 14812 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_161
timestamp 1644511149
transform 1 0 15916 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_167
timestamp 1644511149
transform 1 0 16468 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_61_169
timestamp 1644511149
transform 1 0 16652 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_61_175
timestamp 1644511149
transform 1 0 17204 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_188
timestamp 1644511149
transform 1 0 18400 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_61_208
timestamp 1644511149
transform 1 0 20240 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_61_220
timestamp 1644511149
transform 1 0 21344 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_225
timestamp 1644511149
transform 1 0 21804 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_229
timestamp 1644511149
transform 1 0 22172 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_237
timestamp 1644511149
transform 1 0 22908 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_61_257
timestamp 1644511149
transform 1 0 24748 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_263
timestamp 1644511149
transform 1 0 25300 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_276
timestamp 1644511149
transform 1 0 26496 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_61_289
timestamp 1644511149
transform 1 0 27692 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_61_297
timestamp 1644511149
transform 1 0 28428 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_62_3
timestamp 1644511149
transform 1 0 1380 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_15
timestamp 1644511149
transform 1 0 2484 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_27
timestamp 1644511149
transform 1 0 3588 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_29
timestamp 1644511149
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_41
timestamp 1644511149
transform 1 0 4876 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_53
timestamp 1644511149
transform 1 0 5980 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_65
timestamp 1644511149
transform 1 0 7084 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_77
timestamp 1644511149
transform 1 0 8188 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_83
timestamp 1644511149
transform 1 0 8740 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_85
timestamp 1644511149
transform 1 0 8924 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_97
timestamp 1644511149
transform 1 0 10028 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_109
timestamp 1644511149
transform 1 0 11132 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_121
timestamp 1644511149
transform 1 0 12236 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_133
timestamp 1644511149
transform 1 0 13340 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_139
timestamp 1644511149
transform 1 0 13892 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_141
timestamp 1644511149
transform 1 0 14076 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_153
timestamp 1644511149
transform 1 0 15180 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_165
timestamp 1644511149
transform 1 0 16284 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_177
timestamp 1644511149
transform 1 0 17388 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_62_192
timestamp 1644511149
transform 1 0 18768 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_62_197
timestamp 1644511149
transform 1 0 19228 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_62_205
timestamp 1644511149
transform 1 0 19964 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_210
timestamp 1644511149
transform 1 0 20424 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_62_218
timestamp 1644511149
transform 1 0 21160 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_62_226
timestamp 1644511149
transform 1 0 21896 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_230
timestamp 1644511149
transform 1 0 22264 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_62_242
timestamp 1644511149
transform 1 0 23368 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_62_250
timestamp 1644511149
transform 1 0 24104 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_62_253
timestamp 1644511149
transform 1 0 24380 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_62_265
timestamp 1644511149
transform 1 0 25484 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_62_273
timestamp 1644511149
transform 1 0 26220 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_295
timestamp 1644511149
transform 1 0 28244 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_3
timestamp 1644511149
transform 1 0 1380 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_13
timestamp 1644511149
transform 1 0 2300 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_63_20
timestamp 1644511149
transform 1 0 2944 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_32
timestamp 1644511149
transform 1 0 4048 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_44
timestamp 1644511149
transform 1 0 5152 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_57
timestamp 1644511149
transform 1 0 6348 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_69
timestamp 1644511149
transform 1 0 7452 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_81
timestamp 1644511149
transform 1 0 8556 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_93
timestamp 1644511149
transform 1 0 9660 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_105
timestamp 1644511149
transform 1 0 10764 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_111
timestamp 1644511149
transform 1 0 11316 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_113
timestamp 1644511149
transform 1 0 11500 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_125
timestamp 1644511149
transform 1 0 12604 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_137
timestamp 1644511149
transform 1 0 13708 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_149
timestamp 1644511149
transform 1 0 14812 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_161
timestamp 1644511149
transform 1 0 15916 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_167
timestamp 1644511149
transform 1 0 16468 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_169
timestamp 1644511149
transform 1 0 16652 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_63_181
timestamp 1644511149
transform 1 0 17756 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_63_189
timestamp 1644511149
transform 1 0 18492 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_201
timestamp 1644511149
transform 1 0 19596 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_213
timestamp 1644511149
transform 1 0 20700 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_63_221
timestamp 1644511149
transform 1 0 21436 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_63_225
timestamp 1644511149
transform 1 0 21804 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_231
timestamp 1644511149
transform 1 0 22356 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_236
timestamp 1644511149
transform 1 0 22816 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_248
timestamp 1644511149
transform 1 0 23920 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_260
timestamp 1644511149
transform 1 0 25024 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_272
timestamp 1644511149
transform 1 0 26128 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_63_281
timestamp 1644511149
transform 1 0 26956 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_289
timestamp 1644511149
transform 1 0 27692 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_63_293
timestamp 1644511149
transform 1 0 28060 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_64_24
timestamp 1644511149
transform 1 0 3312 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_64_29
timestamp 1644511149
transform 1 0 3772 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_41
timestamp 1644511149
transform 1 0 4876 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_53
timestamp 1644511149
transform 1 0 5980 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_65
timestamp 1644511149
transform 1 0 7084 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_77
timestamp 1644511149
transform 1 0 8188 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_83
timestamp 1644511149
transform 1 0 8740 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_85
timestamp 1644511149
transform 1 0 8924 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_97
timestamp 1644511149
transform 1 0 10028 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_109
timestamp 1644511149
transform 1 0 11132 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_121
timestamp 1644511149
transform 1 0 12236 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_133
timestamp 1644511149
transform 1 0 13340 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_139
timestamp 1644511149
transform 1 0 13892 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_141
timestamp 1644511149
transform 1 0 14076 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_153
timestamp 1644511149
transform 1 0 15180 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_165
timestamp 1644511149
transform 1 0 16284 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_177
timestamp 1644511149
transform 1 0 17388 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_189
timestamp 1644511149
transform 1 0 18492 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_195
timestamp 1644511149
transform 1 0 19044 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_64_197
timestamp 1644511149
transform 1 0 19228 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_203
timestamp 1644511149
transform 1 0 19780 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_64_208
timestamp 1644511149
transform 1 0 20240 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_214
timestamp 1644511149
transform 1 0 20792 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_221
timestamp 1644511149
transform 1 0 21436 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_64_229
timestamp 1644511149
transform 1 0 22172 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_241
timestamp 1644511149
transform 1 0 23276 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_64_249
timestamp 1644511149
transform 1 0 24012 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_253
timestamp 1644511149
transform 1 0 24380 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_265
timestamp 1644511149
transform 1 0 25484 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_280
timestamp 1644511149
transform 1 0 26864 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_287
timestamp 1644511149
transform 1 0 27508 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_294
timestamp 1644511149
transform 1 0 28152 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_298
timestamp 1644511149
transform 1 0 28520 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_65_6
timestamp 1644511149
transform 1 0 1656 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_65_13
timestamp 1644511149
transform 1 0 2300 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_25
timestamp 1644511149
transform 1 0 3404 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_37
timestamp 1644511149
transform 1 0 4508 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_49
timestamp 1644511149
transform 1 0 5612 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_55
timestamp 1644511149
transform 1 0 6164 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_57
timestamp 1644511149
transform 1 0 6348 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_69
timestamp 1644511149
transform 1 0 7452 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_81
timestamp 1644511149
transform 1 0 8556 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_93
timestamp 1644511149
transform 1 0 9660 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_105
timestamp 1644511149
transform 1 0 10764 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_111
timestamp 1644511149
transform 1 0 11316 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_113
timestamp 1644511149
transform 1 0 11500 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_125
timestamp 1644511149
transform 1 0 12604 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_137
timestamp 1644511149
transform 1 0 13708 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_149
timestamp 1644511149
transform 1 0 14812 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_161
timestamp 1644511149
transform 1 0 15916 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_167
timestamp 1644511149
transform 1 0 16468 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_169
timestamp 1644511149
transform 1 0 16652 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_181
timestamp 1644511149
transform 1 0 17756 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_65_193
timestamp 1644511149
transform 1 0 18860 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_65_201
timestamp 1644511149
transform 1 0 19596 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_65_211
timestamp 1644511149
transform 1 0 20516 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_220
timestamp 1644511149
transform 1 0 21344 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_225
timestamp 1644511149
transform 1 0 21804 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_65_237
timestamp 1644511149
transform 1 0 22908 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_249
timestamp 1644511149
transform 1 0 24012 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_261
timestamp 1644511149
transform 1 0 25116 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_273
timestamp 1644511149
transform 1 0 26220 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_279
timestamp 1644511149
transform 1 0 26772 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_65_281
timestamp 1644511149
transform 1 0 26956 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_287
timestamp 1644511149
transform 1 0 27508 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_65_291
timestamp 1644511149
transform 1 0 27876 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_66_24
timestamp 1644511149
transform 1 0 3312 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_66_29
timestamp 1644511149
transform 1 0 3772 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_41
timestamp 1644511149
transform 1 0 4876 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_53
timestamp 1644511149
transform 1 0 5980 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_65
timestamp 1644511149
transform 1 0 7084 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_77
timestamp 1644511149
transform 1 0 8188 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_83
timestamp 1644511149
transform 1 0 8740 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_85
timestamp 1644511149
transform 1 0 8924 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_97
timestamp 1644511149
transform 1 0 10028 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_109
timestamp 1644511149
transform 1 0 11132 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_121
timestamp 1644511149
transform 1 0 12236 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_133
timestamp 1644511149
transform 1 0 13340 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_139
timestamp 1644511149
transform 1 0 13892 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_141
timestamp 1644511149
transform 1 0 14076 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_153
timestamp 1644511149
transform 1 0 15180 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_165
timestamp 1644511149
transform 1 0 16284 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_177
timestamp 1644511149
transform 1 0 17388 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_189
timestamp 1644511149
transform 1 0 18492 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_195
timestamp 1644511149
transform 1 0 19044 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_66_213
timestamp 1644511149
transform 1 0 20700 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_227
timestamp 1644511149
transform 1 0 21988 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_247
timestamp 1644511149
transform 1 0 23828 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_66_251
timestamp 1644511149
transform 1 0 24196 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_253
timestamp 1644511149
transform 1 0 24380 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_66_265
timestamp 1644511149
transform 1 0 25484 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_66_273
timestamp 1644511149
transform 1 0 26220 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_66_295
timestamp 1644511149
transform 1 0 28244 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_67_3
timestamp 1644511149
transform 1 0 1380 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_67_9
timestamp 1644511149
transform 1 0 1932 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_21
timestamp 1644511149
transform 1 0 3036 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_33
timestamp 1644511149
transform 1 0 4140 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_67_45
timestamp 1644511149
transform 1 0 5244 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_67_53
timestamp 1644511149
transform 1 0 5980 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_67_57
timestamp 1644511149
transform 1 0 6348 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_69
timestamp 1644511149
transform 1 0 7452 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_81
timestamp 1644511149
transform 1 0 8556 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_93
timestamp 1644511149
transform 1 0 9660 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_105
timestamp 1644511149
transform 1 0 10764 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_111
timestamp 1644511149
transform 1 0 11316 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_113
timestamp 1644511149
transform 1 0 11500 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_125
timestamp 1644511149
transform 1 0 12604 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_137
timestamp 1644511149
transform 1 0 13708 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_149
timestamp 1644511149
transform 1 0 14812 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_161
timestamp 1644511149
transform 1 0 15916 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_167
timestamp 1644511149
transform 1 0 16468 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_169
timestamp 1644511149
transform 1 0 16652 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_181
timestamp 1644511149
transform 1 0 17756 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_193
timestamp 1644511149
transform 1 0 18860 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_67_202
timestamp 1644511149
transform 1 0 19688 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_67_216
timestamp 1644511149
transform 1 0 20976 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_67_231
timestamp 1644511149
transform 1 0 22356 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_243
timestamp 1644511149
transform 1 0 23460 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_255
timestamp 1644511149
transform 1 0 24564 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_267
timestamp 1644511149
transform 1 0 25668 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_67_276
timestamp 1644511149
transform 1 0 26496 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_67_281
timestamp 1644511149
transform 1 0 26956 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_67_290
timestamp 1644511149
transform 1 0 27784 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_67_298
timestamp 1644511149
transform 1 0 28520 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_3
timestamp 1644511149
transform 1 0 1380 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_15
timestamp 1644511149
transform 1 0 2484 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_68_27
timestamp 1644511149
transform 1 0 3588 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_29
timestamp 1644511149
transform 1 0 3772 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_41
timestamp 1644511149
transform 1 0 4876 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_53
timestamp 1644511149
transform 1 0 5980 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_65
timestamp 1644511149
transform 1 0 7084 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_77
timestamp 1644511149
transform 1 0 8188 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_83
timestamp 1644511149
transform 1 0 8740 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_85
timestamp 1644511149
transform 1 0 8924 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_97
timestamp 1644511149
transform 1 0 10028 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_109
timestamp 1644511149
transform 1 0 11132 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_121
timestamp 1644511149
transform 1 0 12236 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_133
timestamp 1644511149
transform 1 0 13340 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_139
timestamp 1644511149
transform 1 0 13892 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_141
timestamp 1644511149
transform 1 0 14076 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_153
timestamp 1644511149
transform 1 0 15180 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_165
timestamp 1644511149
transform 1 0 16284 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_177
timestamp 1644511149
transform 1 0 17388 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_189
timestamp 1644511149
transform 1 0 18492 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_195
timestamp 1644511149
transform 1 0 19044 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_197
timestamp 1644511149
transform 1 0 19228 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_68_209
timestamp 1644511149
transform 1 0 20332 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_68_214
timestamp 1644511149
transform 1 0 20792 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_68_222
timestamp 1644511149
transform 1 0 21528 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_234
timestamp 1644511149
transform 1 0 22632 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_246
timestamp 1644511149
transform 1 0 23736 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_68_253
timestamp 1644511149
transform 1 0 24380 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_68_265
timestamp 1644511149
transform 1 0 25484 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_68_273
timestamp 1644511149
transform 1 0 26220 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_68_295
timestamp 1644511149
transform 1 0 28244 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_69_3
timestamp 1644511149
transform 1 0 1380 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_15
timestamp 1644511149
transform 1 0 2484 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_27
timestamp 1644511149
transform 1 0 3588 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_39
timestamp 1644511149
transform 1 0 4692 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_69_51
timestamp 1644511149
transform 1 0 5796 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_55
timestamp 1644511149
transform 1 0 6164 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_57
timestamp 1644511149
transform 1 0 6348 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_69
timestamp 1644511149
transform 1 0 7452 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_81
timestamp 1644511149
transform 1 0 8556 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_93
timestamp 1644511149
transform 1 0 9660 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_105
timestamp 1644511149
transform 1 0 10764 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_111
timestamp 1644511149
transform 1 0 11316 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_113
timestamp 1644511149
transform 1 0 11500 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_125
timestamp 1644511149
transform 1 0 12604 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_137
timestamp 1644511149
transform 1 0 13708 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_149
timestamp 1644511149
transform 1 0 14812 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_161
timestamp 1644511149
transform 1 0 15916 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_167
timestamp 1644511149
transform 1 0 16468 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_169
timestamp 1644511149
transform 1 0 16652 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_181
timestamp 1644511149
transform 1 0 17756 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_193
timestamp 1644511149
transform 1 0 18860 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_205
timestamp 1644511149
transform 1 0 19964 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_217
timestamp 1644511149
transform 1 0 21068 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_223
timestamp 1644511149
transform 1 0 21620 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_225
timestamp 1644511149
transform 1 0 21804 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_237
timestamp 1644511149
transform 1 0 22908 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_249
timestamp 1644511149
transform 1 0 24012 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_261
timestamp 1644511149
transform 1 0 25116 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_273
timestamp 1644511149
transform 1 0 26220 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_279
timestamp 1644511149
transform 1 0 26772 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_69_281
timestamp 1644511149
transform 1 0 26956 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_69_285
timestamp 1644511149
transform 1 0 27324 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_69_292
timestamp 1644511149
transform 1 0 27968 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_298
timestamp 1644511149
transform 1 0 28520 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_70_3
timestamp 1644511149
transform 1 0 1380 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_70_12
timestamp 1644511149
transform 1 0 2208 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_70_19
timestamp 1644511149
transform 1 0 2852 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_70_27
timestamp 1644511149
transform 1 0 3588 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_29
timestamp 1644511149
transform 1 0 3772 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_41
timestamp 1644511149
transform 1 0 4876 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_53
timestamp 1644511149
transform 1 0 5980 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_65
timestamp 1644511149
transform 1 0 7084 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_77
timestamp 1644511149
transform 1 0 8188 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_83
timestamp 1644511149
transform 1 0 8740 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_85
timestamp 1644511149
transform 1 0 8924 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_97
timestamp 1644511149
transform 1 0 10028 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_109
timestamp 1644511149
transform 1 0 11132 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_121
timestamp 1644511149
transform 1 0 12236 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_133
timestamp 1644511149
transform 1 0 13340 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_139
timestamp 1644511149
transform 1 0 13892 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_141
timestamp 1644511149
transform 1 0 14076 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_153
timestamp 1644511149
transform 1 0 15180 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_165
timestamp 1644511149
transform 1 0 16284 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_177
timestamp 1644511149
transform 1 0 17388 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_189
timestamp 1644511149
transform 1 0 18492 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_195
timestamp 1644511149
transform 1 0 19044 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_197
timestamp 1644511149
transform 1 0 19228 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_209
timestamp 1644511149
transform 1 0 20332 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_221
timestamp 1644511149
transform 1 0 21436 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_233
timestamp 1644511149
transform 1 0 22540 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_245
timestamp 1644511149
transform 1 0 23644 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_251
timestamp 1644511149
transform 1 0 24196 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_253
timestamp 1644511149
transform 1 0 24380 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_70_265
timestamp 1644511149
transform 1 0 25484 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_70_273
timestamp 1644511149
transform 1 0 26220 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_70_295
timestamp 1644511149
transform 1 0 28244 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_71_3
timestamp 1644511149
transform 1 0 1380 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_71_26
timestamp 1644511149
transform 1 0 3496 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_38
timestamp 1644511149
transform 1 0 4600 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_50
timestamp 1644511149
transform 1 0 5704 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_71_57
timestamp 1644511149
transform 1 0 6348 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_69
timestamp 1644511149
transform 1 0 7452 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_81
timestamp 1644511149
transform 1 0 8556 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_93
timestamp 1644511149
transform 1 0 9660 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_105
timestamp 1644511149
transform 1 0 10764 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_111
timestamp 1644511149
transform 1 0 11316 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_113
timestamp 1644511149
transform 1 0 11500 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_125
timestamp 1644511149
transform 1 0 12604 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_137
timestamp 1644511149
transform 1 0 13708 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_149
timestamp 1644511149
transform 1 0 14812 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_161
timestamp 1644511149
transform 1 0 15916 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_167
timestamp 1644511149
transform 1 0 16468 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_169
timestamp 1644511149
transform 1 0 16652 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_181
timestamp 1644511149
transform 1 0 17756 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_193
timestamp 1644511149
transform 1 0 18860 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_205
timestamp 1644511149
transform 1 0 19964 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_217
timestamp 1644511149
transform 1 0 21068 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_223
timestamp 1644511149
transform 1 0 21620 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_225
timestamp 1644511149
transform 1 0 21804 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_237
timestamp 1644511149
transform 1 0 22908 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_249
timestamp 1644511149
transform 1 0 24012 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_71_276
timestamp 1644511149
transform 1 0 26496 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_71_284
timestamp 1644511149
transform 1 0 27232 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_290
timestamp 1644511149
transform 1 0 27784 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_71_294
timestamp 1644511149
transform 1 0 28152 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_298
timestamp 1644511149
transform 1 0 28520 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_72_24
timestamp 1644511149
transform 1 0 3312 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_32
timestamp 1644511149
transform 1 0 4048 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_72_39
timestamp 1644511149
transform 1 0 4692 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_51
timestamp 1644511149
transform 1 0 5796 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_63
timestamp 1644511149
transform 1 0 6900 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_72_75
timestamp 1644511149
transform 1 0 8004 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_72_83
timestamp 1644511149
transform 1 0 8740 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_85
timestamp 1644511149
transform 1 0 8924 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_97
timestamp 1644511149
transform 1 0 10028 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_109
timestamp 1644511149
transform 1 0 11132 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_121
timestamp 1644511149
transform 1 0 12236 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_133
timestamp 1644511149
transform 1 0 13340 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_139
timestamp 1644511149
transform 1 0 13892 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_141
timestamp 1644511149
transform 1 0 14076 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_153
timestamp 1644511149
transform 1 0 15180 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_165
timestamp 1644511149
transform 1 0 16284 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_177
timestamp 1644511149
transform 1 0 17388 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_189
timestamp 1644511149
transform 1 0 18492 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_195
timestamp 1644511149
transform 1 0 19044 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_197
timestamp 1644511149
transform 1 0 19228 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_209
timestamp 1644511149
transform 1 0 20332 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_221
timestamp 1644511149
transform 1 0 21436 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_233
timestamp 1644511149
transform 1 0 22540 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_245
timestamp 1644511149
transform 1 0 23644 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_251
timestamp 1644511149
transform 1 0 24196 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_253
timestamp 1644511149
transform 1 0 24380 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_72_265
timestamp 1644511149
transform 1 0 25484 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_72_273
timestamp 1644511149
transform 1 0 26220 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_72_295
timestamp 1644511149
transform 1 0 28244 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_73_3
timestamp 1644511149
transform 1 0 1380 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_73_8
timestamp 1644511149
transform 1 0 1840 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_73_16
timestamp 1644511149
transform 1 0 2576 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_73_39
timestamp 1644511149
transform 1 0 4692 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_73_51
timestamp 1644511149
transform 1 0 5796 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_55
timestamp 1644511149
transform 1 0 6164 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_57
timestamp 1644511149
transform 1 0 6348 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_69
timestamp 1644511149
transform 1 0 7452 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_81
timestamp 1644511149
transform 1 0 8556 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_93
timestamp 1644511149
transform 1 0 9660 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_105
timestamp 1644511149
transform 1 0 10764 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_111
timestamp 1644511149
transform 1 0 11316 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_113
timestamp 1644511149
transform 1 0 11500 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_125
timestamp 1644511149
transform 1 0 12604 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_137
timestamp 1644511149
transform 1 0 13708 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_149
timestamp 1644511149
transform 1 0 14812 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_161
timestamp 1644511149
transform 1 0 15916 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_167
timestamp 1644511149
transform 1 0 16468 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_169
timestamp 1644511149
transform 1 0 16652 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_181
timestamp 1644511149
transform 1 0 17756 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_193
timestamp 1644511149
transform 1 0 18860 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_205
timestamp 1644511149
transform 1 0 19964 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_217
timestamp 1644511149
transform 1 0 21068 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_223
timestamp 1644511149
transform 1 0 21620 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_225
timestamp 1644511149
transform 1 0 21804 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_237
timestamp 1644511149
transform 1 0 22908 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_249
timestamp 1644511149
transform 1 0 24012 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_261
timestamp 1644511149
transform 1 0 25116 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_73_276
timestamp 1644511149
transform 1 0 26496 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_281
timestamp 1644511149
transform 1 0 26956 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_73_285
timestamp 1644511149
transform 1 0 27324 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_73_292
timestamp 1644511149
transform 1 0 27968 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_298
timestamp 1644511149
transform 1 0 28520 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_74_3
timestamp 1644511149
transform 1 0 1380 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_74_8
timestamp 1644511149
transform 1 0 1840 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_74_16
timestamp 1644511149
transform 1 0 2576 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_74_22
timestamp 1644511149
transform 1 0 3128 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_74_29
timestamp 1644511149
transform 1 0 3772 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_41
timestamp 1644511149
transform 1 0 4876 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_53
timestamp 1644511149
transform 1 0 5980 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_65
timestamp 1644511149
transform 1 0 7084 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_77
timestamp 1644511149
transform 1 0 8188 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_83
timestamp 1644511149
transform 1 0 8740 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_85
timestamp 1644511149
transform 1 0 8924 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_97
timestamp 1644511149
transform 1 0 10028 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_109
timestamp 1644511149
transform 1 0 11132 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_121
timestamp 1644511149
transform 1 0 12236 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_133
timestamp 1644511149
transform 1 0 13340 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_139
timestamp 1644511149
transform 1 0 13892 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_141
timestamp 1644511149
transform 1 0 14076 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_153
timestamp 1644511149
transform 1 0 15180 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_165
timestamp 1644511149
transform 1 0 16284 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_177
timestamp 1644511149
transform 1 0 17388 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_189
timestamp 1644511149
transform 1 0 18492 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_195
timestamp 1644511149
transform 1 0 19044 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_197
timestamp 1644511149
transform 1 0 19228 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_209
timestamp 1644511149
transform 1 0 20332 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_221
timestamp 1644511149
transform 1 0 21436 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_233
timestamp 1644511149
transform 1 0 22540 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_245
timestamp 1644511149
transform 1 0 23644 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_251
timestamp 1644511149
transform 1 0 24196 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_253
timestamp 1644511149
transform 1 0 24380 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_74_265
timestamp 1644511149
transform 1 0 25484 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_74_273
timestamp 1644511149
transform 1 0 26220 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_74_295
timestamp 1644511149
transform 1 0 28244 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_75_3
timestamp 1644511149
transform 1 0 1380 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_36
timestamp 1644511149
transform 1 0 4416 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_75_48
timestamp 1644511149
transform 1 0 5520 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_75_57
timestamp 1644511149
transform 1 0 6348 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_69
timestamp 1644511149
transform 1 0 7452 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_81
timestamp 1644511149
transform 1 0 8556 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_93
timestamp 1644511149
transform 1 0 9660 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_105
timestamp 1644511149
transform 1 0 10764 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_111
timestamp 1644511149
transform 1 0 11316 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_113
timestamp 1644511149
transform 1 0 11500 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_125
timestamp 1644511149
transform 1 0 12604 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_137
timestamp 1644511149
transform 1 0 13708 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_149
timestamp 1644511149
transform 1 0 14812 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_161
timestamp 1644511149
transform 1 0 15916 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_167
timestamp 1644511149
transform 1 0 16468 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_169
timestamp 1644511149
transform 1 0 16652 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_181
timestamp 1644511149
transform 1 0 17756 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_193
timestamp 1644511149
transform 1 0 18860 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_205
timestamp 1644511149
transform 1 0 19964 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_217
timestamp 1644511149
transform 1 0 21068 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_223
timestamp 1644511149
transform 1 0 21620 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_225
timestamp 1644511149
transform 1 0 21804 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_237
timestamp 1644511149
transform 1 0 22908 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_249
timestamp 1644511149
transform 1 0 24012 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_261
timestamp 1644511149
transform 1 0 25116 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_273
timestamp 1644511149
transform 1 0 26220 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_279
timestamp 1644511149
transform 1 0 26772 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_75_284
timestamp 1644511149
transform 1 0 27232 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_75_291
timestamp 1644511149
transform 1 0 27876 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_76_24
timestamp 1644511149
transform 1 0 3312 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_76_29
timestamp 1644511149
transform 1 0 3772 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_41
timestamp 1644511149
transform 1 0 4876 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_53
timestamp 1644511149
transform 1 0 5980 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_65
timestamp 1644511149
transform 1 0 7084 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_77
timestamp 1644511149
transform 1 0 8188 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_83
timestamp 1644511149
transform 1 0 8740 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_85
timestamp 1644511149
transform 1 0 8924 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_97
timestamp 1644511149
transform 1 0 10028 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_109
timestamp 1644511149
transform 1 0 11132 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_121
timestamp 1644511149
transform 1 0 12236 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_133
timestamp 1644511149
transform 1 0 13340 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_139
timestamp 1644511149
transform 1 0 13892 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_141
timestamp 1644511149
transform 1 0 14076 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_153
timestamp 1644511149
transform 1 0 15180 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_165
timestamp 1644511149
transform 1 0 16284 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_177
timestamp 1644511149
transform 1 0 17388 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_189
timestamp 1644511149
transform 1 0 18492 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_195
timestamp 1644511149
transform 1 0 19044 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_197
timestamp 1644511149
transform 1 0 19228 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_209
timestamp 1644511149
transform 1 0 20332 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_221
timestamp 1644511149
transform 1 0 21436 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_233
timestamp 1644511149
transform 1 0 22540 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_245
timestamp 1644511149
transform 1 0 23644 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_251
timestamp 1644511149
transform 1 0 24196 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_253
timestamp 1644511149
transform 1 0 24380 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_76_265
timestamp 1644511149
transform 1 0 25484 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_76_270
timestamp 1644511149
transform 1 0 25944 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_295
timestamp 1644511149
transform 1 0 28244 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_3
timestamp 1644511149
transform 1 0 1380 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_77_7
timestamp 1644511149
transform 1 0 1748 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_14
timestamp 1644511149
transform 1 0 2392 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_77_21
timestamp 1644511149
transform 1 0 3036 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_33
timestamp 1644511149
transform 1 0 4140 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_77_45
timestamp 1644511149
transform 1 0 5244 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_77_53
timestamp 1644511149
transform 1 0 5980 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_77_57
timestamp 1644511149
transform 1 0 6348 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_69
timestamp 1644511149
transform 1 0 7452 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_81
timestamp 1644511149
transform 1 0 8556 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_93
timestamp 1644511149
transform 1 0 9660 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_105
timestamp 1644511149
transform 1 0 10764 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_111
timestamp 1644511149
transform 1 0 11316 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_116
timestamp 1644511149
transform 1 0 11776 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_128
timestamp 1644511149
transform 1 0 12880 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_140
timestamp 1644511149
transform 1 0 13984 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_152
timestamp 1644511149
transform 1 0 15088 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_77_164
timestamp 1644511149
transform 1 0 16192 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_77_169
timestamp 1644511149
transform 1 0 16652 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_181
timestamp 1644511149
transform 1 0 17756 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_193
timestamp 1644511149
transform 1 0 18860 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_205
timestamp 1644511149
transform 1 0 19964 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_217
timestamp 1644511149
transform 1 0 21068 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_223
timestamp 1644511149
transform 1 0 21620 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_225
timestamp 1644511149
transform 1 0 21804 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_237
timestamp 1644511149
transform 1 0 22908 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_249
timestamp 1644511149
transform 1 0 24012 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_261
timestamp 1644511149
transform 1 0 25116 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_77_276
timestamp 1644511149
transform 1 0 26496 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_77_281
timestamp 1644511149
transform 1 0 26956 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_77_290
timestamp 1644511149
transform 1 0 27784 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_77_298
timestamp 1644511149
transform 1 0 28520 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_78_3
timestamp 1644511149
transform 1 0 1380 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_78_7
timestamp 1644511149
transform 1 0 1748 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_11
timestamp 1644511149
transform 1 0 2116 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_78_23
timestamp 1644511149
transform 1 0 3220 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_78_27
timestamp 1644511149
transform 1 0 3588 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_29
timestamp 1644511149
transform 1 0 3772 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_41
timestamp 1644511149
transform 1 0 4876 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_53
timestamp 1644511149
transform 1 0 5980 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_65
timestamp 1644511149
transform 1 0 7084 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_77
timestamp 1644511149
transform 1 0 8188 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_83
timestamp 1644511149
transform 1 0 8740 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_85
timestamp 1644511149
transform 1 0 8924 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_78_97
timestamp 1644511149
transform 1 0 10028 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_78_101
timestamp 1644511149
transform 1 0 10396 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_78_105
timestamp 1644511149
transform 1 0 10764 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_78_130
timestamp 1644511149
transform 1 0 13064 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_78_138
timestamp 1644511149
transform 1 0 13800 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_78_141
timestamp 1644511149
transform 1 0 14076 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_153
timestamp 1644511149
transform 1 0 15180 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_165
timestamp 1644511149
transform 1 0 16284 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_177
timestamp 1644511149
transform 1 0 17388 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_189
timestamp 1644511149
transform 1 0 18492 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_195
timestamp 1644511149
transform 1 0 19044 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_78_197
timestamp 1644511149
transform 1 0 19228 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_78_202
timestamp 1644511149
transform 1 0 19688 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_78_206
timestamp 1644511149
transform 1 0 20056 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_210
timestamp 1644511149
transform 1 0 20424 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_222
timestamp 1644511149
transform 1 0 21528 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_237
timestamp 1644511149
transform 1 0 22908 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_78_249
timestamp 1644511149
transform 1 0 24012 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_78_253
timestamp 1644511149
transform 1 0 24380 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_78_265
timestamp 1644511149
transform 1 0 25484 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_78_273
timestamp 1644511149
transform 1 0 26220 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_78_295
timestamp 1644511149
transform 1 0 28244 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_79_3
timestamp 1644511149
transform 1 0 1380 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_79_26
timestamp 1644511149
transform 1 0 3496 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_79_34
timestamp 1644511149
transform 1 0 4232 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_79_39
timestamp 1644511149
transform 1 0 4692 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_79_51
timestamp 1644511149
transform 1 0 5796 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_55
timestamp 1644511149
transform 1 0 6164 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_57
timestamp 1644511149
transform 1 0 6348 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_69
timestamp 1644511149
transform 1 0 7452 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_81
timestamp 1644511149
transform 1 0 8556 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_79_93
timestamp 1644511149
transform 1 0 9660 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_79_97
timestamp 1644511149
transform 1 0 10028 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_79_106
timestamp 1644511149
transform 1 0 10856 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_79_113
timestamp 1644511149
transform 1 0 11500 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_125
timestamp 1644511149
transform 1 0 12604 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_137
timestamp 1644511149
transform 1 0 13708 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_143
timestamp 1644511149
transform 1 0 14260 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_79_147
timestamp 1644511149
transform 1 0 14628 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_79_154
timestamp 1644511149
transform 1 0 15272 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_79_166
timestamp 1644511149
transform 1 0 16376 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_79_169
timestamp 1644511149
transform 1 0 16652 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_79_181
timestamp 1644511149
transform 1 0 17756 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_206
timestamp 1644511149
transform 1 0 20056 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_79_213
timestamp 1644511149
transform 1 0 20700 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_79_221
timestamp 1644511149
transform 1 0 21436 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_79_225
timestamp 1644511149
transform 1 0 21804 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_79_230
timestamp 1644511149
transform 1 0 22264 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_237
timestamp 1644511149
transform 1 0 22908 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_79_244
timestamp 1644511149
transform 1 0 23552 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_79_252
timestamp 1644511149
transform 1 0 24288 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_79_276
timestamp 1644511149
transform 1 0 26496 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_281
timestamp 1644511149
transform 1 0 26956 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_285
timestamp 1644511149
transform 1 0 27324 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_79_289
timestamp 1644511149
transform 1 0 27692 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_79_297
timestamp 1644511149
transform 1 0 28428 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_80_6
timestamp 1644511149
transform 1 0 1656 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_80_13
timestamp 1644511149
transform 1 0 2300 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_80_24
timestamp 1644511149
transform 1 0 3312 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_80_50
timestamp 1644511149
transform 1 0 5704 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_62
timestamp 1644511149
transform 1 0 6808 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_77
timestamp 1644511149
transform 1 0 8188 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_83
timestamp 1644511149
transform 1 0 8740 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_80_85
timestamp 1644511149
transform 1 0 8924 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_91
timestamp 1644511149
transform 1 0 9476 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_113
timestamp 1644511149
transform 1 0 11500 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_80_125
timestamp 1644511149
transform 1 0 12604 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_80_136
timestamp 1644511149
transform 1 0 13616 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_80_141
timestamp 1644511149
transform 1 0 14076 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_80_164
timestamp 1644511149
transform 1 0 16192 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_80_171
timestamp 1644511149
transform 1 0 16836 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_80_183
timestamp 1644511149
transform 1 0 17940 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_80_189
timestamp 1644511149
transform 1 0 18492 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_195
timestamp 1644511149
transform 1 0 19044 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_80_197
timestamp 1644511149
transform 1 0 19228 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_80_201
timestamp 1644511149
transform 1 0 19596 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_80_223
timestamp 1644511149
transform 1 0 21620 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_248
timestamp 1644511149
transform 1 0 23920 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_80_256
timestamp 1644511149
transform 1 0 24656 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_80_264
timestamp 1644511149
transform 1 0 25392 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_80_270
timestamp 1644511149
transform 1 0 25944 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_295
timestamp 1644511149
transform 1 0 28244 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_81_3
timestamp 1644511149
transform 1 0 1380 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_81_27
timestamp 1644511149
transform 1 0 3588 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_52
timestamp 1644511149
transform 1 0 5888 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_81_57
timestamp 1644511149
transform 1 0 6348 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_81_69
timestamp 1644511149
transform 1 0 7452 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_94
timestamp 1644511149
transform 1 0 9752 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_101
timestamp 1644511149
transform 1 0 10396 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_108
timestamp 1644511149
transform 1 0 11040 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_134
timestamp 1644511149
transform 1 0 13432 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_81_159
timestamp 1644511149
transform 1 0 15732 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_81_167
timestamp 1644511149
transform 1 0 16468 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_81_190
timestamp 1644511149
transform 1 0 18584 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_81_198
timestamp 1644511149
transform 1 0 19320 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_81_220
timestamp 1644511149
transform 1 0 21344 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_81_225
timestamp 1644511149
transform 1 0 21804 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_81_231
timestamp 1644511149
transform 1 0 22356 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_237
timestamp 1644511149
transform 1 0 22908 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_81_242
timestamp 1644511149
transform 1 0 23368 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_267
timestamp 1644511149
transform 1 0 25668 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_271
timestamp 1644511149
transform 1 0 26036 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_81_275
timestamp 1644511149
transform 1 0 26404 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_279
timestamp 1644511149
transform 1 0 26772 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_81_284
timestamp 1644511149
transform 1 0 27232 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_288
timestamp 1644511149
transform 1 0 27600 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_81_292
timestamp 1644511149
transform 1 0 27968 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_298
timestamp 1644511149
transform 1 0 28520 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_3
timestamp 1644511149
transform 1 0 1380 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_82_10
timestamp 1644511149
transform 1 0 2024 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_82_21
timestamp 1644511149
transform 1 0 3036 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_27
timestamp 1644511149
transform 1 0 3588 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_82_32
timestamp 1644511149
transform 1 0 4048 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_44
timestamp 1644511149
transform 1 0 5152 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_82_61
timestamp 1644511149
transform 1 0 6716 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_69
timestamp 1644511149
transform 1 0 7452 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_82_76
timestamp 1644511149
transform 1 0 8096 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_82_85
timestamp 1644511149
transform 1 0 8924 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_97
timestamp 1644511149
transform 1 0 10028 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_82_109
timestamp 1644511149
transform 1 0 11132 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_82_113
timestamp 1644511149
transform 1 0 11500 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_125
timestamp 1644511149
transform 1 0 12604 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_82_137
timestamp 1644511149
transform 1 0 13708 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_82_144
timestamp 1644511149
transform 1 0 14352 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_156
timestamp 1644511149
transform 1 0 15456 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_172
timestamp 1644511149
transform 1 0 16928 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_82_184
timestamp 1644511149
transform 1 0 18032 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_82_188
timestamp 1644511149
transform 1 0 18400 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_82_197
timestamp 1644511149
transform 1 0 19228 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_82_202
timestamp 1644511149
transform 1 0 19688 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_82_214
timestamp 1644511149
transform 1 0 20792 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_82_222
timestamp 1644511149
transform 1 0 21528 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_82_225
timestamp 1644511149
transform 1 0 21804 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_82_248
timestamp 1644511149
transform 1 0 23920 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_82_253
timestamp 1644511149
transform 1 0 24380 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_82_276
timestamp 1644511149
transform 1 0 26496 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_82_284
timestamp 1644511149
transform 1 0 27232 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_290
timestamp 1644511149
transform 1 0 27784 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_294
timestamp 1644511149
transform 1 0 28152 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_82_298
timestamp 1644511149
transform 1 0 28520 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1644511149
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1644511149
transform -1 0 28888 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1644511149
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1644511149
transform -1 0 28888 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1644511149
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1644511149
transform -1 0 28888 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1644511149
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1644511149
transform -1 0 28888 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1644511149
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1644511149
transform -1 0 28888 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1644511149
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1644511149
transform -1 0 28888 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1644511149
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1644511149
transform -1 0 28888 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1644511149
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1644511149
transform -1 0 28888 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1644511149
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1644511149
transform -1 0 28888 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1644511149
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1644511149
transform -1 0 28888 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1644511149
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1644511149
transform -1 0 28888 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1644511149
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1644511149
transform -1 0 28888 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1644511149
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1644511149
transform -1 0 28888 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1644511149
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1644511149
transform -1 0 28888 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1644511149
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1644511149
transform -1 0 28888 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1644511149
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1644511149
transform -1 0 28888 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1644511149
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1644511149
transform -1 0 28888 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1644511149
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1644511149
transform -1 0 28888 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1644511149
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1644511149
transform -1 0 28888 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1644511149
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1644511149
transform -1 0 28888 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1644511149
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1644511149
transform -1 0 28888 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1644511149
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1644511149
transform -1 0 28888 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1644511149
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1644511149
transform -1 0 28888 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1644511149
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1644511149
transform -1 0 28888 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1644511149
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1644511149
transform -1 0 28888 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1644511149
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1644511149
transform -1 0 28888 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1644511149
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1644511149
transform -1 0 28888 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1644511149
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1644511149
transform -1 0 28888 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1644511149
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1644511149
transform -1 0 28888 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1644511149
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1644511149
transform -1 0 28888 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1644511149
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1644511149
transform -1 0 28888 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1644511149
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1644511149
transform -1 0 28888 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1644511149
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1644511149
transform -1 0 28888 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1644511149
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1644511149
transform -1 0 28888 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1644511149
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1644511149
transform -1 0 28888 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1644511149
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1644511149
transform -1 0 28888 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1644511149
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1644511149
transform -1 0 28888 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1644511149
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1644511149
transform -1 0 28888 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1644511149
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1644511149
transform -1 0 28888 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1644511149
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1644511149
transform -1 0 28888 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1644511149
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1644511149
transform -1 0 28888 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1644511149
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1644511149
transform -1 0 28888 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1644511149
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1644511149
transform -1 0 28888 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1644511149
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1644511149
transform -1 0 28888 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1644511149
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1644511149
transform -1 0 28888 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1644511149
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1644511149
transform -1 0 28888 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1644511149
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1644511149
transform -1 0 28888 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1644511149
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1644511149
transform -1 0 28888 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1644511149
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1644511149
transform -1 0 28888 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1644511149
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1644511149
transform -1 0 28888 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1644511149
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1644511149
transform -1 0 28888 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1644511149
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1644511149
transform -1 0 28888 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1644511149
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1644511149
transform -1 0 28888 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1644511149
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1644511149
transform -1 0 28888 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1644511149
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1644511149
transform -1 0 28888 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1644511149
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1644511149
transform -1 0 28888 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1644511149
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1644511149
transform -1 0 28888 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1644511149
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1644511149
transform -1 0 28888 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1644511149
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1644511149
transform -1 0 28888 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1644511149
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1644511149
transform -1 0 28888 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1644511149
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1644511149
transform -1 0 28888 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1644511149
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1644511149
transform -1 0 28888 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1644511149
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1644511149
transform -1 0 28888 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1644511149
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1644511149
transform -1 0 28888 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1644511149
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1644511149
transform -1 0 28888 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 1644511149
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 1644511149
transform -1 0 28888 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 1644511149
transform 1 0 1104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 1644511149
transform -1 0 28888 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_134
timestamp 1644511149
transform 1 0 1104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_135
timestamp 1644511149
transform -1 0 28888 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_136
timestamp 1644511149
transform 1 0 1104 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_137
timestamp 1644511149
transform -1 0 28888 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_138
timestamp 1644511149
transform 1 0 1104 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_139
timestamp 1644511149
transform -1 0 28888 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_140
timestamp 1644511149
transform 1 0 1104 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_141
timestamp 1644511149
transform -1 0 28888 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_142
timestamp 1644511149
transform 1 0 1104 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_143
timestamp 1644511149
transform -1 0 28888 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_144
timestamp 1644511149
transform 1 0 1104 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_145
timestamp 1644511149
transform -1 0 28888 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_146
timestamp 1644511149
transform 1 0 1104 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_147
timestamp 1644511149
transform -1 0 28888 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_148
timestamp 1644511149
transform 1 0 1104 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_149
timestamp 1644511149
transform -1 0 28888 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_150
timestamp 1644511149
transform 1 0 1104 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_151
timestamp 1644511149
transform -1 0 28888 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_152
timestamp 1644511149
transform 1 0 1104 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_153
timestamp 1644511149
transform -1 0 28888 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_154
timestamp 1644511149
transform 1 0 1104 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_155
timestamp 1644511149
transform -1 0 28888 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_156
timestamp 1644511149
transform 1 0 1104 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_157
timestamp 1644511149
transform -1 0 28888 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_158
timestamp 1644511149
transform 1 0 1104 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_159
timestamp 1644511149
transform -1 0 28888 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_160
timestamp 1644511149
transform 1 0 1104 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_161
timestamp 1644511149
transform -1 0 28888 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_162
timestamp 1644511149
transform 1 0 1104 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_163
timestamp 1644511149
transform -1 0 28888 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_164
timestamp 1644511149
transform 1 0 1104 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_165
timestamp 1644511149
transform -1 0 28888 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1644511149
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1644511149
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1644511149
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1644511149
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1644511149
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1644511149
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1644511149
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1644511149
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1644511149
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1644511149
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1644511149
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1644511149
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1644511149
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1644511149
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1644511149
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1644511149
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1644511149
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1644511149
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1644511149
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1644511149
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1644511149
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1644511149
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1644511149
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1644511149
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1644511149
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1644511149
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1644511149
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1644511149
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1644511149
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1644511149
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1644511149
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1644511149
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1644511149
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1644511149
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1644511149
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1644511149
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1644511149
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1644511149
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1644511149
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1644511149
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1644511149
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1644511149
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1644511149
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1644511149
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1644511149
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1644511149
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1644511149
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1644511149
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1644511149
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1644511149
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1644511149
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1644511149
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1644511149
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1644511149
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1644511149
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1644511149
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1644511149
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1644511149
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1644511149
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1644511149
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1644511149
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1644511149
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1644511149
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1644511149
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1644511149
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1644511149
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1644511149
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1644511149
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1644511149
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1644511149
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1644511149
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1644511149
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1644511149
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1644511149
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1644511149
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1644511149
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1644511149
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1644511149
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1644511149
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1644511149
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1644511149
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1644511149
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1644511149
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1644511149
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1644511149
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1644511149
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1644511149
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1644511149
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1644511149
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1644511149
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1644511149
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1644511149
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1644511149
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1644511149
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1644511149
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1644511149
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1644511149
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1644511149
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1644511149
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1644511149
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1644511149
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1644511149
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1644511149
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1644511149
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1644511149
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1644511149
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1644511149
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1644511149
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1644511149
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1644511149
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1644511149
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1644511149
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1644511149
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1644511149
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1644511149
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1644511149
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1644511149
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1644511149
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1644511149
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1644511149
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1644511149
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1644511149
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1644511149
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1644511149
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1644511149
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1644511149
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1644511149
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1644511149
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1644511149
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1644511149
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1644511149
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1644511149
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1644511149
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1644511149
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1644511149
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1644511149
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1644511149
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1644511149
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1644511149
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1644511149
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1644511149
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1644511149
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1644511149
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1644511149
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1644511149
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1644511149
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1644511149
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1644511149
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1644511149
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1644511149
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1644511149
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1644511149
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1644511149
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1644511149
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1644511149
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1644511149
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1644511149
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1644511149
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1644511149
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1644511149
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1644511149
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1644511149
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1644511149
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1644511149
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1644511149
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1644511149
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1644511149
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1644511149
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1644511149
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1644511149
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1644511149
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1644511149
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1644511149
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1644511149
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1644511149
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1644511149
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1644511149
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1644511149
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1644511149
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1644511149
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1644511149
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1644511149
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1644511149
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1644511149
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1644511149
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1644511149
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1644511149
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1644511149
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1644511149
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1644511149
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1644511149
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1644511149
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1644511149
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1644511149
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1644511149
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1644511149
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1644511149
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1644511149
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1644511149
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1644511149
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1644511149
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1644511149
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1644511149
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1644511149
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1644511149
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1644511149
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1644511149
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1644511149
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1644511149
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1644511149
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1644511149
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1644511149
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1644511149
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1644511149
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1644511149
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1644511149
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1644511149
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1644511149
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1644511149
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1644511149
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1644511149
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1644511149
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1644511149
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1644511149
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1644511149
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1644511149
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1644511149
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1644511149
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1644511149
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1644511149
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1644511149
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1644511149
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1644511149
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1644511149
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1644511149
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1644511149
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1644511149
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1644511149
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1644511149
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1644511149
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1644511149
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1644511149
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1644511149
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1644511149
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1644511149
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1644511149
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1644511149
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1644511149
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1644511149
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1644511149
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1644511149
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1644511149
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1644511149
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1644511149
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1644511149
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1644511149
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1644511149
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1644511149
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1644511149
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1644511149
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1644511149
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1644511149
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1644511149
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1644511149
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1644511149
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1644511149
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1644511149
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1644511149
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1644511149
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1644511149
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1644511149
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1644511149
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1644511149
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1644511149
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1644511149
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1644511149
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1644511149
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1644511149
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1644511149
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1644511149
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1644511149
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1644511149
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1644511149
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1644511149
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1644511149
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1644511149
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1644511149
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1644511149
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1644511149
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1644511149
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1644511149
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1644511149
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1644511149
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1644511149
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1644511149
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1644511149
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1644511149
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1644511149
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1644511149
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1644511149
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1644511149
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1644511149
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1644511149
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1644511149
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1644511149
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1644511149
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1644511149
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1644511149
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1644511149
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1644511149
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1644511149
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1644511149
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1644511149
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1644511149
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1644511149
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1644511149
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1644511149
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1644511149
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1644511149
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1644511149
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1644511149
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1644511149
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1644511149
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1644511149
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1644511149
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1644511149
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1644511149
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1644511149
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1644511149
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1644511149
transform 1 0 6256 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1644511149
transform 1 0 11408 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1644511149
transform 1 0 16560 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1644511149
transform 1 0 21712 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1644511149
transform 1 0 26864 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1644511149
transform 1 0 3680 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1644511149
transform 1 0 8832 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1644511149
transform 1 0 13984 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1644511149
transform 1 0 19136 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1644511149
transform 1 0 24288 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1644511149
transform 1 0 6256 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1644511149
transform 1 0 11408 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1644511149
transform 1 0 16560 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1644511149
transform 1 0 21712 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1644511149
transform 1 0 26864 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1644511149
transform 1 0 3680 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1644511149
transform 1 0 8832 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1644511149
transform 1 0 13984 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1644511149
transform 1 0 19136 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1644511149
transform 1 0 24288 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1644511149
transform 1 0 6256 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1644511149
transform 1 0 11408 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1644511149
transform 1 0 16560 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1644511149
transform 1 0 21712 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1644511149
transform 1 0 26864 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1644511149
transform 1 0 3680 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1644511149
transform 1 0 8832 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1644511149
transform 1 0 13984 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1644511149
transform 1 0 19136 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1644511149
transform 1 0 24288 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1644511149
transform 1 0 6256 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1644511149
transform 1 0 11408 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1644511149
transform 1 0 16560 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1644511149
transform 1 0 21712 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1644511149
transform 1 0 26864 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1644511149
transform 1 0 3680 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1644511149
transform 1 0 8832 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1644511149
transform 1 0 13984 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1644511149
transform 1 0 19136 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1644511149
transform 1 0 24288 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1644511149
transform 1 0 6256 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1644511149
transform 1 0 11408 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1644511149
transform 1 0 16560 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1644511149
transform 1 0 21712 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1644511149
transform 1 0 26864 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1644511149
transform 1 0 3680 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1644511149
transform 1 0 8832 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1644511149
transform 1 0 13984 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1644511149
transform 1 0 19136 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1644511149
transform 1 0 24288 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1644511149
transform 1 0 6256 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1644511149
transform 1 0 11408 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1644511149
transform 1 0 16560 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1644511149
transform 1 0 21712 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1644511149
transform 1 0 26864 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1644511149
transform 1 0 3680 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1644511149
transform 1 0 8832 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1644511149
transform 1 0 13984 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1644511149
transform 1 0 19136 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1644511149
transform 1 0 24288 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1644511149
transform 1 0 6256 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1644511149
transform 1 0 11408 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1644511149
transform 1 0 16560 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1644511149
transform 1 0 21712 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1644511149
transform 1 0 26864 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1644511149
transform 1 0 3680 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1644511149
transform 1 0 8832 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1644511149
transform 1 0 13984 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1644511149
transform 1 0 19136 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1644511149
transform 1 0 24288 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1644511149
transform 1 0 6256 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1644511149
transform 1 0 11408 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1644511149
transform 1 0 16560 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1644511149
transform 1 0 21712 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1644511149
transform 1 0 26864 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1644511149
transform 1 0 3680 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1644511149
transform 1 0 8832 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1644511149
transform 1 0 13984 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1644511149
transform 1 0 19136 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1644511149
transform 1 0 24288 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1644511149
transform 1 0 6256 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1644511149
transform 1 0 11408 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1644511149
transform 1 0 16560 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1644511149
transform 1 0 21712 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1644511149
transform 1 0 26864 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1644511149
transform 1 0 3680 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1644511149
transform 1 0 6256 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1644511149
transform 1 0 8832 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1644511149
transform 1 0 11408 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1644511149
transform 1 0 13984 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1644511149
transform 1 0 16560 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1644511149
transform 1 0 19136 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1644511149
transform 1 0 21712 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1644511149
transform 1 0 24288 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1644511149
transform 1 0 26864 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _0528_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 16836 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  _0529_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 17940 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _0530_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 22632 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0531_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 23368 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0532_
timestamp 1644511149
transform 1 0 6348 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0533_
timestamp 1644511149
transform -1 0 2116 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0534_
timestamp 1644511149
transform 1 0 16284 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0535_
timestamp 1644511149
transform -1 0 2116 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0536_
timestamp 1644511149
transform 1 0 18216 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0537_
timestamp 1644511149
transform 1 0 27692 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0538_
timestamp 1644511149
transform -1 0 3036 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0539_
timestamp 1644511149
transform 1 0 27968 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0540_
timestamp 1644511149
transform -1 0 2392 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0541_
timestamp 1644511149
transform 1 0 27692 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0542_
timestamp 1644511149
transform 1 0 25116 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  _0543_
timestamp 1644511149
transform 1 0 27692 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0544_
timestamp 1644511149
transform -1 0 27784 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0545_
timestamp 1644511149
transform -1 0 27232 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0546_
timestamp 1644511149
transform 1 0 27692 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0547_
timestamp 1644511149
transform -1 0 25576 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0548_
timestamp 1644511149
transform -1 0 27876 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _0549_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 25392 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0550_
timestamp 1644511149
transform -1 0 2392 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0551_
timestamp 1644511149
transform -1 0 11776 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0552_
timestamp 1644511149
transform -1 0 2484 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0553_
timestamp 1644511149
transform 1 0 27876 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0554_
timestamp 1644511149
transform -1 0 27876 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0555_
timestamp 1644511149
transform 1 0 27692 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0556_
timestamp 1644511149
transform -1 0 2208 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0557_
timestamp 1644511149
transform -1 0 28060 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0558_
timestamp 1644511149
transform 1 0 27784 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0559_
timestamp 1644511149
transform -1 0 2852 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0560_
timestamp 1644511149
transform 1 0 27784 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _0561_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 25484 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0562_
timestamp 1644511149
transform -1 0 4048 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0563_
timestamp 1644511149
transform 1 0 27508 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0564_
timestamp 1644511149
transform 1 0 14352 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0565_
timestamp 1644511149
transform 1 0 9200 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0566_
timestamp 1644511149
transform 1 0 27508 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _0567_
timestamp 1644511149
transform 1 0 26956 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0568_
timestamp 1644511149
transform -1 0 2300 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0569_
timestamp 1644511149
transform 1 0 27784 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0570_
timestamp 1644511149
transform -1 0 2300 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0571_
timestamp 1644511149
transform -1 0 27692 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0572_
timestamp 1644511149
transform -1 0 4416 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0573_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 26956 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_8  _0574_
timestamp 1644511149
transform 1 0 26036 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0575_
timestamp 1644511149
transform -1 0 27416 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0576_
timestamp 1644511149
transform 1 0 27416 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0577_
timestamp 1644511149
transform 1 0 16560 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0578_
timestamp 1644511149
transform 1 0 5244 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0579_
timestamp 1644511149
transform -1 0 2760 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _0580_
timestamp 1644511149
transform 1 0 25392 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0581_
timestamp 1644511149
transform 1 0 27048 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0582_
timestamp 1644511149
transform 1 0 7912 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0583_
timestamp 1644511149
transform 1 0 26956 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0584_
timestamp 1644511149
transform -1 0 4048 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0585_
timestamp 1644511149
transform -1 0 14720 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0586_
timestamp 1644511149
transform -1 0 25668 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0587_
timestamp 1644511149
transform 1 0 24840 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0588_
timestamp 1644511149
transform -1 0 27232 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0589_
timestamp 1644511149
transform -1 0 24748 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0590_
timestamp 1644511149
transform 1 0 25116 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0591_
timestamp 1644511149
transform 1 0 27416 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _0592_
timestamp 1644511149
transform 1 0 27324 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0593_
timestamp 1644511149
transform -1 0 27232 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0594_
timestamp 1644511149
transform 1 0 26956 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0595_
timestamp 1644511149
transform -1 0 27232 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0596_
timestamp 1644511149
transform -1 0 25944 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0597_
timestamp 1644511149
transform -1 0 27416 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _0598_
timestamp 1644511149
transform -1 0 25944 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0599_
timestamp 1644511149
transform -1 0 2024 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0600_
timestamp 1644511149
transform 1 0 21988 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0601_
timestamp 1644511149
transform -1 0 2024 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0602_
timestamp 1644511149
transform -1 0 27876 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0603_
timestamp 1644511149
transform 1 0 27968 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0604_
timestamp 1644511149
transform -1 0 5060 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_8  _0605_
timestamp 1644511149
transform 1 0 4784 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0606_
timestamp 1644511149
transform 1 0 27692 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0607_
timestamp 1644511149
transform -1 0 3036 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0608_
timestamp 1644511149
transform 1 0 27692 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0609_
timestamp 1644511149
transform -1 0 3128 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0610_
timestamp 1644511149
transform 1 0 27692 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _0611_
timestamp 1644511149
transform 1 0 4876 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0612_
timestamp 1644511149
transform -1 0 25944 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0613_
timestamp 1644511149
transform 1 0 26956 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0614_
timestamp 1644511149
transform -1 0 4692 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0615_
timestamp 1644511149
transform -1 0 22908 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0616_
timestamp 1644511149
transform 1 0 19504 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0617_
timestamp 1644511149
transform 1 0 6348 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0618_
timestamp 1644511149
transform -1 0 1840 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0619_
timestamp 1644511149
transform -1 0 27324 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0620_
timestamp 1644511149
transform -1 0 1932 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0621_
timestamp 1644511149
transform -1 0 1840 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0622_
timestamp 1644511149
transform 1 0 27692 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0623_
timestamp 1644511149
transform -1 0 4416 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0624_
timestamp 1644511149
transform -1 0 2024 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0625_
timestamp 1644511149
transform -1 0 2116 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0626_
timestamp 1644511149
transform 1 0 2760 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0627_
timestamp 1644511149
transform 1 0 7452 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0628_
timestamp 1644511149
transform -1 0 2116 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _0629_
timestamp 1644511149
transform -1 0 5704 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0630_
timestamp 1644511149
transform 1 0 27692 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0631_
timestamp 1644511149
transform -1 0 27784 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0632_
timestamp 1644511149
transform 1 0 27692 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0633_
timestamp 1644511149
transform -1 0 2208 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0634_
timestamp 1644511149
transform -1 0 2300 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _0635_
timestamp 1644511149
transform 1 0 17572 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0636_
timestamp 1644511149
transform 1 0 27968 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0637_
timestamp 1644511149
transform 1 0 10488 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0638_
timestamp 1644511149
transform 1 0 18216 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0639_
timestamp 1644511149
transform -1 0 3312 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0640_
timestamp 1644511149
transform 1 0 27600 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _0641_
timestamp 1644511149
transform 1 0 17940 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0642_
timestamp 1644511149
transform -1 0 4048 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0643_
timestamp 1644511149
transform -1 0 4692 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0644_
timestamp 1644511149
transform -1 0 10028 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0645_
timestamp 1644511149
transform 1 0 10580 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0646_
timestamp 1644511149
transform 1 0 25668 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _0647_
timestamp 1644511149
transform 1 0 17940 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0648_
timestamp 1644511149
transform -1 0 27232 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0649_
timestamp 1644511149
transform -1 0 13616 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0650_
timestamp 1644511149
transform 1 0 27232 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0651_
timestamp 1644511149
transform 1 0 20608 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0652_
timestamp 1644511149
transform 1 0 19412 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _0653_
timestamp 1644511149
transform 1 0 17940 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0654_
timestamp 1644511149
transform -1 0 1840 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0655_
timestamp 1644511149
transform 1 0 20424 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0656_
timestamp 1644511149
transform 1 0 13064 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0657_
timestamp 1644511149
transform -1 0 2024 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0658_
timestamp 1644511149
transform 1 0 2668 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _0659_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 17940 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0660_
timestamp 1644511149
transform 1 0 20792 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0661_
timestamp 1644511149
transform 1 0 23276 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0662_
timestamp 1644511149
transform -1 0 19964 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0663_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 18676 0 1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _0664_
timestamp 1644511149
transform 1 0 16836 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _0665_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 17296 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _0666_
timestamp 1644511149
transform 1 0 17480 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0667_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 18216 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _0668_
timestamp 1644511149
transform 1 0 17388 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0669_
timestamp 1644511149
transform 1 0 17480 0 1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__and2b_1  _0670_
timestamp 1644511149
transform 1 0 17296 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0671_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 18308 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _0672_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 17112 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _0673_
timestamp 1644511149
transform 1 0 16560 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _0674_
timestamp 1644511149
transform 1 0 16652 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__a21boi_1  _0675_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 18124 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _0676_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 17572 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0677_
timestamp 1644511149
transform 1 0 18584 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _0678_
timestamp 1644511149
transform 1 0 18676 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _0679_
timestamp 1644511149
transform -1 0 19412 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _0680_
timestamp 1644511149
transform 1 0 17020 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__a2111o_1  _0681_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 17940 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0682_
timestamp 1644511149
transform 1 0 19228 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _0683_
timestamp 1644511149
transform 1 0 19228 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0684_
timestamp 1644511149
transform 1 0 19228 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0685_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 20056 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__or2b_1  _0686_
timestamp 1644511149
transform 1 0 17112 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__and4b_1  _0687_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 18768 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0688_
timestamp 1644511149
transform -1 0 14996 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _0689_
timestamp 1644511149
transform -1 0 14628 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _0690_
timestamp 1644511149
transform -1 0 16008 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _0691_
timestamp 1644511149
transform 1 0 13432 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__a2111o_1  _0692_
timestamp 1644511149
transform -1 0 14904 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0693_
timestamp 1644511149
transform 1 0 14996 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _0694_
timestamp 1644511149
transform -1 0 14720 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0695_
timestamp 1644511149
transform 1 0 15916 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0696_
timestamp 1644511149
transform 1 0 16652 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__or2b_1  _0697_
timestamp 1644511149
transform 1 0 13248 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__and4b_1  _0698_
timestamp 1644511149
transform 1 0 14352 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__nand3b_1  _0699_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 17848 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__o311a_1  _0700_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 14168 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _0701_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 20792 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _0702_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 19872 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _0703_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 18676 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0704_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 17296 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0705_
timestamp 1644511149
transform 1 0 18860 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0706_
timestamp 1644511149
transform -1 0 18492 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__and4_1  _0707_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 17848 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0708_
timestamp 1644511149
transform 1 0 18308 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _0709_
timestamp 1644511149
transform -1 0 24748 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _0710_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 20792 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__or3_2  _0711_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 20976 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _0712_
timestamp 1644511149
transform 1 0 20700 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0713_
timestamp 1644511149
transform 1 0 21620 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _0714_
timestamp 1644511149
transform 1 0 19228 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _0715_
timestamp 1644511149
transform 1 0 19228 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0716_
timestamp 1644511149
transform 1 0 19044 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0717_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 20792 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0718_
timestamp 1644511149
transform -1 0 20056 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0719_
timestamp 1644511149
transform 1 0 19964 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _0720_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 19228 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _0721_
timestamp 1644511149
transform -1 0 21528 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _0722_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 21252 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _0723_
timestamp 1644511149
transform -1 0 20332 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0724_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 25208 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0725_
timestamp 1644511149
transform 1 0 24932 0 -1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  _0726_
timestamp 1644511149
transform -1 0 24748 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0727_
timestamp 1644511149
transform 1 0 25392 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0728_
timestamp 1644511149
transform 1 0 25576 0 -1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__nor2b_1  _0729_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 26956 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0730_
timestamp 1644511149
transform -1 0 25852 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__or2b_1  _0731_
timestamp 1644511149
transform 1 0 25392 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0732_
timestamp 1644511149
transform -1 0 26036 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0733_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 25024 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _0734_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 27324 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0735_
timestamp 1644511149
transform 1 0 25576 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0736_
timestamp 1644511149
transform -1 0 26496 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _0737_
timestamp 1644511149
transform 1 0 25484 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0738_
timestamp 1644511149
transform 1 0 24932 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0739_
timestamp 1644511149
transform -1 0 25760 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _0740_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 25208 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0741_
timestamp 1644511149
transform -1 0 24656 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0742_
timestamp 1644511149
transform -1 0 27876 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _0743_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 26956 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0744_
timestamp 1644511149
transform -1 0 25944 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _0745_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 26956 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0746_
timestamp 1644511149
transform 1 0 26864 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0747_
timestamp 1644511149
transform -1 0 25116 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _0748_
timestamp 1644511149
transform -1 0 27600 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0749_
timestamp 1644511149
transform -1 0 26220 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0750_
timestamp 1644511149
transform 1 0 20148 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0751_
timestamp 1644511149
transform 1 0 20240 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0752_
timestamp 1644511149
transform -1 0 23000 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0753_
timestamp 1644511149
transform -1 0 19872 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_2  _0754_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 20148 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0755_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 19688 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0756_
timestamp 1644511149
transform 1 0 18492 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0757_
timestamp 1644511149
transform -1 0 22816 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0758_
timestamp 1644511149
transform -1 0 20332 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0759_
timestamp 1644511149
transform -1 0 19504 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _0760_
timestamp 1644511149
transform -1 0 20424 0 -1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_2  _0761_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 19964 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0762_
timestamp 1644511149
transform 1 0 21804 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0763_
timestamp 1644511149
transform 1 0 22080 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0764_
timestamp 1644511149
transform 1 0 21252 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0765_
timestamp 1644511149
transform 1 0 21712 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0766_
timestamp 1644511149
transform -1 0 23736 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _0767_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 21804 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__o221ai_1  _0768_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 21896 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _0769_
timestamp 1644511149
transform 1 0 21068 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _0770_
timestamp 1644511149
transform -1 0 23092 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _0771_
timestamp 1644511149
transform -1 0 22816 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0772_
timestamp 1644511149
transform -1 0 23920 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0773_
timestamp 1644511149
transform 1 0 23460 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_1  _0774_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 22264 0 -1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__o32a_1  _0775_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 22448 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0776_
timestamp 1644511149
transform -1 0 22264 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0777_
timestamp 1644511149
transform -1 0 22540 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _0778_
timestamp 1644511149
transform -1 0 23368 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _0779_
timestamp 1644511149
transform -1 0 21160 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _0780_
timestamp 1644511149
transform -1 0 21620 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _0781_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 22264 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0782_
timestamp 1644511149
transform -1 0 21528 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0783_
timestamp 1644511149
transform 1 0 20240 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0784_
timestamp 1644511149
transform -1 0 19872 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _0785_
timestamp 1644511149
transform 1 0 20608 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0786_
timestamp 1644511149
transform -1 0 21252 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__o311a_1  _0787_
timestamp 1644511149
transform 1 0 19688 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0788_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 20792 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0789_
timestamp 1644511149
transform 1 0 21068 0 1 38080
box -38 -48 958 592
use sky130_fd_sc_hd__a21oi_1  _0790_
timestamp 1644511149
transform 1 0 19872 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0791_
timestamp 1644511149
transform 1 0 20056 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _0792_
timestamp 1644511149
transform 1 0 19872 0 -1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0793_
timestamp 1644511149
transform 1 0 19412 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0794_
timestamp 1644511149
transform -1 0 21528 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0795_
timestamp 1644511149
transform -1 0 21344 0 -1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0796_
timestamp 1644511149
transform 1 0 20884 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _0797_
timestamp 1644511149
transform 1 0 20424 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _0798_
timestamp 1644511149
transform -1 0 21436 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__o211ai_1  _0799_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 21804 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _0800_
timestamp 1644511149
transform -1 0 22908 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _0801_
timestamp 1644511149
transform -1 0 20056 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _0802_
timestamp 1644511149
transform 1 0 20424 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _0803_
timestamp 1644511149
transform 1 0 21804 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0804_
timestamp 1644511149
transform 1 0 20148 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__nor3_1  _0805_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 19320 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0806_
timestamp 1644511149
transform 1 0 21160 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _0807_
timestamp 1644511149
transform 1 0 23092 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0808_
timestamp 1644511149
transform 1 0 22264 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0809_
timestamp 1644511149
transform -1 0 23000 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0810_
timestamp 1644511149
transform -1 0 23184 0 1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  _0811_
timestamp 1644511149
transform 1 0 24748 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0812_
timestamp 1644511149
transform 1 0 24288 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0813_
timestamp 1644511149
transform 1 0 25116 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0814_
timestamp 1644511149
transform -1 0 25208 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0815_
timestamp 1644511149
transform -1 0 24932 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _0816_
timestamp 1644511149
transform 1 0 25024 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _0817_
timestamp 1644511149
transform -1 0 21068 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _0818_
timestamp 1644511149
transform 1 0 23460 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0819_
timestamp 1644511149
transform -1 0 23552 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0820_
timestamp 1644511149
transform 1 0 22816 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0821_
timestamp 1644511149
transform -1 0 23368 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0822_
timestamp 1644511149
transform -1 0 23276 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0823_
timestamp 1644511149
transform -1 0 22356 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0824_
timestamp 1644511149
transform 1 0 23460 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0825_
timestamp 1644511149
transform -1 0 24104 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0826_
timestamp 1644511149
transform -1 0 23828 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0827_
timestamp 1644511149
transform -1 0 23092 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0828_
timestamp 1644511149
transform 1 0 23184 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0829_
timestamp 1644511149
transform -1 0 23552 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0830_
timestamp 1644511149
transform -1 0 21344 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _0831_
timestamp 1644511149
transform 1 0 21068 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0832_
timestamp 1644511149
transform 1 0 20792 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0833_
timestamp 1644511149
transform -1 0 21344 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0834_
timestamp 1644511149
transform -1 0 17480 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0835_
timestamp 1644511149
transform 1 0 15916 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _0836_
timestamp 1644511149
transform 1 0 12236 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _0837_
timestamp 1644511149
transform 1 0 12512 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0838_
timestamp 1644511149
transform -1 0 12420 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0839_
timestamp 1644511149
transform 1 0 12696 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _0840_
timestamp 1644511149
transform 1 0 12512 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0841_
timestamp 1644511149
transform 1 0 13340 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0842_
timestamp 1644511149
transform 1 0 17112 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _0843_
timestamp 1644511149
transform -1 0 17296 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0844_
timestamp 1644511149
transform -1 0 16744 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0845_
timestamp 1644511149
transform 1 0 17296 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _0846_
timestamp 1644511149
transform -1 0 17388 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0847_
timestamp 1644511149
transform -1 0 16928 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0848_
timestamp 1644511149
transform 1 0 15364 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _0849_
timestamp 1644511149
transform 1 0 12236 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0850_
timestamp 1644511149
transform -1 0 12604 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0851_
timestamp 1644511149
transform -1 0 11500 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0852_
timestamp 1644511149
transform 1 0 12236 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _0853_
timestamp 1644511149
transform 1 0 12052 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0854_
timestamp 1644511149
transform 1 0 12880 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0855_
timestamp 1644511149
transform 1 0 12328 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0856_
timestamp 1644511149
transform 1 0 11960 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0857_
timestamp 1644511149
transform 1 0 12788 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0858_
timestamp 1644511149
transform 1 0 14168 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _0859_
timestamp 1644511149
transform 1 0 14168 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0860_
timestamp 1644511149
transform -1 0 13616 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0861_
timestamp 1644511149
transform 1 0 16744 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0862_
timestamp 1644511149
transform -1 0 16744 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0863_
timestamp 1644511149
transform -1 0 16192 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0864_
timestamp 1644511149
transform 1 0 20148 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0865_
timestamp 1644511149
transform 1 0 19780 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0866_
timestamp 1644511149
transform 1 0 19872 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0867_
timestamp 1644511149
transform 1 0 14720 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _0868_
timestamp 1644511149
transform 1 0 14628 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0869_
timestamp 1644511149
transform 1 0 15456 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0870_
timestamp 1644511149
transform -1 0 20976 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0871_
timestamp 1644511149
transform 1 0 20424 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0872_
timestamp 1644511149
transform 1 0 21160 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0873_
timestamp 1644511149
transform -1 0 20700 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0874_
timestamp 1644511149
transform 1 0 21068 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0875_
timestamp 1644511149
transform -1 0 19228 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0876_
timestamp 1644511149
transform -1 0 17388 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0877_
timestamp 1644511149
transform 1 0 20240 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__a21boi_1  _0878_
timestamp 1644511149
transform -1 0 22356 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _0879_
timestamp 1644511149
transform 1 0 21804 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _0880_
timestamp 1644511149
transform 1 0 21804 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__a21boi_1  _0881_
timestamp 1644511149
transform -1 0 23276 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _0882_
timestamp 1644511149
transform 1 0 21436 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _0883_
timestamp 1644511149
transform -1 0 22448 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__a21boi_1  _0884_
timestamp 1644511149
transform -1 0 22540 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _0885_
timestamp 1644511149
transform 1 0 21804 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _0886_
timestamp 1644511149
transform 1 0 21804 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__a21boi_1  _0887_
timestamp 1644511149
transform -1 0 21344 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _0888_
timestamp 1644511149
transform 1 0 20608 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _0889_
timestamp 1644511149
transform 1 0 20608 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0890_
timestamp 1644511149
transform 1 0 21804 0 -1 25024
box -38 -48 958 592
use sky130_fd_sc_hd__a21oi_2  _0891_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 20240 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0892_
timestamp 1644511149
transform 1 0 23644 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0893_
timestamp 1644511149
transform -1 0 22816 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0894_
timestamp 1644511149
transform -1 0 23644 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _0895_
timestamp 1644511149
transform -1 0 23920 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0896_
timestamp 1644511149
transform 1 0 22264 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _0897_
timestamp 1644511149
transform -1 0 22448 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0898_
timestamp 1644511149
transform 1 0 22448 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0899_
timestamp 1644511149
transform 1 0 23000 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _0900_
timestamp 1644511149
transform -1 0 23736 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _0901_
timestamp 1644511149
transform -1 0 22172 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _0902_
timestamp 1644511149
transform 1 0 22264 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0903_
timestamp 1644511149
transform -1 0 21896 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0904_
timestamp 1644511149
transform -1 0 24564 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0905_
timestamp 1644511149
transform -1 0 22264 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _0906_
timestamp 1644511149
transform 1 0 22632 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0907_
timestamp 1644511149
transform -1 0 23000 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0908_
timestamp 1644511149
transform -1 0 23736 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _0909_
timestamp 1644511149
transform -1 0 23828 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0910_
timestamp 1644511149
transform -1 0 19136 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _0911_
timestamp 1644511149
transform -1 0 19964 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _0912_
timestamp 1644511149
transform -1 0 16192 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0913_
timestamp 1644511149
transform 1 0 17480 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0914_
timestamp 1644511149
transform -1 0 17112 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _0915_
timestamp 1644511149
transform 1 0 16376 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _0916_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 16008 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _0917_
timestamp 1644511149
transform 1 0 15088 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0918_
timestamp 1644511149
transform -1 0 18584 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0919_
timestamp 1644511149
transform -1 0 16192 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0920_
timestamp 1644511149
transform 1 0 16652 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0921_
timestamp 1644511149
transform 1 0 15732 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0922_
timestamp 1644511149
transform 1 0 16652 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0923_
timestamp 1644511149
transform 1 0 15364 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__and4_1  _0924_
timestamp 1644511149
transform -1 0 16560 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0925_
timestamp 1644511149
transform -1 0 15548 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0926_
timestamp 1644511149
transform -1 0 15364 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0927_
timestamp 1644511149
transform 1 0 14536 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0928_
timestamp 1644511149
transform 1 0 15088 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _0929_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 16008 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0930_
timestamp 1644511149
transform -1 0 15272 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0931_
timestamp 1644511149
transform -1 0 14352 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0932_
timestamp 1644511149
transform 1 0 15640 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0933_
timestamp 1644511149
transform -1 0 15916 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0934_
timestamp 1644511149
transform -1 0 14444 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0935_
timestamp 1644511149
transform -1 0 15272 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0936_
timestamp 1644511149
transform 1 0 14076 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0937_
timestamp 1644511149
transform 1 0 15272 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0938_
timestamp 1644511149
transform -1 0 15916 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0939_
timestamp 1644511149
transform -1 0 15272 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0940_
timestamp 1644511149
transform -1 0 15548 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0941_
timestamp 1644511149
transform 1 0 14076 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0942_
timestamp 1644511149
transform 1 0 16192 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0943_
timestamp 1644511149
transform 1 0 15364 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0944_
timestamp 1644511149
transform 1 0 15364 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0945_
timestamp 1644511149
transform 1 0 15548 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0946_
timestamp 1644511149
transform -1 0 18492 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0947_
timestamp 1644511149
transform -1 0 17112 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _0948_
timestamp 1644511149
transform -1 0 15824 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _0949_
timestamp 1644511149
transform -1 0 16560 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _0950_
timestamp 1644511149
transform -1 0 17204 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0951_
timestamp 1644511149
transform 1 0 16928 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0952_
timestamp 1644511149
transform 1 0 16284 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _0953_
timestamp 1644511149
transform 1 0 17112 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _0954_
timestamp 1644511149
transform -1 0 18400 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0955_
timestamp 1644511149
transform -1 0 17756 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0956_
timestamp 1644511149
transform 1 0 17848 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0957_
timestamp 1644511149
transform 1 0 17020 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0958_
timestamp 1644511149
transform 1 0 17204 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a21boi_1  _0959_
timestamp 1644511149
transform 1 0 17296 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _0960_
timestamp 1644511149
transform 1 0 21528 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _0961_
timestamp 1644511149
transform -1 0 22540 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _0962_
timestamp 1644511149
transform -1 0 25208 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0963_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 23184 0 -1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0964_
timestamp 1644511149
transform -1 0 24748 0 -1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0965_
timestamp 1644511149
transform 1 0 18768 0 -1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0966_
timestamp 1644511149
transform 1 0 19228 0 1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0967_
timestamp 1644511149
transform -1 0 23828 0 1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0968_
timestamp 1644511149
transform 1 0 19228 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0969_
timestamp 1644511149
transform -1 0 20884 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0970_
timestamp 1644511149
transform 1 0 18216 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0971_
timestamp 1644511149
transform 1 0 18860 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0972_
timestamp 1644511149
transform 1 0 22816 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0973_
timestamp 1644511149
transform 1 0 24472 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0974_
timestamp 1644511149
transform 1 0 24932 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0975_
timestamp 1644511149
transform 1 0 22448 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0976_
timestamp 1644511149
transform 1 0 22724 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0977_
timestamp 1644511149
transform 1 0 24380 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0978_
timestamp 1644511149
transform 1 0 23460 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0979_
timestamp 1644511149
transform 1 0 21804 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0980_
timestamp 1644511149
transform 1 0 25852 0 1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0981_
timestamp 1644511149
transform -1 0 26496 0 -1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0982_
timestamp 1644511149
transform 1 0 17940 0 -1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0983_
timestamp 1644511149
transform 1 0 12144 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0984_
timestamp 1644511149
transform -1 0 13616 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0985_
timestamp 1644511149
transform 1 0 16652 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0986_
timestamp 1644511149
transform 1 0 16836 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0987_
timestamp 1644511149
transform 1 0 11868 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0988_
timestamp 1644511149
transform 1 0 11960 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0989_
timestamp 1644511149
transform 1 0 11960 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0990_
timestamp 1644511149
transform 1 0 13340 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0991_
timestamp 1644511149
transform 1 0 16652 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0992_
timestamp 1644511149
transform 1 0 19504 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _0993_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 14628 0 -1 30464
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _0994_
timestamp 1644511149
transform -1 0 20792 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0995_
timestamp 1644511149
transform 1 0 19688 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0996_
timestamp 1644511149
transform 1 0 20976 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0997_
timestamp 1644511149
transform 1 0 21988 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0998_
timestamp 1644511149
transform 1 0 21436 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0999_
timestamp 1644511149
transform 1 0 19780 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1000_
timestamp 1644511149
transform -1 0 25852 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1001_
timestamp 1644511149
transform 1 0 24104 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1002_
timestamp 1644511149
transform 1 0 24380 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1003_
timestamp 1644511149
transform -1 0 25852 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1004_
timestamp 1644511149
transform -1 0 19964 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1005_
timestamp 1644511149
transform 1 0 14720 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1006_
timestamp 1644511149
transform 1 0 15640 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1007_
timestamp 1644511149
transform 1 0 13984 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1008_
timestamp 1644511149
transform -1 0 14812 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1009_
timestamp 1644511149
transform 1 0 13800 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1010_
timestamp 1644511149
transform 1 0 13340 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1011_
timestamp 1644511149
transform 1 0 14720 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1012_
timestamp 1644511149
transform -1 0 17664 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1013_
timestamp 1644511149
transform 1 0 18032 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1014_
timestamp 1644511149
transform 1 0 16928 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1015_
timestamp 1644511149
transform 1 0 17296 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1016_
timestamp 1644511149
transform 1 0 22540 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1017_
timestamp 1644511149
transform 1 0 24840 0 -1 30464
box -38 -48 1602 592
use sky130_fd_sc_hd__conb_1  _1018__17 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 6624 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1019__18
timestamp 1644511149
transform -1 0 1748 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1020__19
timestamp 1644511149
transform -1 0 17204 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1021__20
timestamp 1644511149
transform -1 0 1840 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1022__21
timestamp 1644511149
transform 1 0 27876 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1023__22
timestamp 1644511149
transform 1 0 1840 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1024__23
timestamp 1644511149
transform 1 0 27876 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1025__24
timestamp 1644511149
transform 1 0 1472 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1026__25
timestamp 1644511149
transform -1 0 27324 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1027__26
timestamp 1644511149
transform 1 0 25668 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1028__27
timestamp 1644511149
transform 1 0 27232 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1029__28
timestamp 1644511149
transform 1 0 18124 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1030__29
timestamp 1644511149
transform 1 0 26220 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1031__30
timestamp 1644511149
transform -1 0 1748 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1032__31
timestamp 1644511149
transform 1 0 10488 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1033__32
timestamp 1644511149
transform 1 0 2852 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1034__33
timestamp 1644511149
transform 1 0 27876 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1035__34
timestamp 1644511149
transform 1 0 26220 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1036__35
timestamp 1644511149
transform -1 0 1840 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1037__36
timestamp 1644511149
transform 1 0 27876 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1038__37
timestamp 1644511149
transform -1 0 3220 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1039__38
timestamp 1644511149
transform 1 0 27692 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1040__39
timestamp 1644511149
transform -1 0 15272 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1041__40
timestamp 1644511149
transform 1 0 8188 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1042__41
timestamp 1644511149
transform 1 0 27876 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1043__42
timestamp 1644511149
transform 1 0 1380 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1044__43
timestamp 1644511149
transform 1 0 27784 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1045__44
timestamp 1644511149
transform -1 0 1932 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1046__45
timestamp 1644511149
transform -1 0 27324 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1047__46
timestamp 1644511149
transform -1 0 4324 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1048__47
timestamp 1644511149
transform 1 0 26220 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1049__48
timestamp 1644511149
transform 1 0 27876 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1050__49
timestamp 1644511149
transform -1 0 24656 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1051__50
timestamp 1644511149
transform -1 0 16928 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1052__51
timestamp 1644511149
transform -1 0 5520 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1053__52
timestamp 1644511149
transform 1 0 2116 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1054__53
timestamp 1644511149
transform 1 0 27876 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1055__54
timestamp 1644511149
transform -1 0 8096 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1056__55
timestamp 1644511149
transform -1 0 27232 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1057__56
timestamp 1644511149
transform 1 0 2484 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1058__57
timestamp 1644511149
transform -1 0 15364 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1059__58
timestamp 1644511149
transform 1 0 26220 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1060__59
timestamp 1644511149
transform 1 0 27784 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1061__60
timestamp 1644511149
transform -1 0 1748 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1062__61
timestamp 1644511149
transform -1 0 22356 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1063__62
timestamp 1644511149
transform -1 0 1748 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1064__63
timestamp 1644511149
transform -1 0 24656 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1065__64
timestamp 1644511149
transform 1 0 27784 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1066__65
timestamp 1644511149
transform -1 0 22080 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1067__66
timestamp 1644511149
transform -1 0 19688 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1068__67
timestamp 1644511149
transform 1 0 2208 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1069__68
timestamp 1644511149
transform -1 0 20424 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1070__69
timestamp 1644511149
transform 1 0 12420 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1071__70
timestamp 1644511149
transform 1 0 27140 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1072__71
timestamp 1644511149
transform 1 0 4784 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1073__72
timestamp 1644511149
transform -1 0 1748 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1074__73
timestamp 1644511149
transform 1 0 1380 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1075__74
timestamp 1644511149
transform 1 0 24840 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1076__75
timestamp 1644511149
transform -1 0 27324 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1077__76
timestamp 1644511149
transform 1 0 27876 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1078__77
timestamp 1644511149
transform -1 0 3036 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1079__78
timestamp 1644511149
transform 1 0 26128 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1080__79
timestamp 1644511149
transform -1 0 22080 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1081__80
timestamp 1644511149
transform -1 0 27232 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1082__81
timestamp 1644511149
transform -1 0 22908 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1083__82
timestamp 1644511149
transform -1 0 19688 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1084__83
timestamp 1644511149
transform -1 0 27324 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1085__84
timestamp 1644511149
transform -1 0 1748 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1086__85
timestamp 1644511149
transform -1 0 27508 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1087__86
timestamp 1644511149
transform 1 0 1380 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1088__87
timestamp 1644511149
transform -1 0 3128 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1089__88
timestamp 1644511149
transform 1 0 7268 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1090__89
timestamp 1644511149
transform -1 0 1840 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1091__90
timestamp 1644511149
transform 1 0 25576 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1092__91
timestamp 1644511149
transform 1 0 23644 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1093__92
timestamp 1644511149
transform 1 0 23920 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1094__93
timestamp 1644511149
transform -1 0 1840 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1095__94
timestamp 1644511149
transform -1 0 2024 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1096__95
timestamp 1644511149
transform 1 0 25668 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1097__96
timestamp 1644511149
transform 1 0 11408 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1098__97
timestamp 1644511149
transform -1 0 18400 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1099__98
timestamp 1644511149
transform 1 0 2760 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1100__99
timestamp 1644511149
transform 1 0 27876 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1101__100
timestamp 1644511149
transform 1 0 4416 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1102__101
timestamp 1644511149
transform -1 0 4048 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1103__102
timestamp 1644511149
transform -1 0 10396 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1104__103
timestamp 1644511149
transform 1 0 10764 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1105__104
timestamp 1644511149
transform -1 0 27232 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1106__105
timestamp 1644511149
transform 1 0 26220 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1107__106
timestamp 1644511149
transform -1 0 14352 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1108__107
timestamp 1644511149
transform 1 0 27876 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1109__108
timestamp 1644511149
transform 1 0 27232 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1110__109
timestamp 1644511149
transform 1 0 1564 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1111__110
timestamp 1644511149
transform 1 0 26220 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1112__111
timestamp 1644511149
transform 1 0 2116 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1113__112
timestamp 1644511149
transform 1 0 24472 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1114__113
timestamp 1644511149
transform -1 0 4048 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1115__114
timestamp 1644511149
transform -1 0 1656 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1116__115
timestamp 1644511149
transform -1 0 1748 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1117__116
timestamp 1644511149
transform -1 0 1748 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1118_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 6348 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1119_
timestamp 1644511149
transform 1 0 1380 0 1 34816
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1120_
timestamp 1644511149
transform 1 0 16652 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1121_
timestamp 1644511149
transform 1 0 1472 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1122_
timestamp 1644511149
transform -1 0 28244 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1123_
timestamp 1644511149
transform 1 0 2484 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1124_
timestamp 1644511149
transform -1 0 28244 0 1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1125_
timestamp 1644511149
transform 1 0 2116 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1126_
timestamp 1644511149
transform 1 0 26312 0 1 39168
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1127_
timestamp 1644511149
transform 1 0 26312 0 1 43520
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1128_
timestamp 1644511149
transform -1 0 28244 0 1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1129_
timestamp 1644511149
transform -1 0 19964 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1130_
timestamp 1644511149
transform 1 0 26312 0 1 42432
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1131_
timestamp 1644511149
transform 1 0 1380 0 1 43520
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1132_
timestamp 1644511149
transform 1 0 11132 0 1 44608
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1133_
timestamp 1644511149
transform -1 0 3864 0 -1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1134_
timestamp 1644511149
transform -1 0 28244 0 1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1135_
timestamp 1644511149
transform 1 0 26312 0 1 38080
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1136_
timestamp 1644511149
transform 1 0 1564 0 -1 41344
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1137_
timestamp 1644511149
transform -1 0 28244 0 1 30464
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1138_
timestamp 1644511149
transform 1 0 2944 0 -1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1139_
timestamp 1644511149
transform -1 0 28244 0 1 44608
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1140_
timestamp 1644511149
transform 1 0 14260 0 1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1141_
timestamp 1644511149
transform 1 0 9108 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1142_
timestamp 1644511149
transform -1 0 28244 0 1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1143_
timestamp 1644511149
transform 1 0 1656 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1144_
timestamp 1644511149
transform -1 0 28244 0 1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1145_
timestamp 1644511149
transform 1 0 1380 0 1 38080
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1146_
timestamp 1644511149
transform 1 0 26312 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1147_
timestamp 1644511149
transform 1 0 3956 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1148_
timestamp 1644511149
transform 1 0 26312 0 1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1149_
timestamp 1644511149
transform -1 0 28244 0 1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1150_
timestamp 1644511149
transform 1 0 23736 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1151_
timestamp 1644511149
transform 1 0 16652 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1152_
timestamp 1644511149
transform 1 0 5152 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1153_
timestamp 1644511149
transform -1 0 3680 0 -1 34816
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1154_
timestamp 1644511149
transform -1 0 28244 0 1 33728
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1155_
timestamp 1644511149
transform 1 0 7820 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1156_
timestamp 1644511149
transform -1 0 26496 0 1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1157_
timestamp 1644511149
transform -1 0 4416 0 -1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1158_
timestamp 1644511149
transform 1 0 14260 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1159_
timestamp 1644511149
transform -1 0 26496 0 1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1160_
timestamp 1644511149
transform 1 0 26312 0 1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1161_
timestamp 1644511149
transform -1 0 27048 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1162_
timestamp 1644511149
transform -1 0 26496 0 -1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1163_
timestamp 1644511149
transform 1 0 26312 0 1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1164_
timestamp 1644511149
transform 1 0 26312 0 1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1165_
timestamp 1644511149
transform -1 0 27508 0 1 31552
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1166_
timestamp 1644511149
transform 1 0 26312 0 1 29376
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1167_
timestamp 1644511149
transform 1 0 26312 0 1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1168_
timestamp 1644511149
transform -1 0 28244 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1169_
timestamp 1644511149
transform 1 0 1380 0 -1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1170_
timestamp 1644511149
transform 1 0 21988 0 1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1171_
timestamp 1644511149
transform 1 0 1380 0 1 31552
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1172_
timestamp 1644511149
transform 1 0 24012 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1173_
timestamp 1644511149
transform -1 0 28244 0 1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1174_
timestamp 1644511149
transform 1 0 21252 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1175_
timestamp 1644511149
transform 1 0 19412 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1176_
timestamp 1644511149
transform -1 0 3312 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1177_
timestamp 1644511149
transform 1 0 19688 0 1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1178_
timestamp 1644511149
transform 1 0 12972 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1179_
timestamp 1644511149
transform -1 0 28244 0 1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1180_
timestamp 1644511149
transform -1 0 6348 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1181_
timestamp 1644511149
transform 1 0 1472 0 -1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1182_
timestamp 1644511149
transform -1 0 3312 0 1 36992
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1183_
timestamp 1644511149
transform 1 0 26312 0 1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1184_
timestamp 1644511149
transform 1 0 26312 0 1 41344
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1185_
timestamp 1644511149
transform -1 0 28244 0 1 40256
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1186_
timestamp 1644511149
transform 1 0 2484 0 -1 43520
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1187_
timestamp 1644511149
transform -1 0 26496 0 -1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1188_
timestamp 1644511149
transform 1 0 20700 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1189_
timestamp 1644511149
transform 1 0 26312 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1190_
timestamp 1644511149
transform 1 0 21988 0 1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1191_
timestamp 1644511149
transform 1 0 19412 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1192_
timestamp 1644511149
transform -1 0 26496 0 -1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1193_
timestamp 1644511149
transform 1 0 1380 0 1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1194_
timestamp 1644511149
transform -1 0 26496 0 -1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1195_
timestamp 1644511149
transform 1 0 1564 0 -1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1196_
timestamp 1644511149
transform 1 0 2852 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1197_
timestamp 1644511149
transform 1 0 8648 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1198_
timestamp 1644511149
transform 1 0 1472 0 -1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1199_
timestamp 1644511149
transform -1 0 26496 0 -1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1200_
timestamp 1644511149
transform 1 0 26312 0 1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1201_
timestamp 1644511149
transform 1 0 24564 0 -1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1202_
timestamp 1644511149
transform 1 0 1380 0 1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1203_
timestamp 1644511149
transform 1 0 1656 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1204_
timestamp 1644511149
transform 1 0 26312 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1205_
timestamp 1644511149
transform 1 0 11500 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1206_
timestamp 1644511149
transform 1 0 18124 0 -1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1207_
timestamp 1644511149
transform 1 0 3956 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1208_
timestamp 1644511149
transform -1 0 28244 0 1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1209_
timestamp 1644511149
transform -1 0 4692 0 -1 42432
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1210_
timestamp 1644511149
transform 1 0 3772 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1211_
timestamp 1644511149
transform 1 0 9568 0 1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1212_
timestamp 1644511149
transform 1 0 11500 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1213_
timestamp 1644511149
transform -1 0 26496 0 -1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1214_
timestamp 1644511149
transform -1 0 26496 0 -1 41344
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1215_
timestamp 1644511149
transform 1 0 13800 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1216_
timestamp 1644511149
transform -1 0 28244 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1217_
timestamp 1644511149
transform -1 0 28244 0 1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1218_
timestamp 1644511149
transform -1 0 3312 0 1 41344
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1219_
timestamp 1644511149
transform -1 0 26496 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1220_
timestamp 1644511149
transform 1 0 2300 0 -1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1221_
timestamp 1644511149
transform 1 0 24564 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1222_
timestamp 1644511149
transform 1 0 3772 0 1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1223_
timestamp 1644511149
transform 1 0 1380 0 1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1224_
timestamp 1644511149
transform 1 0 1380 0 1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1225_
timestamp 1644511149
transform 1 0 1380 0 1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_wb_clk_i $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 21344 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_2_0_0_wb_clk_i
timestamp 1644511149
transform -1 0 18124 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_2_1_0_wb_clk_i
timestamp 1644511149
transform -1 0 20792 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_2_2_0_wb_clk_i
timestamp 1644511149
transform -1 0 19596 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_2_3_0_wb_clk_i
timestamp 1644511149
transform 1 0 22908 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 27692 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold2 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 25852 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_4  input1
timestamp 1644511149
transform 1 0 1748 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1644511149
transform 1 0 26588 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input3
timestamp 1644511149
transform -1 0 28244 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1644511149
transform 1 0 17480 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1644511149
transform 1 0 24564 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1644511149
transform -1 0 1656 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input7
timestamp 1644511149
transform 1 0 27140 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  input8
timestamp 1644511149
transform 1 0 16652 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input9
timestamp 1644511149
transform 1 0 9292 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1644511149
transform -1 0 1656 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input11
timestamp 1644511149
transform -1 0 23368 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1644511149
transform 1 0 27140 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input13
timestamp 1644511149
transform 1 0 6348 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1644511149
transform -1 0 2668 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input15
timestamp 1644511149
transform 1 0 7084 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input16
timestamp 1644511149
transform -1 0 1656 0 -1 28288
box -38 -48 314 592
<< labels >>
rlabel metal3 s 0 36668 800 36908 6 active
port 0 nsew signal input
rlabel metal2 s 12226 0 12338 800 6 io_in[0]
port 1 nsew signal input
rlabel metal2 s 12226 49200 12338 50000 6 io_in[10]
port 2 nsew signal input
rlabel metal3 s 0 40068 800 40308 6 io_in[11]
port 3 nsew signal input
rlabel metal3 s 29200 43468 30000 43708 6 io_in[12]
port 4 nsew signal input
rlabel metal2 s 18666 0 18778 800 6 io_in[13]
port 5 nsew signal input
rlabel metal2 s 5142 49200 5254 50000 6 io_in[14]
port 6 nsew signal input
rlabel metal3 s 29200 45508 30000 45748 6 io_in[15]
port 7 nsew signal input
rlabel metal3 s 29200 13548 30000 13788 6 io_in[16]
port 8 nsew signal input
rlabel metal3 s 0 48228 800 48468 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s -10 49200 102 50000 6 io_in[18]
port 10 nsew signal input
rlabel metal3 s 29200 4028 30000 4268 6 io_in[19]
port 11 nsew signal input
rlabel metal3 s 0 12868 800 13108 6 io_in[1]
port 12 nsew signal input
rlabel metal3 s 0 23068 800 23308 6 io_in[20]
port 13 nsew signal input
rlabel metal3 s 0 14908 800 15148 6 io_in[21]
port 14 nsew signal input
rlabel metal3 s 29200 23068 30000 23308 6 io_in[22]
port 15 nsew signal input
rlabel metal3 s 0 47548 800 47788 6 io_in[23]
port 16 nsew signal input
rlabel metal3 s 0 45508 800 45748 6 io_in[24]
port 17 nsew signal input
rlabel metal2 s 29614 0 29726 800 6 io_in[25]
port 18 nsew signal input
rlabel metal2 s 28970 0 29082 800 6 io_in[26]
port 19 nsew signal input
rlabel metal3 s 29200 18988 30000 19228 6 io_in[27]
port 20 nsew signal input
rlabel metal2 s 26394 0 26506 800 6 io_in[28]
port 21 nsew signal input
rlabel metal2 s 29614 49200 29726 50000 6 io_in[29]
port 22 nsew signal input
rlabel metal2 s 12870 0 12982 800 6 io_in[2]
port 23 nsew signal input
rlabel metal3 s 29200 25788 30000 26028 6 io_in[30]
port 24 nsew signal input
rlabel metal3 s 0 35308 800 35548 6 io_in[31]
port 25 nsew signal input
rlabel metal2 s 24462 0 24574 800 6 io_in[32]
port 26 nsew signal input
rlabel metal3 s 0 20348 800 20588 6 io_in[33]
port 27 nsew signal input
rlabel metal2 s 20598 49200 20710 50000 6 io_in[34]
port 28 nsew signal input
rlabel metal2 s 25106 49200 25218 50000 6 io_in[35]
port 29 nsew signal input
rlabel metal3 s 29200 35308 30000 35548 6 io_in[36]
port 30 nsew signal input
rlabel metal2 s 25750 49200 25862 50000 6 io_in[37]
port 31 nsew signal input
rlabel metal2 s 12870 49200 12982 50000 6 io_in[3]
port 32 nsew signal input
rlabel metal3 s 29200 34628 30000 34868 6 io_in[4]
port 33 nsew signal input
rlabel metal3 s 29200 48228 30000 48468 6 io_in[5]
port 34 nsew signal input
rlabel metal3 s 0 24428 800 24668 6 io_in[6]
port 35 nsew signal input
rlabel metal3 s 0 16948 800 17188 6 io_in[7]
port 36 nsew signal input
rlabel metal3 s 29200 36668 30000 36908 6 io_in[8]
port 37 nsew signal input
rlabel metal3 s 0 46868 800 47108 6 io_in[9]
port 38 nsew signal input
rlabel metal2 s 21242 0 21354 800 6 io_oeb[0]
port 39 nsew signal tristate
rlabel metal3 s 0 13548 800 13788 6 io_oeb[10]
port 40 nsew signal tristate
rlabel metal3 s 29200 32588 30000 32828 6 io_oeb[11]
port 41 nsew signal tristate
rlabel metal3 s 29200 21708 30000 21948 6 io_oeb[12]
port 42 nsew signal tristate
rlabel metal3 s 29200 21028 30000 21268 6 io_oeb[13]
port 43 nsew signal tristate
rlabel metal3 s 0 3348 800 3588 6 io_oeb[14]
port 44 nsew signal tristate
rlabel metal2 s 1278 49200 1390 50000 6 io_oeb[15]
port 45 nsew signal tristate
rlabel metal3 s 29200 12188 30000 12428 6 io_oeb[16]
port 46 nsew signal tristate
rlabel metal2 s 10938 0 11050 800 6 io_oeb[17]
port 47 nsew signal tristate
rlabel metal2 s 18666 49200 18778 50000 6 io_oeb[18]
port 48 nsew signal tristate
rlabel metal2 s 1922 49200 2034 50000 6 io_oeb[19]
port 49 nsew signal tristate
rlabel metal3 s 29200 1308 30000 1548 6 io_oeb[1]
port 50 nsew signal tristate
rlabel metal3 s 29200 27148 30000 27388 6 io_oeb[20]
port 51 nsew signal tristate
rlabel metal3 s 0 41428 800 41668 6 io_oeb[21]
port 52 nsew signal tristate
rlabel metal2 s 3854 0 3966 800 6 io_oeb[22]
port 53 nsew signal tristate
rlabel metal2 s 10294 49200 10406 50000 6 io_oeb[23]
port 54 nsew signal tristate
rlabel metal2 s 10938 49200 11050 50000 6 io_oeb[24]
port 55 nsew signal tristate
rlabel metal3 s 29200 8108 30000 8348 6 io_oeb[25]
port 56 nsew signal tristate
rlabel metal3 s 29200 41428 30000 41668 6 io_oeb[26]
port 57 nsew signal tristate
rlabel metal2 s 13514 49200 13626 50000 6 io_oeb[27]
port 58 nsew signal tristate
rlabel metal3 s 29200 3348 30000 3588 6 io_oeb[28]
port 59 nsew signal tristate
rlabel metal3 s 29200 35988 30000 36228 6 io_oeb[29]
port 60 nsew signal tristate
rlabel metal2 s 23174 49200 23286 50000 6 io_oeb[2]
port 61 nsew signal tristate
rlabel metal3 s 0 42108 800 42348 6 io_oeb[30]
port 62 nsew signal tristate
rlabel metal3 s 29200 2668 30000 2908 6 io_oeb[31]
port 63 nsew signal tristate
rlabel metal3 s 0 19668 800 19908 6 io_oeb[32]
port 64 nsew signal tristate
rlabel metal3 s 29200 8788 30000 9028 6 io_oeb[33]
port 65 nsew signal tristate
rlabel metal3 s 0 49588 800 49828 6 io_oeb[34]
port 66 nsew signal tristate
rlabel metal3 s 0 17628 800 17868 6 io_oeb[35]
port 67 nsew signal tristate
rlabel metal3 s 0 8788 800 9028 6 io_oeb[36]
port 68 nsew signal tristate
rlabel metal3 s 0 14228 800 14468 6 io_oeb[37]
port 69 nsew signal tristate
rlabel metal2 s 19954 0 20066 800 6 io_oeb[3]
port 70 nsew signal tristate
rlabel metal3 s 29200 10148 30000 10388 6 io_oeb[4]
port 71 nsew signal tristate
rlabel metal3 s 0 25788 800 26028 6 io_oeb[5]
port 72 nsew signal tristate
rlabel metal3 s 29200 24428 30000 24668 6 io_oeb[6]
port 73 nsew signal tristate
rlabel metal2 s 634 49200 746 50000 6 io_oeb[7]
port 74 nsew signal tristate
rlabel metal2 s 3210 0 3322 800 6 io_oeb[8]
port 75 nsew signal tristate
rlabel metal2 s 8362 0 8474 800 6 io_oeb[9]
port 76 nsew signal tristate
rlabel metal3 s 29200 47548 30000 47788 6 io_out[0]
port 77 nsew signal tristate
rlabel metal3 s 29200 31908 30000 32148 6 io_out[10]
port 78 nsew signal tristate
rlabel metal3 s 0 1988 800 2228 6 io_out[11]
port 79 nsew signal tristate
rlabel metal3 s 0 6068 800 6308 6 io_out[12]
port 80 nsew signal tristate
rlabel metal3 s 29200 1988 30000 2228 6 io_out[13]
port 81 nsew signal tristate
rlabel metal3 s 29200 42108 30000 42348 6 io_out[14]
port 82 nsew signal tristate
rlabel metal3 s 0 33268 800 33508 6 io_out[15]
port 83 nsew signal tristate
rlabel metal3 s 29200 31228 30000 31468 6 io_out[16]
port 84 nsew signal tristate
rlabel metal2 s 27038 49200 27150 50000 6 io_out[17]
port 85 nsew signal tristate
rlabel metal3 s 29200 7428 30000 7668 6 io_out[18]
port 86 nsew signal tristate
rlabel metal3 s 0 18988 800 19228 6 io_out[19]
port 87 nsew signal tristate
rlabel metal2 s 16734 49200 16846 50000 6 io_out[1]
port 88 nsew signal tristate
rlabel metal2 s 22530 49200 22642 50000 6 io_out[20]
port 89 nsew signal tristate
rlabel metal3 s 0 31908 800 32148 6 io_out[21]
port 90 nsew signal tristate
rlabel metal2 s 25106 0 25218 800 6 io_out[22]
port 91 nsew signal tristate
rlabel metal3 s 29200 28508 30000 28748 6 io_out[23]
port 92 nsew signal tristate
rlabel metal2 s 21886 0 21998 800 6 io_out[24]
port 93 nsew signal tristate
rlabel metal2 s 19954 49200 20066 50000 6 io_out[25]
port 94 nsew signal tristate
rlabel metal3 s 0 4028 800 4268 6 io_out[26]
port 95 nsew signal tristate
rlabel metal2 s 21242 49200 21354 50000 6 io_out[27]
port 96 nsew signal tristate
rlabel metal2 s 13514 0 13626 800 6 io_out[28]
port 97 nsew signal tristate
rlabel metal3 s 29200 10828 30000 11068 6 io_out[29]
port 98 nsew signal tristate
rlabel metal2 s 5786 0 5898 800 6 io_out[2]
port 99 nsew signal tristate
rlabel metal3 s 0 4708 800 4948 6 io_out[30]
port 100 nsew signal tristate
rlabel metal3 s 0 11508 800 11748 6 io_out[31]
port 101 nsew signal tristate
rlabel metal3 s 0 37348 800 37588 6 io_out[32]
port 102 nsew signal tristate
rlabel metal3 s 29200 15588 30000 15828 6 io_out[33]
port 103 nsew signal tristate
rlabel metal3 s 29200 42788 30000 43028 6 io_out[34]
port 104 nsew signal tristate
rlabel metal3 s 29200 40748 30000 40988 6 io_out[35]
port 105 nsew signal tristate
rlabel metal2 s 2566 49200 2678 50000 6 io_out[36]
port 106 nsew signal tristate
rlabel metal3 s 29200 46188 30000 46428 6 io_out[37]
port 107 nsew signal tristate
rlabel metal3 s 0 34628 800 34868 6 io_out[3]
port 108 nsew signal tristate
rlabel metal3 s 29200 33948 30000 34188 6 io_out[4]
port 109 nsew signal tristate
rlabel metal2 s 8362 49200 8474 50000 6 io_out[5]
port 110 nsew signal tristate
rlabel metal2 s 28326 49200 28438 50000 6 io_out[6]
port 111 nsew signal tristate
rlabel metal3 s 0 15588 800 15828 6 io_out[7]
port 112 nsew signal tristate
rlabel metal2 s 14802 0 14914 800 6 io_out[8]
port 113 nsew signal tristate
rlabel metal3 s 0 12188 800 12428 6 io_out[9]
port 114 nsew signal tristate
rlabel metal3 s 29200 16268 30000 16508 6 la1_data_in[0]
port 115 nsew signal input
rlabel metal2 s 17378 0 17490 800 6 la1_data_in[10]
port 116 nsew signal input
rlabel metal3 s 29200 14908 30000 15148 6 la1_data_in[11]
port 117 nsew signal input
rlabel metal3 s 0 29868 800 30108 6 la1_data_in[12]
port 118 nsew signal input
rlabel metal2 s 27038 0 27150 800 6 la1_data_in[13]
port 119 nsew signal input
rlabel metal3 s 0 10148 800 10388 6 la1_data_in[14]
port 120 nsew signal input
rlabel metal2 s 3210 49200 3322 50000 6 la1_data_in[15]
port 121 nsew signal input
rlabel metal2 s 15446 49200 15558 50000 6 la1_data_in[16]
port 122 nsew signal input
rlabel metal2 s 9650 49200 9762 50000 6 la1_data_in[17]
port 123 nsew signal input
rlabel metal3 s 29200 4708 30000 4948 6 la1_data_in[18]
port 124 nsew signal input
rlabel metal2 s 4498 49200 4610 50000 6 la1_data_in[19]
port 125 nsew signal input
rlabel metal2 s 16090 0 16202 800 6 la1_data_in[1]
port 126 nsew signal input
rlabel metal3 s 0 29188 800 29428 6 la1_data_in[20]
port 127 nsew signal input
rlabel metal2 s 28970 49200 29082 50000 6 la1_data_in[21]
port 128 nsew signal input
rlabel metal3 s 29200 17628 30000 17868 6 la1_data_in[22]
port 129 nsew signal input
rlabel metal3 s 0 628 800 868 6 la1_data_in[23]
port 130 nsew signal input
rlabel metal2 s 11582 0 11694 800 6 la1_data_in[24]
port 131 nsew signal input
rlabel metal3 s 0 30548 800 30788 6 la1_data_in[25]
port 132 nsew signal input
rlabel metal3 s 29200 12868 30000 13108 6 la1_data_in[26]
port 133 nsew signal input
rlabel metal2 s 23174 0 23286 800 6 la1_data_in[27]
port 134 nsew signal input
rlabel metal3 s 0 26468 800 26708 6 la1_data_in[28]
port 135 nsew signal input
rlabel metal3 s 0 40748 800 40988 6 la1_data_in[29]
port 136 nsew signal input
rlabel metal2 s 9006 0 9118 800 6 la1_data_in[2]
port 137 nsew signal input
rlabel metal2 s 1278 0 1390 800 6 la1_data_in[30]
port 138 nsew signal input
rlabel metal3 s 29200 -52 30000 188 6 la1_data_in[31]
port 139 nsew signal input
rlabel metal3 s 0 25108 800 25348 6 la1_data_in[3]
port 140 nsew signal input
rlabel metal2 s 23818 49200 23930 50000 6 la1_data_in[4]
port 141 nsew signal input
rlabel metal3 s 29200 29868 30000 30108 6 la1_data_in[5]
port 142 nsew signal input
rlabel metal2 s 5786 49200 5898 50000 6 la1_data_in[6]
port 143 nsew signal input
rlabel metal3 s 0 18308 800 18548 6 la1_data_in[7]
port 144 nsew signal input
rlabel metal2 s 6430 49200 6542 50000 6 la1_data_in[8]
port 145 nsew signal input
rlabel metal3 s 0 27828 800 28068 6 la1_data_in[9]
port 146 nsew signal input
rlabel metal2 s 6430 0 6542 800 6 la1_data_out[0]
port 147 nsew signal tristate
rlabel metal3 s 29200 19668 30000 19908 6 la1_data_out[10]
port 148 nsew signal tristate
rlabel metal2 s 18022 0 18134 800 6 la1_data_out[11]
port 149 nsew signal tristate
rlabel metal3 s 29200 46868 30000 47108 6 la1_data_out[12]
port 150 nsew signal tristate
rlabel metal3 s 0 44148 800 44388 6 la1_data_out[13]
port 151 nsew signal tristate
rlabel metal2 s 11582 49200 11694 50000 6 la1_data_out[14]
port 152 nsew signal tristate
rlabel metal3 s 0 1308 800 1548 6 la1_data_out[15]
port 153 nsew signal tristate
rlabel metal3 s 29200 23748 30000 23988 6 la1_data_out[16]
port 154 nsew signal tristate
rlabel metal3 s 29200 39388 30000 39628 6 la1_data_out[17]
port 155 nsew signal tristate
rlabel metal3 s 0 44828 800 45068 6 la1_data_out[18]
port 156 nsew signal tristate
rlabel metal3 s 29200 30548 30000 30788 6 la1_data_out[19]
port 157 nsew signal tristate
rlabel metal3 s 0 35988 800 36228 6 la1_data_out[1]
port 158 nsew signal tristate
rlabel metal3 s 0 8108 800 8348 6 la1_data_out[20]
port 159 nsew signal tristate
rlabel metal3 s 29200 44828 30000 45068 6 la1_data_out[21]
port 160 nsew signal tristate
rlabel metal2 s 14802 49200 14914 50000 6 la1_data_out[22]
port 161 nsew signal tristate
rlabel metal2 s 9650 0 9762 800 6 la1_data_out[23]
port 162 nsew signal tristate
rlabel metal3 s 29200 25108 30000 25348 6 la1_data_out[24]
port 163 nsew signal tristate
rlabel metal3 s 0 2668 800 2908 6 la1_data_out[25]
port 164 nsew signal tristate
rlabel metal3 s 29200 14228 30000 14468 6 la1_data_out[26]
port 165 nsew signal tristate
rlabel metal3 s 0 38708 800 38948 6 la1_data_out[27]
port 166 nsew signal tristate
rlabel metal3 s 29200 5388 30000 5628 6 la1_data_out[28]
port 167 nsew signal tristate
rlabel metal2 s 4498 0 4610 800 6 la1_data_out[29]
port 168 nsew signal tristate
rlabel metal2 s 16734 0 16846 800 6 la1_data_out[2]
port 169 nsew signal tristate
rlabel metal3 s 29200 20348 30000 20588 6 la1_data_out[30]
port 170 nsew signal tristate
rlabel metal3 s 29200 48908 30000 49148 6 la1_data_out[31]
port 171 nsew signal tristate
rlabel metal3 s 0 7428 800 7668 6 la1_data_out[3]
port 172 nsew signal tristate
rlabel metal3 s 29200 6748 30000 6988 6 la1_data_out[4]
port 173 nsew signal tristate
rlabel metal2 s 2566 0 2678 800 6 la1_data_out[5]
port 174 nsew signal tristate
rlabel metal3 s 29200 26468 30000 26708 6 la1_data_out[6]
port 175 nsew signal tristate
rlabel metal2 s 634 0 746 800 6 la1_data_out[7]
port 176 nsew signal tristate
rlabel metal3 s 29200 40068 30000 40308 6 la1_data_out[8]
port 177 nsew signal tristate
rlabel metal2 s 27682 49200 27794 50000 6 la1_data_out[9]
port 178 nsew signal tristate
rlabel metal3 s 29200 9468 30000 9708 6 la1_oenb[0]
port 179 nsew signal input
rlabel metal2 s 26394 49200 26506 50000 6 la1_oenb[10]
port 180 nsew signal input
rlabel metal3 s 0 22388 800 22628 6 la1_oenb[11]
port 181 nsew signal input
rlabel metal3 s 0 23748 800 23988 6 la1_oenb[12]
port 182 nsew signal input
rlabel metal2 s 23818 0 23930 800 6 la1_oenb[13]
port 183 nsew signal input
rlabel metal2 s -10 0 102 800 6 la1_oenb[14]
port 184 nsew signal input
rlabel metal2 s 28326 0 28438 800 6 la1_oenb[15]
port 185 nsew signal input
rlabel metal3 s 0 28508 800 28748 6 la1_oenb[16]
port 186 nsew signal input
rlabel metal3 s 0 42788 800 43028 6 la1_oenb[17]
port 187 nsew signal input
rlabel metal2 s 7718 49200 7830 50000 6 la1_oenb[18]
port 188 nsew signal input
rlabel metal3 s 0 21028 800 21268 6 la1_oenb[19]
port 189 nsew signal input
rlabel metal2 s 7074 0 7186 800 6 la1_oenb[1]
port 190 nsew signal input
rlabel metal2 s 1922 0 2034 800 6 la1_oenb[20]
port 191 nsew signal input
rlabel metal2 s 16090 49200 16202 50000 6 la1_oenb[21]
port 192 nsew signal input
rlabel metal2 s 7074 49200 7186 50000 6 la1_oenb[22]
port 193 nsew signal input
rlabel metal2 s 19310 0 19422 800 6 la1_oenb[23]
port 194 nsew signal input
rlabel metal2 s 21886 49200 21998 50000 6 la1_oenb[24]
port 195 nsew signal input
rlabel metal3 s 29200 18308 30000 18548 6 la1_oenb[25]
port 196 nsew signal input
rlabel metal3 s 0 31228 800 31468 6 la1_oenb[26]
port 197 nsew signal input
rlabel metal3 s 29200 38028 30000 38268 6 la1_oenb[27]
port 198 nsew signal input
rlabel metal2 s 7718 0 7830 800 6 la1_oenb[28]
port 199 nsew signal input
rlabel metal2 s 14158 0 14270 800 6 la1_oenb[29]
port 200 nsew signal input
rlabel metal3 s 0 6748 800 6988 6 la1_oenb[2]
port 201 nsew signal input
rlabel metal3 s 29200 37348 30000 37588 6 la1_oenb[30]
port 202 nsew signal input
rlabel metal2 s 22530 0 22642 800 6 la1_oenb[31]
port 203 nsew signal input
rlabel metal2 s 18022 49200 18134 50000 6 la1_oenb[3]
port 204 nsew signal input
rlabel metal2 s 17378 49200 17490 50000 6 la1_oenb[4]
port 205 nsew signal input
rlabel metal3 s 0 39388 800 39628 6 la1_oenb[5]
port 206 nsew signal input
rlabel metal3 s 0 46188 800 46428 6 la1_oenb[6]
port 207 nsew signal input
rlabel metal2 s 27682 0 27794 800 6 la1_oenb[7]
port 208 nsew signal input
rlabel metal3 s 0 9468 800 9708 6 la1_oenb[8]
port 209 nsew signal input
rlabel metal3 s 0 33948 800 34188 6 la1_oenb[9]
port 210 nsew signal input
rlabel metal4 s 5576 2128 5896 47376 6 vccd1
port 211 nsew power input
rlabel metal4 s 14840 2128 15160 47376 6 vccd1
port 211 nsew power input
rlabel metal4 s 24104 2128 24424 47376 6 vccd1
port 211 nsew power input
rlabel metal4 s 10208 2128 10528 47376 6 vssd1
port 212 nsew ground input
rlabel metal4 s 19472 2128 19792 47376 6 vssd1
port 212 nsew ground input
rlabel metal3 s 29200 29188 30000 29428 6 wb_clk_i
port 213 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 30000 50000
<< end >>
